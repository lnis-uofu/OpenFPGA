//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Top-level Verilog module for FPGA
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Sun May  3 00:45:58 2020
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

// ----- Verilog module for fpga_top -----
module fpga_core(pReset,
                prog_clk,
                Reset,
                Test_en,
		clk,
lut4_out_0, lut4_out_1, lut4_out_2, lut4_out_3, lut5_out_0, lut5_out_1, lut6_out_0, sc_head, sc_tail, cc_spypad_0, cc_spypad_1, cc_spypad_2, sc_spypad_0, shiftreg_spypad_0, cout_spypad_0, perf_spypad_0,


                gfpga_pad_GPIO_A,
                gfpga_pad_GPIO_IE,
                gfpga_pad_GPIO_OE,
                gfpga_pad_GPIO_Y,
                ccff_head,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] pReset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- GLOBAL PORTS -----
input [0:0] Reset;
//----- GLOBAL PORTS -----
input [0:0] Test_en;
//----- GLOBAL PORTS -----
input [0:0] clk;
//----- GPOUT PORTS -----
wire [0:3] gfpga_pad_frac_lut6_spypad_lut4_spy;
//----- GPOUT PORTS -----
wire [0:1] gfpga_pad_frac_lut6_spypad_lut5_spy;
//----- GPOUT PORTS -----
wire [0:0] gfpga_pad_frac_lut6_spypad_lut6_spy;
//----- GPOUT PORTS -----
output [0:7] gfpga_pad_GPIO_A;
//----- GPOUT PORTS -----
output [0:7] gfpga_pad_GPIO_IE;
//----- GPOUT PORTS -----
output [0:7] gfpga_pad_GPIO_OE;
//----- GPIO PORTS -----
inout [0:7] gfpga_pad_GPIO_Y;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;


output [0:0] lut4_out_0; output [0:0] lut4_out_1; output [0:0] lut4_out_2; output [0:0] lut4_out_3; output [0:0] lut5_out_0; output [0:0] lut5_out_1; output [0:0] lut6_out_0; input [0:0] sc_head; output [0:0] sc_tail; output [0:0] cc_spypad_0; output [0:0] cc_spypad_1; output [0:0] cc_spypad_2; output [0:0] sc_spypad_0; output [0:0] shiftreg_spypad_0; output [0:0] cout_spypad_0; output [0:0] perf_spypad_0;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:0] cbx_1__0__0_bottom_grid_pin_0_;
wire [0:0] cbx_1__0__0_ccff_tail;
wire [0:0] cbx_1__0__0_chanx_out_0_;
wire [0:0] cbx_1__0__0_chanx_out_100_;
wire [0:0] cbx_1__0__0_chanx_out_101_;
wire [0:0] cbx_1__0__0_chanx_out_102_;
wire [0:0] cbx_1__0__0_chanx_out_103_;
wire [0:0] cbx_1__0__0_chanx_out_104_;
wire [0:0] cbx_1__0__0_chanx_out_105_;
wire [0:0] cbx_1__0__0_chanx_out_106_;
wire [0:0] cbx_1__0__0_chanx_out_107_;
wire [0:0] cbx_1__0__0_chanx_out_108_;
wire [0:0] cbx_1__0__0_chanx_out_109_;
wire [0:0] cbx_1__0__0_chanx_out_10_;
wire [0:0] cbx_1__0__0_chanx_out_110_;
wire [0:0] cbx_1__0__0_chanx_out_111_;
wire [0:0] cbx_1__0__0_chanx_out_112_;
wire [0:0] cbx_1__0__0_chanx_out_113_;
wire [0:0] cbx_1__0__0_chanx_out_114_;
wire [0:0] cbx_1__0__0_chanx_out_115_;
wire [0:0] cbx_1__0__0_chanx_out_116_;
wire [0:0] cbx_1__0__0_chanx_out_117_;
wire [0:0] cbx_1__0__0_chanx_out_118_;
wire [0:0] cbx_1__0__0_chanx_out_119_;
wire [0:0] cbx_1__0__0_chanx_out_11_;
wire [0:0] cbx_1__0__0_chanx_out_120_;
wire [0:0] cbx_1__0__0_chanx_out_121_;
wire [0:0] cbx_1__0__0_chanx_out_122_;
wire [0:0] cbx_1__0__0_chanx_out_123_;
wire [0:0] cbx_1__0__0_chanx_out_124_;
wire [0:0] cbx_1__0__0_chanx_out_125_;
wire [0:0] cbx_1__0__0_chanx_out_126_;
wire [0:0] cbx_1__0__0_chanx_out_127_;
wire [0:0] cbx_1__0__0_chanx_out_128_;
wire [0:0] cbx_1__0__0_chanx_out_129_;
wire [0:0] cbx_1__0__0_chanx_out_12_;
wire [0:0] cbx_1__0__0_chanx_out_130_;
wire [0:0] cbx_1__0__0_chanx_out_131_;
wire [0:0] cbx_1__0__0_chanx_out_132_;
wire [0:0] cbx_1__0__0_chanx_out_133_;
wire [0:0] cbx_1__0__0_chanx_out_134_;
wire [0:0] cbx_1__0__0_chanx_out_135_;
wire [0:0] cbx_1__0__0_chanx_out_136_;
wire [0:0] cbx_1__0__0_chanx_out_137_;
wire [0:0] cbx_1__0__0_chanx_out_138_;
wire [0:0] cbx_1__0__0_chanx_out_139_;
wire [0:0] cbx_1__0__0_chanx_out_13_;
wire [0:0] cbx_1__0__0_chanx_out_140_;
wire [0:0] cbx_1__0__0_chanx_out_141_;
wire [0:0] cbx_1__0__0_chanx_out_142_;
wire [0:0] cbx_1__0__0_chanx_out_143_;
wire [0:0] cbx_1__0__0_chanx_out_144_;
wire [0:0] cbx_1__0__0_chanx_out_145_;
wire [0:0] cbx_1__0__0_chanx_out_146_;
wire [0:0] cbx_1__0__0_chanx_out_147_;
wire [0:0] cbx_1__0__0_chanx_out_148_;
wire [0:0] cbx_1__0__0_chanx_out_149_;
wire [0:0] cbx_1__0__0_chanx_out_14_;
wire [0:0] cbx_1__0__0_chanx_out_150_;
wire [0:0] cbx_1__0__0_chanx_out_151_;
wire [0:0] cbx_1__0__0_chanx_out_152_;
wire [0:0] cbx_1__0__0_chanx_out_153_;
wire [0:0] cbx_1__0__0_chanx_out_154_;
wire [0:0] cbx_1__0__0_chanx_out_155_;
wire [0:0] cbx_1__0__0_chanx_out_156_;
wire [0:0] cbx_1__0__0_chanx_out_157_;
wire [0:0] cbx_1__0__0_chanx_out_158_;
wire [0:0] cbx_1__0__0_chanx_out_159_;
wire [0:0] cbx_1__0__0_chanx_out_15_;
wire [0:0] cbx_1__0__0_chanx_out_160_;
wire [0:0] cbx_1__0__0_chanx_out_161_;
wire [0:0] cbx_1__0__0_chanx_out_162_;
wire [0:0] cbx_1__0__0_chanx_out_163_;
wire [0:0] cbx_1__0__0_chanx_out_164_;
wire [0:0] cbx_1__0__0_chanx_out_165_;
wire [0:0] cbx_1__0__0_chanx_out_166_;
wire [0:0] cbx_1__0__0_chanx_out_167_;
wire [0:0] cbx_1__0__0_chanx_out_168_;
wire [0:0] cbx_1__0__0_chanx_out_169_;
wire [0:0] cbx_1__0__0_chanx_out_16_;
wire [0:0] cbx_1__0__0_chanx_out_170_;
wire [0:0] cbx_1__0__0_chanx_out_171_;
wire [0:0] cbx_1__0__0_chanx_out_172_;
wire [0:0] cbx_1__0__0_chanx_out_173_;
wire [0:0] cbx_1__0__0_chanx_out_174_;
wire [0:0] cbx_1__0__0_chanx_out_175_;
wire [0:0] cbx_1__0__0_chanx_out_176_;
wire [0:0] cbx_1__0__0_chanx_out_177_;
wire [0:0] cbx_1__0__0_chanx_out_178_;
wire [0:0] cbx_1__0__0_chanx_out_179_;
wire [0:0] cbx_1__0__0_chanx_out_17_;
wire [0:0] cbx_1__0__0_chanx_out_180_;
wire [0:0] cbx_1__0__0_chanx_out_181_;
wire [0:0] cbx_1__0__0_chanx_out_182_;
wire [0:0] cbx_1__0__0_chanx_out_183_;
wire [0:0] cbx_1__0__0_chanx_out_184_;
wire [0:0] cbx_1__0__0_chanx_out_185_;
wire [0:0] cbx_1__0__0_chanx_out_186_;
wire [0:0] cbx_1__0__0_chanx_out_187_;
wire [0:0] cbx_1__0__0_chanx_out_188_;
wire [0:0] cbx_1__0__0_chanx_out_189_;
wire [0:0] cbx_1__0__0_chanx_out_18_;
wire [0:0] cbx_1__0__0_chanx_out_190_;
wire [0:0] cbx_1__0__0_chanx_out_191_;
wire [0:0] cbx_1__0__0_chanx_out_192_;
wire [0:0] cbx_1__0__0_chanx_out_193_;
wire [0:0] cbx_1__0__0_chanx_out_194_;
wire [0:0] cbx_1__0__0_chanx_out_195_;
wire [0:0] cbx_1__0__0_chanx_out_196_;
wire [0:0] cbx_1__0__0_chanx_out_197_;
wire [0:0] cbx_1__0__0_chanx_out_198_;
wire [0:0] cbx_1__0__0_chanx_out_199_;
wire [0:0] cbx_1__0__0_chanx_out_19_;
wire [0:0] cbx_1__0__0_chanx_out_1_;
wire [0:0] cbx_1__0__0_chanx_out_20_;
wire [0:0] cbx_1__0__0_chanx_out_21_;
wire [0:0] cbx_1__0__0_chanx_out_22_;
wire [0:0] cbx_1__0__0_chanx_out_23_;
wire [0:0] cbx_1__0__0_chanx_out_24_;
wire [0:0] cbx_1__0__0_chanx_out_25_;
wire [0:0] cbx_1__0__0_chanx_out_26_;
wire [0:0] cbx_1__0__0_chanx_out_27_;
wire [0:0] cbx_1__0__0_chanx_out_28_;
wire [0:0] cbx_1__0__0_chanx_out_29_;
wire [0:0] cbx_1__0__0_chanx_out_2_;
wire [0:0] cbx_1__0__0_chanx_out_30_;
wire [0:0] cbx_1__0__0_chanx_out_31_;
wire [0:0] cbx_1__0__0_chanx_out_32_;
wire [0:0] cbx_1__0__0_chanx_out_33_;
wire [0:0] cbx_1__0__0_chanx_out_34_;
wire [0:0] cbx_1__0__0_chanx_out_35_;
wire [0:0] cbx_1__0__0_chanx_out_36_;
wire [0:0] cbx_1__0__0_chanx_out_37_;
wire [0:0] cbx_1__0__0_chanx_out_38_;
wire [0:0] cbx_1__0__0_chanx_out_39_;
wire [0:0] cbx_1__0__0_chanx_out_3_;
wire [0:0] cbx_1__0__0_chanx_out_40_;
wire [0:0] cbx_1__0__0_chanx_out_41_;
wire [0:0] cbx_1__0__0_chanx_out_42_;
wire [0:0] cbx_1__0__0_chanx_out_43_;
wire [0:0] cbx_1__0__0_chanx_out_44_;
wire [0:0] cbx_1__0__0_chanx_out_45_;
wire [0:0] cbx_1__0__0_chanx_out_46_;
wire [0:0] cbx_1__0__0_chanx_out_47_;
wire [0:0] cbx_1__0__0_chanx_out_48_;
wire [0:0] cbx_1__0__0_chanx_out_49_;
wire [0:0] cbx_1__0__0_chanx_out_4_;
wire [0:0] cbx_1__0__0_chanx_out_50_;
wire [0:0] cbx_1__0__0_chanx_out_51_;
wire [0:0] cbx_1__0__0_chanx_out_52_;
wire [0:0] cbx_1__0__0_chanx_out_53_;
wire [0:0] cbx_1__0__0_chanx_out_54_;
wire [0:0] cbx_1__0__0_chanx_out_55_;
wire [0:0] cbx_1__0__0_chanx_out_56_;
wire [0:0] cbx_1__0__0_chanx_out_57_;
wire [0:0] cbx_1__0__0_chanx_out_58_;
wire [0:0] cbx_1__0__0_chanx_out_59_;
wire [0:0] cbx_1__0__0_chanx_out_5_;
wire [0:0] cbx_1__0__0_chanx_out_60_;
wire [0:0] cbx_1__0__0_chanx_out_61_;
wire [0:0] cbx_1__0__0_chanx_out_62_;
wire [0:0] cbx_1__0__0_chanx_out_63_;
wire [0:0] cbx_1__0__0_chanx_out_64_;
wire [0:0] cbx_1__0__0_chanx_out_65_;
wire [0:0] cbx_1__0__0_chanx_out_66_;
wire [0:0] cbx_1__0__0_chanx_out_67_;
wire [0:0] cbx_1__0__0_chanx_out_68_;
wire [0:0] cbx_1__0__0_chanx_out_69_;
wire [0:0] cbx_1__0__0_chanx_out_6_;
wire [0:0] cbx_1__0__0_chanx_out_70_;
wire [0:0] cbx_1__0__0_chanx_out_71_;
wire [0:0] cbx_1__0__0_chanx_out_72_;
wire [0:0] cbx_1__0__0_chanx_out_73_;
wire [0:0] cbx_1__0__0_chanx_out_74_;
wire [0:0] cbx_1__0__0_chanx_out_75_;
wire [0:0] cbx_1__0__0_chanx_out_76_;
wire [0:0] cbx_1__0__0_chanx_out_77_;
wire [0:0] cbx_1__0__0_chanx_out_78_;
wire [0:0] cbx_1__0__0_chanx_out_79_;
wire [0:0] cbx_1__0__0_chanx_out_7_;
wire [0:0] cbx_1__0__0_chanx_out_80_;
wire [0:0] cbx_1__0__0_chanx_out_81_;
wire [0:0] cbx_1__0__0_chanx_out_82_;
wire [0:0] cbx_1__0__0_chanx_out_83_;
wire [0:0] cbx_1__0__0_chanx_out_84_;
wire [0:0] cbx_1__0__0_chanx_out_85_;
wire [0:0] cbx_1__0__0_chanx_out_86_;
wire [0:0] cbx_1__0__0_chanx_out_87_;
wire [0:0] cbx_1__0__0_chanx_out_88_;
wire [0:0] cbx_1__0__0_chanx_out_89_;
wire [0:0] cbx_1__0__0_chanx_out_8_;
wire [0:0] cbx_1__0__0_chanx_out_90_;
wire [0:0] cbx_1__0__0_chanx_out_91_;
wire [0:0] cbx_1__0__0_chanx_out_92_;
wire [0:0] cbx_1__0__0_chanx_out_93_;
wire [0:0] cbx_1__0__0_chanx_out_94_;
wire [0:0] cbx_1__0__0_chanx_out_95_;
wire [0:0] cbx_1__0__0_chanx_out_96_;
wire [0:0] cbx_1__0__0_chanx_out_97_;
wire [0:0] cbx_1__0__0_chanx_out_98_;
wire [0:0] cbx_1__0__0_chanx_out_99_;
wire [0:0] cbx_1__0__0_chanx_out_9_;
wire [0:0] cbx_1__0__0_top_grid_pin_20_;
wire [0:0] cbx_1__0__0_top_grid_pin_21_;
wire [0:0] cbx_1__0__0_top_grid_pin_22_;
wire [0:0] cbx_1__0__0_top_grid_pin_23_;
wire [0:0] cbx_1__0__0_top_grid_pin_24_;
wire [0:0] cbx_1__0__0_top_grid_pin_25_;
wire [0:0] cbx_1__0__0_top_grid_pin_26_;
wire [0:0] cbx_1__0__0_top_grid_pin_27_;
wire [0:0] cbx_1__0__0_top_grid_pin_28_;
wire [0:0] cbx_1__0__0_top_grid_pin_29_;
wire [0:0] cbx_1__0__0_top_grid_pin_30_;
wire [0:0] cbx_1__0__0_top_grid_pin_31_;
wire [0:0] cbx_1__0__0_top_grid_pin_32_;
wire [0:0] cbx_1__0__0_top_grid_pin_33_;
wire [0:0] cbx_1__0__0_top_grid_pin_34_;
wire [0:0] cbx_1__0__0_top_grid_pin_35_;
wire [0:0] cbx_1__0__0_top_grid_pin_36_;
wire [0:0] cbx_1__0__0_top_grid_pin_37_;
wire [0:0] cbx_1__0__0_top_grid_pin_38_;
wire [0:0] cbx_1__0__0_top_grid_pin_39_;
wire [0:0] cbx_1__0__1_bottom_grid_pin_0_;
wire [0:0] cbx_1__0__1_ccff_tail;
wire [0:0] cbx_1__0__1_chanx_out_0_;
wire [0:0] cbx_1__0__1_chanx_out_100_;
wire [0:0] cbx_1__0__1_chanx_out_101_;
wire [0:0] cbx_1__0__1_chanx_out_102_;
wire [0:0] cbx_1__0__1_chanx_out_103_;
wire [0:0] cbx_1__0__1_chanx_out_104_;
wire [0:0] cbx_1__0__1_chanx_out_105_;
wire [0:0] cbx_1__0__1_chanx_out_106_;
wire [0:0] cbx_1__0__1_chanx_out_107_;
wire [0:0] cbx_1__0__1_chanx_out_108_;
wire [0:0] cbx_1__0__1_chanx_out_109_;
wire [0:0] cbx_1__0__1_chanx_out_10_;
wire [0:0] cbx_1__0__1_chanx_out_110_;
wire [0:0] cbx_1__0__1_chanx_out_111_;
wire [0:0] cbx_1__0__1_chanx_out_112_;
wire [0:0] cbx_1__0__1_chanx_out_113_;
wire [0:0] cbx_1__0__1_chanx_out_114_;
wire [0:0] cbx_1__0__1_chanx_out_115_;
wire [0:0] cbx_1__0__1_chanx_out_116_;
wire [0:0] cbx_1__0__1_chanx_out_117_;
wire [0:0] cbx_1__0__1_chanx_out_118_;
wire [0:0] cbx_1__0__1_chanx_out_119_;
wire [0:0] cbx_1__0__1_chanx_out_11_;
wire [0:0] cbx_1__0__1_chanx_out_120_;
wire [0:0] cbx_1__0__1_chanx_out_121_;
wire [0:0] cbx_1__0__1_chanx_out_122_;
wire [0:0] cbx_1__0__1_chanx_out_123_;
wire [0:0] cbx_1__0__1_chanx_out_124_;
wire [0:0] cbx_1__0__1_chanx_out_125_;
wire [0:0] cbx_1__0__1_chanx_out_126_;
wire [0:0] cbx_1__0__1_chanx_out_127_;
wire [0:0] cbx_1__0__1_chanx_out_128_;
wire [0:0] cbx_1__0__1_chanx_out_129_;
wire [0:0] cbx_1__0__1_chanx_out_12_;
wire [0:0] cbx_1__0__1_chanx_out_130_;
wire [0:0] cbx_1__0__1_chanx_out_131_;
wire [0:0] cbx_1__0__1_chanx_out_132_;
wire [0:0] cbx_1__0__1_chanx_out_133_;
wire [0:0] cbx_1__0__1_chanx_out_134_;
wire [0:0] cbx_1__0__1_chanx_out_135_;
wire [0:0] cbx_1__0__1_chanx_out_136_;
wire [0:0] cbx_1__0__1_chanx_out_137_;
wire [0:0] cbx_1__0__1_chanx_out_138_;
wire [0:0] cbx_1__0__1_chanx_out_139_;
wire [0:0] cbx_1__0__1_chanx_out_13_;
wire [0:0] cbx_1__0__1_chanx_out_140_;
wire [0:0] cbx_1__0__1_chanx_out_141_;
wire [0:0] cbx_1__0__1_chanx_out_142_;
wire [0:0] cbx_1__0__1_chanx_out_143_;
wire [0:0] cbx_1__0__1_chanx_out_144_;
wire [0:0] cbx_1__0__1_chanx_out_145_;
wire [0:0] cbx_1__0__1_chanx_out_146_;
wire [0:0] cbx_1__0__1_chanx_out_147_;
wire [0:0] cbx_1__0__1_chanx_out_148_;
wire [0:0] cbx_1__0__1_chanx_out_149_;
wire [0:0] cbx_1__0__1_chanx_out_14_;
wire [0:0] cbx_1__0__1_chanx_out_150_;
wire [0:0] cbx_1__0__1_chanx_out_151_;
wire [0:0] cbx_1__0__1_chanx_out_152_;
wire [0:0] cbx_1__0__1_chanx_out_153_;
wire [0:0] cbx_1__0__1_chanx_out_154_;
wire [0:0] cbx_1__0__1_chanx_out_155_;
wire [0:0] cbx_1__0__1_chanx_out_156_;
wire [0:0] cbx_1__0__1_chanx_out_157_;
wire [0:0] cbx_1__0__1_chanx_out_158_;
wire [0:0] cbx_1__0__1_chanx_out_159_;
wire [0:0] cbx_1__0__1_chanx_out_15_;
wire [0:0] cbx_1__0__1_chanx_out_160_;
wire [0:0] cbx_1__0__1_chanx_out_161_;
wire [0:0] cbx_1__0__1_chanx_out_162_;
wire [0:0] cbx_1__0__1_chanx_out_163_;
wire [0:0] cbx_1__0__1_chanx_out_164_;
wire [0:0] cbx_1__0__1_chanx_out_165_;
wire [0:0] cbx_1__0__1_chanx_out_166_;
wire [0:0] cbx_1__0__1_chanx_out_167_;
wire [0:0] cbx_1__0__1_chanx_out_168_;
wire [0:0] cbx_1__0__1_chanx_out_169_;
wire [0:0] cbx_1__0__1_chanx_out_16_;
wire [0:0] cbx_1__0__1_chanx_out_170_;
wire [0:0] cbx_1__0__1_chanx_out_171_;
wire [0:0] cbx_1__0__1_chanx_out_172_;
wire [0:0] cbx_1__0__1_chanx_out_173_;
wire [0:0] cbx_1__0__1_chanx_out_174_;
wire [0:0] cbx_1__0__1_chanx_out_175_;
wire [0:0] cbx_1__0__1_chanx_out_176_;
wire [0:0] cbx_1__0__1_chanx_out_177_;
wire [0:0] cbx_1__0__1_chanx_out_178_;
wire [0:0] cbx_1__0__1_chanx_out_179_;
wire [0:0] cbx_1__0__1_chanx_out_17_;
wire [0:0] cbx_1__0__1_chanx_out_180_;
wire [0:0] cbx_1__0__1_chanx_out_181_;
wire [0:0] cbx_1__0__1_chanx_out_182_;
wire [0:0] cbx_1__0__1_chanx_out_183_;
wire [0:0] cbx_1__0__1_chanx_out_184_;
wire [0:0] cbx_1__0__1_chanx_out_185_;
wire [0:0] cbx_1__0__1_chanx_out_186_;
wire [0:0] cbx_1__0__1_chanx_out_187_;
wire [0:0] cbx_1__0__1_chanx_out_188_;
wire [0:0] cbx_1__0__1_chanx_out_189_;
wire [0:0] cbx_1__0__1_chanx_out_18_;
wire [0:0] cbx_1__0__1_chanx_out_190_;
wire [0:0] cbx_1__0__1_chanx_out_191_;
wire [0:0] cbx_1__0__1_chanx_out_192_;
wire [0:0] cbx_1__0__1_chanx_out_193_;
wire [0:0] cbx_1__0__1_chanx_out_194_;
wire [0:0] cbx_1__0__1_chanx_out_195_;
wire [0:0] cbx_1__0__1_chanx_out_196_;
wire [0:0] cbx_1__0__1_chanx_out_197_;
wire [0:0] cbx_1__0__1_chanx_out_198_;
wire [0:0] cbx_1__0__1_chanx_out_199_;
wire [0:0] cbx_1__0__1_chanx_out_19_;
wire [0:0] cbx_1__0__1_chanx_out_1_;
wire [0:0] cbx_1__0__1_chanx_out_20_;
wire [0:0] cbx_1__0__1_chanx_out_21_;
wire [0:0] cbx_1__0__1_chanx_out_22_;
wire [0:0] cbx_1__0__1_chanx_out_23_;
wire [0:0] cbx_1__0__1_chanx_out_24_;
wire [0:0] cbx_1__0__1_chanx_out_25_;
wire [0:0] cbx_1__0__1_chanx_out_26_;
wire [0:0] cbx_1__0__1_chanx_out_27_;
wire [0:0] cbx_1__0__1_chanx_out_28_;
wire [0:0] cbx_1__0__1_chanx_out_29_;
wire [0:0] cbx_1__0__1_chanx_out_2_;
wire [0:0] cbx_1__0__1_chanx_out_30_;
wire [0:0] cbx_1__0__1_chanx_out_31_;
wire [0:0] cbx_1__0__1_chanx_out_32_;
wire [0:0] cbx_1__0__1_chanx_out_33_;
wire [0:0] cbx_1__0__1_chanx_out_34_;
wire [0:0] cbx_1__0__1_chanx_out_35_;
wire [0:0] cbx_1__0__1_chanx_out_36_;
wire [0:0] cbx_1__0__1_chanx_out_37_;
wire [0:0] cbx_1__0__1_chanx_out_38_;
wire [0:0] cbx_1__0__1_chanx_out_39_;
wire [0:0] cbx_1__0__1_chanx_out_3_;
wire [0:0] cbx_1__0__1_chanx_out_40_;
wire [0:0] cbx_1__0__1_chanx_out_41_;
wire [0:0] cbx_1__0__1_chanx_out_42_;
wire [0:0] cbx_1__0__1_chanx_out_43_;
wire [0:0] cbx_1__0__1_chanx_out_44_;
wire [0:0] cbx_1__0__1_chanx_out_45_;
wire [0:0] cbx_1__0__1_chanx_out_46_;
wire [0:0] cbx_1__0__1_chanx_out_47_;
wire [0:0] cbx_1__0__1_chanx_out_48_;
wire [0:0] cbx_1__0__1_chanx_out_49_;
wire [0:0] cbx_1__0__1_chanx_out_4_;
wire [0:0] cbx_1__0__1_chanx_out_50_;
wire [0:0] cbx_1__0__1_chanx_out_51_;
wire [0:0] cbx_1__0__1_chanx_out_52_;
wire [0:0] cbx_1__0__1_chanx_out_53_;
wire [0:0] cbx_1__0__1_chanx_out_54_;
wire [0:0] cbx_1__0__1_chanx_out_55_;
wire [0:0] cbx_1__0__1_chanx_out_56_;
wire [0:0] cbx_1__0__1_chanx_out_57_;
wire [0:0] cbx_1__0__1_chanx_out_58_;
wire [0:0] cbx_1__0__1_chanx_out_59_;
wire [0:0] cbx_1__0__1_chanx_out_5_;
wire [0:0] cbx_1__0__1_chanx_out_60_;
wire [0:0] cbx_1__0__1_chanx_out_61_;
wire [0:0] cbx_1__0__1_chanx_out_62_;
wire [0:0] cbx_1__0__1_chanx_out_63_;
wire [0:0] cbx_1__0__1_chanx_out_64_;
wire [0:0] cbx_1__0__1_chanx_out_65_;
wire [0:0] cbx_1__0__1_chanx_out_66_;
wire [0:0] cbx_1__0__1_chanx_out_67_;
wire [0:0] cbx_1__0__1_chanx_out_68_;
wire [0:0] cbx_1__0__1_chanx_out_69_;
wire [0:0] cbx_1__0__1_chanx_out_6_;
wire [0:0] cbx_1__0__1_chanx_out_70_;
wire [0:0] cbx_1__0__1_chanx_out_71_;
wire [0:0] cbx_1__0__1_chanx_out_72_;
wire [0:0] cbx_1__0__1_chanx_out_73_;
wire [0:0] cbx_1__0__1_chanx_out_74_;
wire [0:0] cbx_1__0__1_chanx_out_75_;
wire [0:0] cbx_1__0__1_chanx_out_76_;
wire [0:0] cbx_1__0__1_chanx_out_77_;
wire [0:0] cbx_1__0__1_chanx_out_78_;
wire [0:0] cbx_1__0__1_chanx_out_79_;
wire [0:0] cbx_1__0__1_chanx_out_7_;
wire [0:0] cbx_1__0__1_chanx_out_80_;
wire [0:0] cbx_1__0__1_chanx_out_81_;
wire [0:0] cbx_1__0__1_chanx_out_82_;
wire [0:0] cbx_1__0__1_chanx_out_83_;
wire [0:0] cbx_1__0__1_chanx_out_84_;
wire [0:0] cbx_1__0__1_chanx_out_85_;
wire [0:0] cbx_1__0__1_chanx_out_86_;
wire [0:0] cbx_1__0__1_chanx_out_87_;
wire [0:0] cbx_1__0__1_chanx_out_88_;
wire [0:0] cbx_1__0__1_chanx_out_89_;
wire [0:0] cbx_1__0__1_chanx_out_8_;
wire [0:0] cbx_1__0__1_chanx_out_90_;
wire [0:0] cbx_1__0__1_chanx_out_91_;
wire [0:0] cbx_1__0__1_chanx_out_92_;
wire [0:0] cbx_1__0__1_chanx_out_93_;
wire [0:0] cbx_1__0__1_chanx_out_94_;
wire [0:0] cbx_1__0__1_chanx_out_95_;
wire [0:0] cbx_1__0__1_chanx_out_96_;
wire [0:0] cbx_1__0__1_chanx_out_97_;
wire [0:0] cbx_1__0__1_chanx_out_98_;
wire [0:0] cbx_1__0__1_chanx_out_99_;
wire [0:0] cbx_1__0__1_chanx_out_9_;
wire [0:0] cbx_1__0__1_top_grid_pin_20_;
wire [0:0] cbx_1__0__1_top_grid_pin_21_;
wire [0:0] cbx_1__0__1_top_grid_pin_22_;
wire [0:0] cbx_1__0__1_top_grid_pin_23_;
wire [0:0] cbx_1__0__1_top_grid_pin_24_;
wire [0:0] cbx_1__0__1_top_grid_pin_25_;
wire [0:0] cbx_1__0__1_top_grid_pin_26_;
wire [0:0] cbx_1__0__1_top_grid_pin_27_;
wire [0:0] cbx_1__0__1_top_grid_pin_28_;
wire [0:0] cbx_1__0__1_top_grid_pin_29_;
wire [0:0] cbx_1__0__1_top_grid_pin_30_;
wire [0:0] cbx_1__0__1_top_grid_pin_31_;
wire [0:0] cbx_1__0__1_top_grid_pin_32_;
wire [0:0] cbx_1__0__1_top_grid_pin_33_;
wire [0:0] cbx_1__0__1_top_grid_pin_34_;
wire [0:0] cbx_1__0__1_top_grid_pin_35_;
wire [0:0] cbx_1__0__1_top_grid_pin_36_;
wire [0:0] cbx_1__0__1_top_grid_pin_37_;
wire [0:0] cbx_1__0__1_top_grid_pin_38_;
wire [0:0] cbx_1__0__1_top_grid_pin_39_;
wire [0:0] cbx_1__1__0_bottom_grid_pin_42_;
wire [0:0] cbx_1__1__0_bottom_grid_pin_43_;
wire [0:0] cbx_1__1__0_bottom_grid_pin_69_;
wire [0:0] cbx_1__1__0_ccff_tail;
wire [0:0] cbx_1__1__0_chanx_out_0_;
wire [0:0] cbx_1__1__0_chanx_out_100_;
wire [0:0] cbx_1__1__0_chanx_out_101_;
wire [0:0] cbx_1__1__0_chanx_out_102_;
wire [0:0] cbx_1__1__0_chanx_out_103_;
wire [0:0] cbx_1__1__0_chanx_out_104_;
wire [0:0] cbx_1__1__0_chanx_out_105_;
wire [0:0] cbx_1__1__0_chanx_out_106_;
wire [0:0] cbx_1__1__0_chanx_out_107_;
wire [0:0] cbx_1__1__0_chanx_out_108_;
wire [0:0] cbx_1__1__0_chanx_out_109_;
wire [0:0] cbx_1__1__0_chanx_out_10_;
wire [0:0] cbx_1__1__0_chanx_out_110_;
wire [0:0] cbx_1__1__0_chanx_out_111_;
wire [0:0] cbx_1__1__0_chanx_out_112_;
wire [0:0] cbx_1__1__0_chanx_out_113_;
wire [0:0] cbx_1__1__0_chanx_out_114_;
wire [0:0] cbx_1__1__0_chanx_out_115_;
wire [0:0] cbx_1__1__0_chanx_out_116_;
wire [0:0] cbx_1__1__0_chanx_out_117_;
wire [0:0] cbx_1__1__0_chanx_out_118_;
wire [0:0] cbx_1__1__0_chanx_out_119_;
wire [0:0] cbx_1__1__0_chanx_out_11_;
wire [0:0] cbx_1__1__0_chanx_out_120_;
wire [0:0] cbx_1__1__0_chanx_out_121_;
wire [0:0] cbx_1__1__0_chanx_out_122_;
wire [0:0] cbx_1__1__0_chanx_out_123_;
wire [0:0] cbx_1__1__0_chanx_out_124_;
wire [0:0] cbx_1__1__0_chanx_out_125_;
wire [0:0] cbx_1__1__0_chanx_out_126_;
wire [0:0] cbx_1__1__0_chanx_out_127_;
wire [0:0] cbx_1__1__0_chanx_out_128_;
wire [0:0] cbx_1__1__0_chanx_out_129_;
wire [0:0] cbx_1__1__0_chanx_out_12_;
wire [0:0] cbx_1__1__0_chanx_out_130_;
wire [0:0] cbx_1__1__0_chanx_out_131_;
wire [0:0] cbx_1__1__0_chanx_out_132_;
wire [0:0] cbx_1__1__0_chanx_out_133_;
wire [0:0] cbx_1__1__0_chanx_out_134_;
wire [0:0] cbx_1__1__0_chanx_out_135_;
wire [0:0] cbx_1__1__0_chanx_out_136_;
wire [0:0] cbx_1__1__0_chanx_out_137_;
wire [0:0] cbx_1__1__0_chanx_out_138_;
wire [0:0] cbx_1__1__0_chanx_out_139_;
wire [0:0] cbx_1__1__0_chanx_out_13_;
wire [0:0] cbx_1__1__0_chanx_out_140_;
wire [0:0] cbx_1__1__0_chanx_out_141_;
wire [0:0] cbx_1__1__0_chanx_out_142_;
wire [0:0] cbx_1__1__0_chanx_out_143_;
wire [0:0] cbx_1__1__0_chanx_out_144_;
wire [0:0] cbx_1__1__0_chanx_out_145_;
wire [0:0] cbx_1__1__0_chanx_out_146_;
wire [0:0] cbx_1__1__0_chanx_out_147_;
wire [0:0] cbx_1__1__0_chanx_out_148_;
wire [0:0] cbx_1__1__0_chanx_out_149_;
wire [0:0] cbx_1__1__0_chanx_out_14_;
wire [0:0] cbx_1__1__0_chanx_out_150_;
wire [0:0] cbx_1__1__0_chanx_out_151_;
wire [0:0] cbx_1__1__0_chanx_out_152_;
wire [0:0] cbx_1__1__0_chanx_out_153_;
wire [0:0] cbx_1__1__0_chanx_out_154_;
wire [0:0] cbx_1__1__0_chanx_out_155_;
wire [0:0] cbx_1__1__0_chanx_out_156_;
wire [0:0] cbx_1__1__0_chanx_out_157_;
wire [0:0] cbx_1__1__0_chanx_out_158_;
wire [0:0] cbx_1__1__0_chanx_out_159_;
wire [0:0] cbx_1__1__0_chanx_out_15_;
wire [0:0] cbx_1__1__0_chanx_out_160_;
wire [0:0] cbx_1__1__0_chanx_out_161_;
wire [0:0] cbx_1__1__0_chanx_out_162_;
wire [0:0] cbx_1__1__0_chanx_out_163_;
wire [0:0] cbx_1__1__0_chanx_out_164_;
wire [0:0] cbx_1__1__0_chanx_out_165_;
wire [0:0] cbx_1__1__0_chanx_out_166_;
wire [0:0] cbx_1__1__0_chanx_out_167_;
wire [0:0] cbx_1__1__0_chanx_out_168_;
wire [0:0] cbx_1__1__0_chanx_out_169_;
wire [0:0] cbx_1__1__0_chanx_out_16_;
wire [0:0] cbx_1__1__0_chanx_out_170_;
wire [0:0] cbx_1__1__0_chanx_out_171_;
wire [0:0] cbx_1__1__0_chanx_out_172_;
wire [0:0] cbx_1__1__0_chanx_out_173_;
wire [0:0] cbx_1__1__0_chanx_out_174_;
wire [0:0] cbx_1__1__0_chanx_out_175_;
wire [0:0] cbx_1__1__0_chanx_out_176_;
wire [0:0] cbx_1__1__0_chanx_out_177_;
wire [0:0] cbx_1__1__0_chanx_out_178_;
wire [0:0] cbx_1__1__0_chanx_out_179_;
wire [0:0] cbx_1__1__0_chanx_out_17_;
wire [0:0] cbx_1__1__0_chanx_out_180_;
wire [0:0] cbx_1__1__0_chanx_out_181_;
wire [0:0] cbx_1__1__0_chanx_out_182_;
wire [0:0] cbx_1__1__0_chanx_out_183_;
wire [0:0] cbx_1__1__0_chanx_out_184_;
wire [0:0] cbx_1__1__0_chanx_out_185_;
wire [0:0] cbx_1__1__0_chanx_out_186_;
wire [0:0] cbx_1__1__0_chanx_out_187_;
wire [0:0] cbx_1__1__0_chanx_out_188_;
wire [0:0] cbx_1__1__0_chanx_out_189_;
wire [0:0] cbx_1__1__0_chanx_out_18_;
wire [0:0] cbx_1__1__0_chanx_out_190_;
wire [0:0] cbx_1__1__0_chanx_out_191_;
wire [0:0] cbx_1__1__0_chanx_out_192_;
wire [0:0] cbx_1__1__0_chanx_out_193_;
wire [0:0] cbx_1__1__0_chanx_out_194_;
wire [0:0] cbx_1__1__0_chanx_out_195_;
wire [0:0] cbx_1__1__0_chanx_out_196_;
wire [0:0] cbx_1__1__0_chanx_out_197_;
wire [0:0] cbx_1__1__0_chanx_out_198_;
wire [0:0] cbx_1__1__0_chanx_out_199_;
wire [0:0] cbx_1__1__0_chanx_out_19_;
wire [0:0] cbx_1__1__0_chanx_out_1_;
wire [0:0] cbx_1__1__0_chanx_out_20_;
wire [0:0] cbx_1__1__0_chanx_out_21_;
wire [0:0] cbx_1__1__0_chanx_out_22_;
wire [0:0] cbx_1__1__0_chanx_out_23_;
wire [0:0] cbx_1__1__0_chanx_out_24_;
wire [0:0] cbx_1__1__0_chanx_out_25_;
wire [0:0] cbx_1__1__0_chanx_out_26_;
wire [0:0] cbx_1__1__0_chanx_out_27_;
wire [0:0] cbx_1__1__0_chanx_out_28_;
wire [0:0] cbx_1__1__0_chanx_out_29_;
wire [0:0] cbx_1__1__0_chanx_out_2_;
wire [0:0] cbx_1__1__0_chanx_out_30_;
wire [0:0] cbx_1__1__0_chanx_out_31_;
wire [0:0] cbx_1__1__0_chanx_out_32_;
wire [0:0] cbx_1__1__0_chanx_out_33_;
wire [0:0] cbx_1__1__0_chanx_out_34_;
wire [0:0] cbx_1__1__0_chanx_out_35_;
wire [0:0] cbx_1__1__0_chanx_out_36_;
wire [0:0] cbx_1__1__0_chanx_out_37_;
wire [0:0] cbx_1__1__0_chanx_out_38_;
wire [0:0] cbx_1__1__0_chanx_out_39_;
wire [0:0] cbx_1__1__0_chanx_out_3_;
wire [0:0] cbx_1__1__0_chanx_out_40_;
wire [0:0] cbx_1__1__0_chanx_out_41_;
wire [0:0] cbx_1__1__0_chanx_out_42_;
wire [0:0] cbx_1__1__0_chanx_out_43_;
wire [0:0] cbx_1__1__0_chanx_out_44_;
wire [0:0] cbx_1__1__0_chanx_out_45_;
wire [0:0] cbx_1__1__0_chanx_out_46_;
wire [0:0] cbx_1__1__0_chanx_out_47_;
wire [0:0] cbx_1__1__0_chanx_out_48_;
wire [0:0] cbx_1__1__0_chanx_out_49_;
wire [0:0] cbx_1__1__0_chanx_out_4_;
wire [0:0] cbx_1__1__0_chanx_out_50_;
wire [0:0] cbx_1__1__0_chanx_out_51_;
wire [0:0] cbx_1__1__0_chanx_out_52_;
wire [0:0] cbx_1__1__0_chanx_out_53_;
wire [0:0] cbx_1__1__0_chanx_out_54_;
wire [0:0] cbx_1__1__0_chanx_out_55_;
wire [0:0] cbx_1__1__0_chanx_out_56_;
wire [0:0] cbx_1__1__0_chanx_out_57_;
wire [0:0] cbx_1__1__0_chanx_out_58_;
wire [0:0] cbx_1__1__0_chanx_out_59_;
wire [0:0] cbx_1__1__0_chanx_out_5_;
wire [0:0] cbx_1__1__0_chanx_out_60_;
wire [0:0] cbx_1__1__0_chanx_out_61_;
wire [0:0] cbx_1__1__0_chanx_out_62_;
wire [0:0] cbx_1__1__0_chanx_out_63_;
wire [0:0] cbx_1__1__0_chanx_out_64_;
wire [0:0] cbx_1__1__0_chanx_out_65_;
wire [0:0] cbx_1__1__0_chanx_out_66_;
wire [0:0] cbx_1__1__0_chanx_out_67_;
wire [0:0] cbx_1__1__0_chanx_out_68_;
wire [0:0] cbx_1__1__0_chanx_out_69_;
wire [0:0] cbx_1__1__0_chanx_out_6_;
wire [0:0] cbx_1__1__0_chanx_out_70_;
wire [0:0] cbx_1__1__0_chanx_out_71_;
wire [0:0] cbx_1__1__0_chanx_out_72_;
wire [0:0] cbx_1__1__0_chanx_out_73_;
wire [0:0] cbx_1__1__0_chanx_out_74_;
wire [0:0] cbx_1__1__0_chanx_out_75_;
wire [0:0] cbx_1__1__0_chanx_out_76_;
wire [0:0] cbx_1__1__0_chanx_out_77_;
wire [0:0] cbx_1__1__0_chanx_out_78_;
wire [0:0] cbx_1__1__0_chanx_out_79_;
wire [0:0] cbx_1__1__0_chanx_out_7_;
wire [0:0] cbx_1__1__0_chanx_out_80_;
wire [0:0] cbx_1__1__0_chanx_out_81_;
wire [0:0] cbx_1__1__0_chanx_out_82_;
wire [0:0] cbx_1__1__0_chanx_out_83_;
wire [0:0] cbx_1__1__0_chanx_out_84_;
wire [0:0] cbx_1__1__0_chanx_out_85_;
wire [0:0] cbx_1__1__0_chanx_out_86_;
wire [0:0] cbx_1__1__0_chanx_out_87_;
wire [0:0] cbx_1__1__0_chanx_out_88_;
wire [0:0] cbx_1__1__0_chanx_out_89_;
wire [0:0] cbx_1__1__0_chanx_out_8_;
wire [0:0] cbx_1__1__0_chanx_out_90_;
wire [0:0] cbx_1__1__0_chanx_out_91_;
wire [0:0] cbx_1__1__0_chanx_out_92_;
wire [0:0] cbx_1__1__0_chanx_out_93_;
wire [0:0] cbx_1__1__0_chanx_out_94_;
wire [0:0] cbx_1__1__0_chanx_out_95_;
wire [0:0] cbx_1__1__0_chanx_out_96_;
wire [0:0] cbx_1__1__0_chanx_out_97_;
wire [0:0] cbx_1__1__0_chanx_out_98_;
wire [0:0] cbx_1__1__0_chanx_out_99_;
wire [0:0] cbx_1__1__0_chanx_out_9_;
wire [0:0] cbx_1__1__0_top_grid_pin_20_;
wire [0:0] cbx_1__1__0_top_grid_pin_21_;
wire [0:0] cbx_1__1__0_top_grid_pin_22_;
wire [0:0] cbx_1__1__0_top_grid_pin_23_;
wire [0:0] cbx_1__1__0_top_grid_pin_24_;
wire [0:0] cbx_1__1__0_top_grid_pin_25_;
wire [0:0] cbx_1__1__0_top_grid_pin_26_;
wire [0:0] cbx_1__1__0_top_grid_pin_27_;
wire [0:0] cbx_1__1__0_top_grid_pin_28_;
wire [0:0] cbx_1__1__0_top_grid_pin_29_;
wire [0:0] cbx_1__1__0_top_grid_pin_30_;
wire [0:0] cbx_1__1__0_top_grid_pin_31_;
wire [0:0] cbx_1__1__0_top_grid_pin_32_;
wire [0:0] cbx_1__1__0_top_grid_pin_33_;
wire [0:0] cbx_1__1__0_top_grid_pin_34_;
wire [0:0] cbx_1__1__0_top_grid_pin_35_;
wire [0:0] cbx_1__1__0_top_grid_pin_36_;
wire [0:0] cbx_1__1__0_top_grid_pin_37_;
wire [0:0] cbx_1__1__0_top_grid_pin_38_;
wire [0:0] cbx_1__1__0_top_grid_pin_39_;
wire [0:0] cbx_1__1__1_bottom_grid_pin_42_;
wire [0:0] cbx_1__1__1_bottom_grid_pin_43_;
wire [0:0] cbx_1__1__1_bottom_grid_pin_69_;
wire [0:0] cbx_1__1__1_ccff_tail;
wire [0:0] cbx_1__1__1_chanx_out_0_;
wire [0:0] cbx_1__1__1_chanx_out_100_;
wire [0:0] cbx_1__1__1_chanx_out_101_;
wire [0:0] cbx_1__1__1_chanx_out_102_;
wire [0:0] cbx_1__1__1_chanx_out_103_;
wire [0:0] cbx_1__1__1_chanx_out_104_;
wire [0:0] cbx_1__1__1_chanx_out_105_;
wire [0:0] cbx_1__1__1_chanx_out_106_;
wire [0:0] cbx_1__1__1_chanx_out_107_;
wire [0:0] cbx_1__1__1_chanx_out_108_;
wire [0:0] cbx_1__1__1_chanx_out_109_;
wire [0:0] cbx_1__1__1_chanx_out_10_;
wire [0:0] cbx_1__1__1_chanx_out_110_;
wire [0:0] cbx_1__1__1_chanx_out_111_;
wire [0:0] cbx_1__1__1_chanx_out_112_;
wire [0:0] cbx_1__1__1_chanx_out_113_;
wire [0:0] cbx_1__1__1_chanx_out_114_;
wire [0:0] cbx_1__1__1_chanx_out_115_;
wire [0:0] cbx_1__1__1_chanx_out_116_;
wire [0:0] cbx_1__1__1_chanx_out_117_;
wire [0:0] cbx_1__1__1_chanx_out_118_;
wire [0:0] cbx_1__1__1_chanx_out_119_;
wire [0:0] cbx_1__1__1_chanx_out_11_;
wire [0:0] cbx_1__1__1_chanx_out_120_;
wire [0:0] cbx_1__1__1_chanx_out_121_;
wire [0:0] cbx_1__1__1_chanx_out_122_;
wire [0:0] cbx_1__1__1_chanx_out_123_;
wire [0:0] cbx_1__1__1_chanx_out_124_;
wire [0:0] cbx_1__1__1_chanx_out_125_;
wire [0:0] cbx_1__1__1_chanx_out_126_;
wire [0:0] cbx_1__1__1_chanx_out_127_;
wire [0:0] cbx_1__1__1_chanx_out_128_;
wire [0:0] cbx_1__1__1_chanx_out_129_;
wire [0:0] cbx_1__1__1_chanx_out_12_;
wire [0:0] cbx_1__1__1_chanx_out_130_;
wire [0:0] cbx_1__1__1_chanx_out_131_;
wire [0:0] cbx_1__1__1_chanx_out_132_;
wire [0:0] cbx_1__1__1_chanx_out_133_;
wire [0:0] cbx_1__1__1_chanx_out_134_;
wire [0:0] cbx_1__1__1_chanx_out_135_;
wire [0:0] cbx_1__1__1_chanx_out_136_;
wire [0:0] cbx_1__1__1_chanx_out_137_;
wire [0:0] cbx_1__1__1_chanx_out_138_;
wire [0:0] cbx_1__1__1_chanx_out_139_;
wire [0:0] cbx_1__1__1_chanx_out_13_;
wire [0:0] cbx_1__1__1_chanx_out_140_;
wire [0:0] cbx_1__1__1_chanx_out_141_;
wire [0:0] cbx_1__1__1_chanx_out_142_;
wire [0:0] cbx_1__1__1_chanx_out_143_;
wire [0:0] cbx_1__1__1_chanx_out_144_;
wire [0:0] cbx_1__1__1_chanx_out_145_;
wire [0:0] cbx_1__1__1_chanx_out_146_;
wire [0:0] cbx_1__1__1_chanx_out_147_;
wire [0:0] cbx_1__1__1_chanx_out_148_;
wire [0:0] cbx_1__1__1_chanx_out_149_;
wire [0:0] cbx_1__1__1_chanx_out_14_;
wire [0:0] cbx_1__1__1_chanx_out_150_;
wire [0:0] cbx_1__1__1_chanx_out_151_;
wire [0:0] cbx_1__1__1_chanx_out_152_;
wire [0:0] cbx_1__1__1_chanx_out_153_;
wire [0:0] cbx_1__1__1_chanx_out_154_;
wire [0:0] cbx_1__1__1_chanx_out_155_;
wire [0:0] cbx_1__1__1_chanx_out_156_;
wire [0:0] cbx_1__1__1_chanx_out_157_;
wire [0:0] cbx_1__1__1_chanx_out_158_;
wire [0:0] cbx_1__1__1_chanx_out_159_;
wire [0:0] cbx_1__1__1_chanx_out_15_;
wire [0:0] cbx_1__1__1_chanx_out_160_;
wire [0:0] cbx_1__1__1_chanx_out_161_;
wire [0:0] cbx_1__1__1_chanx_out_162_;
wire [0:0] cbx_1__1__1_chanx_out_163_;
wire [0:0] cbx_1__1__1_chanx_out_164_;
wire [0:0] cbx_1__1__1_chanx_out_165_;
wire [0:0] cbx_1__1__1_chanx_out_166_;
wire [0:0] cbx_1__1__1_chanx_out_167_;
wire [0:0] cbx_1__1__1_chanx_out_168_;
wire [0:0] cbx_1__1__1_chanx_out_169_;
wire [0:0] cbx_1__1__1_chanx_out_16_;
wire [0:0] cbx_1__1__1_chanx_out_170_;
wire [0:0] cbx_1__1__1_chanx_out_171_;
wire [0:0] cbx_1__1__1_chanx_out_172_;
wire [0:0] cbx_1__1__1_chanx_out_173_;
wire [0:0] cbx_1__1__1_chanx_out_174_;
wire [0:0] cbx_1__1__1_chanx_out_175_;
wire [0:0] cbx_1__1__1_chanx_out_176_;
wire [0:0] cbx_1__1__1_chanx_out_177_;
wire [0:0] cbx_1__1__1_chanx_out_178_;
wire [0:0] cbx_1__1__1_chanx_out_179_;
wire [0:0] cbx_1__1__1_chanx_out_17_;
wire [0:0] cbx_1__1__1_chanx_out_180_;
wire [0:0] cbx_1__1__1_chanx_out_181_;
wire [0:0] cbx_1__1__1_chanx_out_182_;
wire [0:0] cbx_1__1__1_chanx_out_183_;
wire [0:0] cbx_1__1__1_chanx_out_184_;
wire [0:0] cbx_1__1__1_chanx_out_185_;
wire [0:0] cbx_1__1__1_chanx_out_186_;
wire [0:0] cbx_1__1__1_chanx_out_187_;
wire [0:0] cbx_1__1__1_chanx_out_188_;
wire [0:0] cbx_1__1__1_chanx_out_189_;
wire [0:0] cbx_1__1__1_chanx_out_18_;
wire [0:0] cbx_1__1__1_chanx_out_190_;
wire [0:0] cbx_1__1__1_chanx_out_191_;
wire [0:0] cbx_1__1__1_chanx_out_192_;
wire [0:0] cbx_1__1__1_chanx_out_193_;
wire [0:0] cbx_1__1__1_chanx_out_194_;
wire [0:0] cbx_1__1__1_chanx_out_195_;
wire [0:0] cbx_1__1__1_chanx_out_196_;
wire [0:0] cbx_1__1__1_chanx_out_197_;
wire [0:0] cbx_1__1__1_chanx_out_198_;
wire [0:0] cbx_1__1__1_chanx_out_199_;
wire [0:0] cbx_1__1__1_chanx_out_19_;
wire [0:0] cbx_1__1__1_chanx_out_1_;
wire [0:0] cbx_1__1__1_chanx_out_20_;
wire [0:0] cbx_1__1__1_chanx_out_21_;
wire [0:0] cbx_1__1__1_chanx_out_22_;
wire [0:0] cbx_1__1__1_chanx_out_23_;
wire [0:0] cbx_1__1__1_chanx_out_24_;
wire [0:0] cbx_1__1__1_chanx_out_25_;
wire [0:0] cbx_1__1__1_chanx_out_26_;
wire [0:0] cbx_1__1__1_chanx_out_27_;
wire [0:0] cbx_1__1__1_chanx_out_28_;
wire [0:0] cbx_1__1__1_chanx_out_29_;
wire [0:0] cbx_1__1__1_chanx_out_2_;
wire [0:0] cbx_1__1__1_chanx_out_30_;
wire [0:0] cbx_1__1__1_chanx_out_31_;
wire [0:0] cbx_1__1__1_chanx_out_32_;
wire [0:0] cbx_1__1__1_chanx_out_33_;
wire [0:0] cbx_1__1__1_chanx_out_34_;
wire [0:0] cbx_1__1__1_chanx_out_35_;
wire [0:0] cbx_1__1__1_chanx_out_36_;
wire [0:0] cbx_1__1__1_chanx_out_37_;
wire [0:0] cbx_1__1__1_chanx_out_38_;
wire [0:0] cbx_1__1__1_chanx_out_39_;
wire [0:0] cbx_1__1__1_chanx_out_3_;
wire [0:0] cbx_1__1__1_chanx_out_40_;
wire [0:0] cbx_1__1__1_chanx_out_41_;
wire [0:0] cbx_1__1__1_chanx_out_42_;
wire [0:0] cbx_1__1__1_chanx_out_43_;
wire [0:0] cbx_1__1__1_chanx_out_44_;
wire [0:0] cbx_1__1__1_chanx_out_45_;
wire [0:0] cbx_1__1__1_chanx_out_46_;
wire [0:0] cbx_1__1__1_chanx_out_47_;
wire [0:0] cbx_1__1__1_chanx_out_48_;
wire [0:0] cbx_1__1__1_chanx_out_49_;
wire [0:0] cbx_1__1__1_chanx_out_4_;
wire [0:0] cbx_1__1__1_chanx_out_50_;
wire [0:0] cbx_1__1__1_chanx_out_51_;
wire [0:0] cbx_1__1__1_chanx_out_52_;
wire [0:0] cbx_1__1__1_chanx_out_53_;
wire [0:0] cbx_1__1__1_chanx_out_54_;
wire [0:0] cbx_1__1__1_chanx_out_55_;
wire [0:0] cbx_1__1__1_chanx_out_56_;
wire [0:0] cbx_1__1__1_chanx_out_57_;
wire [0:0] cbx_1__1__1_chanx_out_58_;
wire [0:0] cbx_1__1__1_chanx_out_59_;
wire [0:0] cbx_1__1__1_chanx_out_5_;
wire [0:0] cbx_1__1__1_chanx_out_60_;
wire [0:0] cbx_1__1__1_chanx_out_61_;
wire [0:0] cbx_1__1__1_chanx_out_62_;
wire [0:0] cbx_1__1__1_chanx_out_63_;
wire [0:0] cbx_1__1__1_chanx_out_64_;
wire [0:0] cbx_1__1__1_chanx_out_65_;
wire [0:0] cbx_1__1__1_chanx_out_66_;
wire [0:0] cbx_1__1__1_chanx_out_67_;
wire [0:0] cbx_1__1__1_chanx_out_68_;
wire [0:0] cbx_1__1__1_chanx_out_69_;
wire [0:0] cbx_1__1__1_chanx_out_6_;
wire [0:0] cbx_1__1__1_chanx_out_70_;
wire [0:0] cbx_1__1__1_chanx_out_71_;
wire [0:0] cbx_1__1__1_chanx_out_72_;
wire [0:0] cbx_1__1__1_chanx_out_73_;
wire [0:0] cbx_1__1__1_chanx_out_74_;
wire [0:0] cbx_1__1__1_chanx_out_75_;
wire [0:0] cbx_1__1__1_chanx_out_76_;
wire [0:0] cbx_1__1__1_chanx_out_77_;
wire [0:0] cbx_1__1__1_chanx_out_78_;
wire [0:0] cbx_1__1__1_chanx_out_79_;
wire [0:0] cbx_1__1__1_chanx_out_7_;
wire [0:0] cbx_1__1__1_chanx_out_80_;
wire [0:0] cbx_1__1__1_chanx_out_81_;
wire [0:0] cbx_1__1__1_chanx_out_82_;
wire [0:0] cbx_1__1__1_chanx_out_83_;
wire [0:0] cbx_1__1__1_chanx_out_84_;
wire [0:0] cbx_1__1__1_chanx_out_85_;
wire [0:0] cbx_1__1__1_chanx_out_86_;
wire [0:0] cbx_1__1__1_chanx_out_87_;
wire [0:0] cbx_1__1__1_chanx_out_88_;
wire [0:0] cbx_1__1__1_chanx_out_89_;
wire [0:0] cbx_1__1__1_chanx_out_8_;
wire [0:0] cbx_1__1__1_chanx_out_90_;
wire [0:0] cbx_1__1__1_chanx_out_91_;
wire [0:0] cbx_1__1__1_chanx_out_92_;
wire [0:0] cbx_1__1__1_chanx_out_93_;
wire [0:0] cbx_1__1__1_chanx_out_94_;
wire [0:0] cbx_1__1__1_chanx_out_95_;
wire [0:0] cbx_1__1__1_chanx_out_96_;
wire [0:0] cbx_1__1__1_chanx_out_97_;
wire [0:0] cbx_1__1__1_chanx_out_98_;
wire [0:0] cbx_1__1__1_chanx_out_99_;
wire [0:0] cbx_1__1__1_chanx_out_9_;
wire [0:0] cbx_1__1__1_top_grid_pin_20_;
wire [0:0] cbx_1__1__1_top_grid_pin_21_;
wire [0:0] cbx_1__1__1_top_grid_pin_22_;
wire [0:0] cbx_1__1__1_top_grid_pin_23_;
wire [0:0] cbx_1__1__1_top_grid_pin_24_;
wire [0:0] cbx_1__1__1_top_grid_pin_25_;
wire [0:0] cbx_1__1__1_top_grid_pin_26_;
wire [0:0] cbx_1__1__1_top_grid_pin_27_;
wire [0:0] cbx_1__1__1_top_grid_pin_28_;
wire [0:0] cbx_1__1__1_top_grid_pin_29_;
wire [0:0] cbx_1__1__1_top_grid_pin_30_;
wire [0:0] cbx_1__1__1_top_grid_pin_31_;
wire [0:0] cbx_1__1__1_top_grid_pin_32_;
wire [0:0] cbx_1__1__1_top_grid_pin_33_;
wire [0:0] cbx_1__1__1_top_grid_pin_34_;
wire [0:0] cbx_1__1__1_top_grid_pin_35_;
wire [0:0] cbx_1__1__1_top_grid_pin_36_;
wire [0:0] cbx_1__1__1_top_grid_pin_37_;
wire [0:0] cbx_1__1__1_top_grid_pin_38_;
wire [0:0] cbx_1__1__1_top_grid_pin_39_;
wire [0:0] cbx_1__2__0_bottom_grid_pin_42_;
wire [0:0] cbx_1__2__0_bottom_grid_pin_43_;
wire [0:0] cbx_1__2__0_bottom_grid_pin_68_;
wire [0:0] cbx_1__2__0_ccff_tail;
wire [0:0] cbx_1__2__0_chanx_out_0_;
wire [0:0] cbx_1__2__0_chanx_out_100_;
wire [0:0] cbx_1__2__0_chanx_out_101_;
wire [0:0] cbx_1__2__0_chanx_out_102_;
wire [0:0] cbx_1__2__0_chanx_out_103_;
wire [0:0] cbx_1__2__0_chanx_out_104_;
wire [0:0] cbx_1__2__0_chanx_out_105_;
wire [0:0] cbx_1__2__0_chanx_out_106_;
wire [0:0] cbx_1__2__0_chanx_out_107_;
wire [0:0] cbx_1__2__0_chanx_out_108_;
wire [0:0] cbx_1__2__0_chanx_out_109_;
wire [0:0] cbx_1__2__0_chanx_out_10_;
wire [0:0] cbx_1__2__0_chanx_out_110_;
wire [0:0] cbx_1__2__0_chanx_out_111_;
wire [0:0] cbx_1__2__0_chanx_out_112_;
wire [0:0] cbx_1__2__0_chanx_out_113_;
wire [0:0] cbx_1__2__0_chanx_out_114_;
wire [0:0] cbx_1__2__0_chanx_out_115_;
wire [0:0] cbx_1__2__0_chanx_out_116_;
wire [0:0] cbx_1__2__0_chanx_out_117_;
wire [0:0] cbx_1__2__0_chanx_out_118_;
wire [0:0] cbx_1__2__0_chanx_out_119_;
wire [0:0] cbx_1__2__0_chanx_out_11_;
wire [0:0] cbx_1__2__0_chanx_out_120_;
wire [0:0] cbx_1__2__0_chanx_out_121_;
wire [0:0] cbx_1__2__0_chanx_out_122_;
wire [0:0] cbx_1__2__0_chanx_out_123_;
wire [0:0] cbx_1__2__0_chanx_out_124_;
wire [0:0] cbx_1__2__0_chanx_out_125_;
wire [0:0] cbx_1__2__0_chanx_out_126_;
wire [0:0] cbx_1__2__0_chanx_out_127_;
wire [0:0] cbx_1__2__0_chanx_out_128_;
wire [0:0] cbx_1__2__0_chanx_out_129_;
wire [0:0] cbx_1__2__0_chanx_out_12_;
wire [0:0] cbx_1__2__0_chanx_out_130_;
wire [0:0] cbx_1__2__0_chanx_out_131_;
wire [0:0] cbx_1__2__0_chanx_out_132_;
wire [0:0] cbx_1__2__0_chanx_out_133_;
wire [0:0] cbx_1__2__0_chanx_out_134_;
wire [0:0] cbx_1__2__0_chanx_out_135_;
wire [0:0] cbx_1__2__0_chanx_out_136_;
wire [0:0] cbx_1__2__0_chanx_out_137_;
wire [0:0] cbx_1__2__0_chanx_out_138_;
wire [0:0] cbx_1__2__0_chanx_out_139_;
wire [0:0] cbx_1__2__0_chanx_out_13_;
wire [0:0] cbx_1__2__0_chanx_out_140_;
wire [0:0] cbx_1__2__0_chanx_out_141_;
wire [0:0] cbx_1__2__0_chanx_out_142_;
wire [0:0] cbx_1__2__0_chanx_out_143_;
wire [0:0] cbx_1__2__0_chanx_out_144_;
wire [0:0] cbx_1__2__0_chanx_out_145_;
wire [0:0] cbx_1__2__0_chanx_out_146_;
wire [0:0] cbx_1__2__0_chanx_out_147_;
wire [0:0] cbx_1__2__0_chanx_out_148_;
wire [0:0] cbx_1__2__0_chanx_out_149_;
wire [0:0] cbx_1__2__0_chanx_out_14_;
wire [0:0] cbx_1__2__0_chanx_out_150_;
wire [0:0] cbx_1__2__0_chanx_out_151_;
wire [0:0] cbx_1__2__0_chanx_out_152_;
wire [0:0] cbx_1__2__0_chanx_out_153_;
wire [0:0] cbx_1__2__0_chanx_out_154_;
wire [0:0] cbx_1__2__0_chanx_out_155_;
wire [0:0] cbx_1__2__0_chanx_out_156_;
wire [0:0] cbx_1__2__0_chanx_out_157_;
wire [0:0] cbx_1__2__0_chanx_out_158_;
wire [0:0] cbx_1__2__0_chanx_out_159_;
wire [0:0] cbx_1__2__0_chanx_out_15_;
wire [0:0] cbx_1__2__0_chanx_out_160_;
wire [0:0] cbx_1__2__0_chanx_out_161_;
wire [0:0] cbx_1__2__0_chanx_out_162_;
wire [0:0] cbx_1__2__0_chanx_out_163_;
wire [0:0] cbx_1__2__0_chanx_out_164_;
wire [0:0] cbx_1__2__0_chanx_out_165_;
wire [0:0] cbx_1__2__0_chanx_out_166_;
wire [0:0] cbx_1__2__0_chanx_out_167_;
wire [0:0] cbx_1__2__0_chanx_out_168_;
wire [0:0] cbx_1__2__0_chanx_out_169_;
wire [0:0] cbx_1__2__0_chanx_out_16_;
wire [0:0] cbx_1__2__0_chanx_out_170_;
wire [0:0] cbx_1__2__0_chanx_out_171_;
wire [0:0] cbx_1__2__0_chanx_out_172_;
wire [0:0] cbx_1__2__0_chanx_out_173_;
wire [0:0] cbx_1__2__0_chanx_out_174_;
wire [0:0] cbx_1__2__0_chanx_out_175_;
wire [0:0] cbx_1__2__0_chanx_out_176_;
wire [0:0] cbx_1__2__0_chanx_out_177_;
wire [0:0] cbx_1__2__0_chanx_out_178_;
wire [0:0] cbx_1__2__0_chanx_out_179_;
wire [0:0] cbx_1__2__0_chanx_out_17_;
wire [0:0] cbx_1__2__0_chanx_out_180_;
wire [0:0] cbx_1__2__0_chanx_out_181_;
wire [0:0] cbx_1__2__0_chanx_out_182_;
wire [0:0] cbx_1__2__0_chanx_out_183_;
wire [0:0] cbx_1__2__0_chanx_out_184_;
wire [0:0] cbx_1__2__0_chanx_out_185_;
wire [0:0] cbx_1__2__0_chanx_out_186_;
wire [0:0] cbx_1__2__0_chanx_out_187_;
wire [0:0] cbx_1__2__0_chanx_out_188_;
wire [0:0] cbx_1__2__0_chanx_out_189_;
wire [0:0] cbx_1__2__0_chanx_out_18_;
wire [0:0] cbx_1__2__0_chanx_out_190_;
wire [0:0] cbx_1__2__0_chanx_out_191_;
wire [0:0] cbx_1__2__0_chanx_out_192_;
wire [0:0] cbx_1__2__0_chanx_out_193_;
wire [0:0] cbx_1__2__0_chanx_out_194_;
wire [0:0] cbx_1__2__0_chanx_out_195_;
wire [0:0] cbx_1__2__0_chanx_out_196_;
wire [0:0] cbx_1__2__0_chanx_out_197_;
wire [0:0] cbx_1__2__0_chanx_out_198_;
wire [0:0] cbx_1__2__0_chanx_out_199_;
wire [0:0] cbx_1__2__0_chanx_out_19_;
wire [0:0] cbx_1__2__0_chanx_out_1_;
wire [0:0] cbx_1__2__0_chanx_out_20_;
wire [0:0] cbx_1__2__0_chanx_out_21_;
wire [0:0] cbx_1__2__0_chanx_out_22_;
wire [0:0] cbx_1__2__0_chanx_out_23_;
wire [0:0] cbx_1__2__0_chanx_out_24_;
wire [0:0] cbx_1__2__0_chanx_out_25_;
wire [0:0] cbx_1__2__0_chanx_out_26_;
wire [0:0] cbx_1__2__0_chanx_out_27_;
wire [0:0] cbx_1__2__0_chanx_out_28_;
wire [0:0] cbx_1__2__0_chanx_out_29_;
wire [0:0] cbx_1__2__0_chanx_out_2_;
wire [0:0] cbx_1__2__0_chanx_out_30_;
wire [0:0] cbx_1__2__0_chanx_out_31_;
wire [0:0] cbx_1__2__0_chanx_out_32_;
wire [0:0] cbx_1__2__0_chanx_out_33_;
wire [0:0] cbx_1__2__0_chanx_out_34_;
wire [0:0] cbx_1__2__0_chanx_out_35_;
wire [0:0] cbx_1__2__0_chanx_out_36_;
wire [0:0] cbx_1__2__0_chanx_out_37_;
wire [0:0] cbx_1__2__0_chanx_out_38_;
wire [0:0] cbx_1__2__0_chanx_out_39_;
wire [0:0] cbx_1__2__0_chanx_out_3_;
wire [0:0] cbx_1__2__0_chanx_out_40_;
wire [0:0] cbx_1__2__0_chanx_out_41_;
wire [0:0] cbx_1__2__0_chanx_out_42_;
wire [0:0] cbx_1__2__0_chanx_out_43_;
wire [0:0] cbx_1__2__0_chanx_out_44_;
wire [0:0] cbx_1__2__0_chanx_out_45_;
wire [0:0] cbx_1__2__0_chanx_out_46_;
wire [0:0] cbx_1__2__0_chanx_out_47_;
wire [0:0] cbx_1__2__0_chanx_out_48_;
wire [0:0] cbx_1__2__0_chanx_out_49_;
wire [0:0] cbx_1__2__0_chanx_out_4_;
wire [0:0] cbx_1__2__0_chanx_out_50_;
wire [0:0] cbx_1__2__0_chanx_out_51_;
wire [0:0] cbx_1__2__0_chanx_out_52_;
wire [0:0] cbx_1__2__0_chanx_out_53_;
wire [0:0] cbx_1__2__0_chanx_out_54_;
wire [0:0] cbx_1__2__0_chanx_out_55_;
wire [0:0] cbx_1__2__0_chanx_out_56_;
wire [0:0] cbx_1__2__0_chanx_out_57_;
wire [0:0] cbx_1__2__0_chanx_out_58_;
wire [0:0] cbx_1__2__0_chanx_out_59_;
wire [0:0] cbx_1__2__0_chanx_out_5_;
wire [0:0] cbx_1__2__0_chanx_out_60_;
wire [0:0] cbx_1__2__0_chanx_out_61_;
wire [0:0] cbx_1__2__0_chanx_out_62_;
wire [0:0] cbx_1__2__0_chanx_out_63_;
wire [0:0] cbx_1__2__0_chanx_out_64_;
wire [0:0] cbx_1__2__0_chanx_out_65_;
wire [0:0] cbx_1__2__0_chanx_out_66_;
wire [0:0] cbx_1__2__0_chanx_out_67_;
wire [0:0] cbx_1__2__0_chanx_out_68_;
wire [0:0] cbx_1__2__0_chanx_out_69_;
wire [0:0] cbx_1__2__0_chanx_out_6_;
wire [0:0] cbx_1__2__0_chanx_out_70_;
wire [0:0] cbx_1__2__0_chanx_out_71_;
wire [0:0] cbx_1__2__0_chanx_out_72_;
wire [0:0] cbx_1__2__0_chanx_out_73_;
wire [0:0] cbx_1__2__0_chanx_out_74_;
wire [0:0] cbx_1__2__0_chanx_out_75_;
wire [0:0] cbx_1__2__0_chanx_out_76_;
wire [0:0] cbx_1__2__0_chanx_out_77_;
wire [0:0] cbx_1__2__0_chanx_out_78_;
wire [0:0] cbx_1__2__0_chanx_out_79_;
wire [0:0] cbx_1__2__0_chanx_out_7_;
wire [0:0] cbx_1__2__0_chanx_out_80_;
wire [0:0] cbx_1__2__0_chanx_out_81_;
wire [0:0] cbx_1__2__0_chanx_out_82_;
wire [0:0] cbx_1__2__0_chanx_out_83_;
wire [0:0] cbx_1__2__0_chanx_out_84_;
wire [0:0] cbx_1__2__0_chanx_out_85_;
wire [0:0] cbx_1__2__0_chanx_out_86_;
wire [0:0] cbx_1__2__0_chanx_out_87_;
wire [0:0] cbx_1__2__0_chanx_out_88_;
wire [0:0] cbx_1__2__0_chanx_out_89_;
wire [0:0] cbx_1__2__0_chanx_out_8_;
wire [0:0] cbx_1__2__0_chanx_out_90_;
wire [0:0] cbx_1__2__0_chanx_out_91_;
wire [0:0] cbx_1__2__0_chanx_out_92_;
wire [0:0] cbx_1__2__0_chanx_out_93_;
wire [0:0] cbx_1__2__0_chanx_out_94_;
wire [0:0] cbx_1__2__0_chanx_out_95_;
wire [0:0] cbx_1__2__0_chanx_out_96_;
wire [0:0] cbx_1__2__0_chanx_out_97_;
wire [0:0] cbx_1__2__0_chanx_out_98_;
wire [0:0] cbx_1__2__0_chanx_out_99_;
wire [0:0] cbx_1__2__0_chanx_out_9_;
wire [0:0] cbx_1__2__0_top_grid_pin_0_;
wire [0:0] cbx_1__2__1_bottom_grid_pin_42_;
wire [0:0] cbx_1__2__1_bottom_grid_pin_43_;
wire [0:0] cbx_1__2__1_bottom_grid_pin_68_;
wire [0:0] cbx_1__2__1_ccff_tail;
wire [0:0] cbx_1__2__1_chanx_out_0_;
wire [0:0] cbx_1__2__1_chanx_out_100_;
wire [0:0] cbx_1__2__1_chanx_out_101_;
wire [0:0] cbx_1__2__1_chanx_out_102_;
wire [0:0] cbx_1__2__1_chanx_out_103_;
wire [0:0] cbx_1__2__1_chanx_out_104_;
wire [0:0] cbx_1__2__1_chanx_out_105_;
wire [0:0] cbx_1__2__1_chanx_out_106_;
wire [0:0] cbx_1__2__1_chanx_out_107_;
wire [0:0] cbx_1__2__1_chanx_out_108_;
wire [0:0] cbx_1__2__1_chanx_out_109_;
wire [0:0] cbx_1__2__1_chanx_out_10_;
wire [0:0] cbx_1__2__1_chanx_out_110_;
wire [0:0] cbx_1__2__1_chanx_out_111_;
wire [0:0] cbx_1__2__1_chanx_out_112_;
wire [0:0] cbx_1__2__1_chanx_out_113_;
wire [0:0] cbx_1__2__1_chanx_out_114_;
wire [0:0] cbx_1__2__1_chanx_out_115_;
wire [0:0] cbx_1__2__1_chanx_out_116_;
wire [0:0] cbx_1__2__1_chanx_out_117_;
wire [0:0] cbx_1__2__1_chanx_out_118_;
wire [0:0] cbx_1__2__1_chanx_out_119_;
wire [0:0] cbx_1__2__1_chanx_out_11_;
wire [0:0] cbx_1__2__1_chanx_out_120_;
wire [0:0] cbx_1__2__1_chanx_out_121_;
wire [0:0] cbx_1__2__1_chanx_out_122_;
wire [0:0] cbx_1__2__1_chanx_out_123_;
wire [0:0] cbx_1__2__1_chanx_out_124_;
wire [0:0] cbx_1__2__1_chanx_out_125_;
wire [0:0] cbx_1__2__1_chanx_out_126_;
wire [0:0] cbx_1__2__1_chanx_out_127_;
wire [0:0] cbx_1__2__1_chanx_out_128_;
wire [0:0] cbx_1__2__1_chanx_out_129_;
wire [0:0] cbx_1__2__1_chanx_out_12_;
wire [0:0] cbx_1__2__1_chanx_out_130_;
wire [0:0] cbx_1__2__1_chanx_out_131_;
wire [0:0] cbx_1__2__1_chanx_out_132_;
wire [0:0] cbx_1__2__1_chanx_out_133_;
wire [0:0] cbx_1__2__1_chanx_out_134_;
wire [0:0] cbx_1__2__1_chanx_out_135_;
wire [0:0] cbx_1__2__1_chanx_out_136_;
wire [0:0] cbx_1__2__1_chanx_out_137_;
wire [0:0] cbx_1__2__1_chanx_out_138_;
wire [0:0] cbx_1__2__1_chanx_out_139_;
wire [0:0] cbx_1__2__1_chanx_out_13_;
wire [0:0] cbx_1__2__1_chanx_out_140_;
wire [0:0] cbx_1__2__1_chanx_out_141_;
wire [0:0] cbx_1__2__1_chanx_out_142_;
wire [0:0] cbx_1__2__1_chanx_out_143_;
wire [0:0] cbx_1__2__1_chanx_out_144_;
wire [0:0] cbx_1__2__1_chanx_out_145_;
wire [0:0] cbx_1__2__1_chanx_out_146_;
wire [0:0] cbx_1__2__1_chanx_out_147_;
wire [0:0] cbx_1__2__1_chanx_out_148_;
wire [0:0] cbx_1__2__1_chanx_out_149_;
wire [0:0] cbx_1__2__1_chanx_out_14_;
wire [0:0] cbx_1__2__1_chanx_out_150_;
wire [0:0] cbx_1__2__1_chanx_out_151_;
wire [0:0] cbx_1__2__1_chanx_out_152_;
wire [0:0] cbx_1__2__1_chanx_out_153_;
wire [0:0] cbx_1__2__1_chanx_out_154_;
wire [0:0] cbx_1__2__1_chanx_out_155_;
wire [0:0] cbx_1__2__1_chanx_out_156_;
wire [0:0] cbx_1__2__1_chanx_out_157_;
wire [0:0] cbx_1__2__1_chanx_out_158_;
wire [0:0] cbx_1__2__1_chanx_out_159_;
wire [0:0] cbx_1__2__1_chanx_out_15_;
wire [0:0] cbx_1__2__1_chanx_out_160_;
wire [0:0] cbx_1__2__1_chanx_out_161_;
wire [0:0] cbx_1__2__1_chanx_out_162_;
wire [0:0] cbx_1__2__1_chanx_out_163_;
wire [0:0] cbx_1__2__1_chanx_out_164_;
wire [0:0] cbx_1__2__1_chanx_out_165_;
wire [0:0] cbx_1__2__1_chanx_out_166_;
wire [0:0] cbx_1__2__1_chanx_out_167_;
wire [0:0] cbx_1__2__1_chanx_out_168_;
wire [0:0] cbx_1__2__1_chanx_out_169_;
wire [0:0] cbx_1__2__1_chanx_out_16_;
wire [0:0] cbx_1__2__1_chanx_out_170_;
wire [0:0] cbx_1__2__1_chanx_out_171_;
wire [0:0] cbx_1__2__1_chanx_out_172_;
wire [0:0] cbx_1__2__1_chanx_out_173_;
wire [0:0] cbx_1__2__1_chanx_out_174_;
wire [0:0] cbx_1__2__1_chanx_out_175_;
wire [0:0] cbx_1__2__1_chanx_out_176_;
wire [0:0] cbx_1__2__1_chanx_out_177_;
wire [0:0] cbx_1__2__1_chanx_out_178_;
wire [0:0] cbx_1__2__1_chanx_out_179_;
wire [0:0] cbx_1__2__1_chanx_out_17_;
wire [0:0] cbx_1__2__1_chanx_out_180_;
wire [0:0] cbx_1__2__1_chanx_out_181_;
wire [0:0] cbx_1__2__1_chanx_out_182_;
wire [0:0] cbx_1__2__1_chanx_out_183_;
wire [0:0] cbx_1__2__1_chanx_out_184_;
wire [0:0] cbx_1__2__1_chanx_out_185_;
wire [0:0] cbx_1__2__1_chanx_out_186_;
wire [0:0] cbx_1__2__1_chanx_out_187_;
wire [0:0] cbx_1__2__1_chanx_out_188_;
wire [0:0] cbx_1__2__1_chanx_out_189_;
wire [0:0] cbx_1__2__1_chanx_out_18_;
wire [0:0] cbx_1__2__1_chanx_out_190_;
wire [0:0] cbx_1__2__1_chanx_out_191_;
wire [0:0] cbx_1__2__1_chanx_out_192_;
wire [0:0] cbx_1__2__1_chanx_out_193_;
wire [0:0] cbx_1__2__1_chanx_out_194_;
wire [0:0] cbx_1__2__1_chanx_out_195_;
wire [0:0] cbx_1__2__1_chanx_out_196_;
wire [0:0] cbx_1__2__1_chanx_out_197_;
wire [0:0] cbx_1__2__1_chanx_out_198_;
wire [0:0] cbx_1__2__1_chanx_out_199_;
wire [0:0] cbx_1__2__1_chanx_out_19_;
wire [0:0] cbx_1__2__1_chanx_out_1_;
wire [0:0] cbx_1__2__1_chanx_out_20_;
wire [0:0] cbx_1__2__1_chanx_out_21_;
wire [0:0] cbx_1__2__1_chanx_out_22_;
wire [0:0] cbx_1__2__1_chanx_out_23_;
wire [0:0] cbx_1__2__1_chanx_out_24_;
wire [0:0] cbx_1__2__1_chanx_out_25_;
wire [0:0] cbx_1__2__1_chanx_out_26_;
wire [0:0] cbx_1__2__1_chanx_out_27_;
wire [0:0] cbx_1__2__1_chanx_out_28_;
wire [0:0] cbx_1__2__1_chanx_out_29_;
wire [0:0] cbx_1__2__1_chanx_out_2_;
wire [0:0] cbx_1__2__1_chanx_out_30_;
wire [0:0] cbx_1__2__1_chanx_out_31_;
wire [0:0] cbx_1__2__1_chanx_out_32_;
wire [0:0] cbx_1__2__1_chanx_out_33_;
wire [0:0] cbx_1__2__1_chanx_out_34_;
wire [0:0] cbx_1__2__1_chanx_out_35_;
wire [0:0] cbx_1__2__1_chanx_out_36_;
wire [0:0] cbx_1__2__1_chanx_out_37_;
wire [0:0] cbx_1__2__1_chanx_out_38_;
wire [0:0] cbx_1__2__1_chanx_out_39_;
wire [0:0] cbx_1__2__1_chanx_out_3_;
wire [0:0] cbx_1__2__1_chanx_out_40_;
wire [0:0] cbx_1__2__1_chanx_out_41_;
wire [0:0] cbx_1__2__1_chanx_out_42_;
wire [0:0] cbx_1__2__1_chanx_out_43_;
wire [0:0] cbx_1__2__1_chanx_out_44_;
wire [0:0] cbx_1__2__1_chanx_out_45_;
wire [0:0] cbx_1__2__1_chanx_out_46_;
wire [0:0] cbx_1__2__1_chanx_out_47_;
wire [0:0] cbx_1__2__1_chanx_out_48_;
wire [0:0] cbx_1__2__1_chanx_out_49_;
wire [0:0] cbx_1__2__1_chanx_out_4_;
wire [0:0] cbx_1__2__1_chanx_out_50_;
wire [0:0] cbx_1__2__1_chanx_out_51_;
wire [0:0] cbx_1__2__1_chanx_out_52_;
wire [0:0] cbx_1__2__1_chanx_out_53_;
wire [0:0] cbx_1__2__1_chanx_out_54_;
wire [0:0] cbx_1__2__1_chanx_out_55_;
wire [0:0] cbx_1__2__1_chanx_out_56_;
wire [0:0] cbx_1__2__1_chanx_out_57_;
wire [0:0] cbx_1__2__1_chanx_out_58_;
wire [0:0] cbx_1__2__1_chanx_out_59_;
wire [0:0] cbx_1__2__1_chanx_out_5_;
wire [0:0] cbx_1__2__1_chanx_out_60_;
wire [0:0] cbx_1__2__1_chanx_out_61_;
wire [0:0] cbx_1__2__1_chanx_out_62_;
wire [0:0] cbx_1__2__1_chanx_out_63_;
wire [0:0] cbx_1__2__1_chanx_out_64_;
wire [0:0] cbx_1__2__1_chanx_out_65_;
wire [0:0] cbx_1__2__1_chanx_out_66_;
wire [0:0] cbx_1__2__1_chanx_out_67_;
wire [0:0] cbx_1__2__1_chanx_out_68_;
wire [0:0] cbx_1__2__1_chanx_out_69_;
wire [0:0] cbx_1__2__1_chanx_out_6_;
wire [0:0] cbx_1__2__1_chanx_out_70_;
wire [0:0] cbx_1__2__1_chanx_out_71_;
wire [0:0] cbx_1__2__1_chanx_out_72_;
wire [0:0] cbx_1__2__1_chanx_out_73_;
wire [0:0] cbx_1__2__1_chanx_out_74_;
wire [0:0] cbx_1__2__1_chanx_out_75_;
wire [0:0] cbx_1__2__1_chanx_out_76_;
wire [0:0] cbx_1__2__1_chanx_out_77_;
wire [0:0] cbx_1__2__1_chanx_out_78_;
wire [0:0] cbx_1__2__1_chanx_out_79_;
wire [0:0] cbx_1__2__1_chanx_out_7_;
wire [0:0] cbx_1__2__1_chanx_out_80_;
wire [0:0] cbx_1__2__1_chanx_out_81_;
wire [0:0] cbx_1__2__1_chanx_out_82_;
wire [0:0] cbx_1__2__1_chanx_out_83_;
wire [0:0] cbx_1__2__1_chanx_out_84_;
wire [0:0] cbx_1__2__1_chanx_out_85_;
wire [0:0] cbx_1__2__1_chanx_out_86_;
wire [0:0] cbx_1__2__1_chanx_out_87_;
wire [0:0] cbx_1__2__1_chanx_out_88_;
wire [0:0] cbx_1__2__1_chanx_out_89_;
wire [0:0] cbx_1__2__1_chanx_out_8_;
wire [0:0] cbx_1__2__1_chanx_out_90_;
wire [0:0] cbx_1__2__1_chanx_out_91_;
wire [0:0] cbx_1__2__1_chanx_out_92_;
wire [0:0] cbx_1__2__1_chanx_out_93_;
wire [0:0] cbx_1__2__1_chanx_out_94_;
wire [0:0] cbx_1__2__1_chanx_out_95_;
wire [0:0] cbx_1__2__1_chanx_out_96_;
wire [0:0] cbx_1__2__1_chanx_out_97_;
wire [0:0] cbx_1__2__1_chanx_out_98_;
wire [0:0] cbx_1__2__1_chanx_out_99_;
wire [0:0] cbx_1__2__1_chanx_out_9_;
wire [0:0] cbx_1__2__1_top_grid_pin_0_;
wire [0:0] cby_0__1__0_ccff_tail;
wire [0:0] cby_0__1__0_chany_out_0_;
wire [0:0] cby_0__1__0_chany_out_100_;
wire [0:0] cby_0__1__0_chany_out_101_;
wire [0:0] cby_0__1__0_chany_out_102_;
wire [0:0] cby_0__1__0_chany_out_103_;
wire [0:0] cby_0__1__0_chany_out_104_;
wire [0:0] cby_0__1__0_chany_out_105_;
wire [0:0] cby_0__1__0_chany_out_106_;
wire [0:0] cby_0__1__0_chany_out_107_;
wire [0:0] cby_0__1__0_chany_out_108_;
wire [0:0] cby_0__1__0_chany_out_109_;
wire [0:0] cby_0__1__0_chany_out_10_;
wire [0:0] cby_0__1__0_chany_out_110_;
wire [0:0] cby_0__1__0_chany_out_111_;
wire [0:0] cby_0__1__0_chany_out_112_;
wire [0:0] cby_0__1__0_chany_out_113_;
wire [0:0] cby_0__1__0_chany_out_114_;
wire [0:0] cby_0__1__0_chany_out_115_;
wire [0:0] cby_0__1__0_chany_out_116_;
wire [0:0] cby_0__1__0_chany_out_117_;
wire [0:0] cby_0__1__0_chany_out_118_;
wire [0:0] cby_0__1__0_chany_out_119_;
wire [0:0] cby_0__1__0_chany_out_11_;
wire [0:0] cby_0__1__0_chany_out_120_;
wire [0:0] cby_0__1__0_chany_out_121_;
wire [0:0] cby_0__1__0_chany_out_122_;
wire [0:0] cby_0__1__0_chany_out_123_;
wire [0:0] cby_0__1__0_chany_out_124_;
wire [0:0] cby_0__1__0_chany_out_125_;
wire [0:0] cby_0__1__0_chany_out_126_;
wire [0:0] cby_0__1__0_chany_out_127_;
wire [0:0] cby_0__1__0_chany_out_128_;
wire [0:0] cby_0__1__0_chany_out_129_;
wire [0:0] cby_0__1__0_chany_out_12_;
wire [0:0] cby_0__1__0_chany_out_130_;
wire [0:0] cby_0__1__0_chany_out_131_;
wire [0:0] cby_0__1__0_chany_out_132_;
wire [0:0] cby_0__1__0_chany_out_133_;
wire [0:0] cby_0__1__0_chany_out_134_;
wire [0:0] cby_0__1__0_chany_out_135_;
wire [0:0] cby_0__1__0_chany_out_136_;
wire [0:0] cby_0__1__0_chany_out_137_;
wire [0:0] cby_0__1__0_chany_out_138_;
wire [0:0] cby_0__1__0_chany_out_139_;
wire [0:0] cby_0__1__0_chany_out_13_;
wire [0:0] cby_0__1__0_chany_out_140_;
wire [0:0] cby_0__1__0_chany_out_141_;
wire [0:0] cby_0__1__0_chany_out_142_;
wire [0:0] cby_0__1__0_chany_out_143_;
wire [0:0] cby_0__1__0_chany_out_144_;
wire [0:0] cby_0__1__0_chany_out_145_;
wire [0:0] cby_0__1__0_chany_out_146_;
wire [0:0] cby_0__1__0_chany_out_147_;
wire [0:0] cby_0__1__0_chany_out_148_;
wire [0:0] cby_0__1__0_chany_out_149_;
wire [0:0] cby_0__1__0_chany_out_14_;
wire [0:0] cby_0__1__0_chany_out_150_;
wire [0:0] cby_0__1__0_chany_out_151_;
wire [0:0] cby_0__1__0_chany_out_152_;
wire [0:0] cby_0__1__0_chany_out_153_;
wire [0:0] cby_0__1__0_chany_out_154_;
wire [0:0] cby_0__1__0_chany_out_155_;
wire [0:0] cby_0__1__0_chany_out_156_;
wire [0:0] cby_0__1__0_chany_out_157_;
wire [0:0] cby_0__1__0_chany_out_158_;
wire [0:0] cby_0__1__0_chany_out_159_;
wire [0:0] cby_0__1__0_chany_out_15_;
wire [0:0] cby_0__1__0_chany_out_160_;
wire [0:0] cby_0__1__0_chany_out_161_;
wire [0:0] cby_0__1__0_chany_out_162_;
wire [0:0] cby_0__1__0_chany_out_163_;
wire [0:0] cby_0__1__0_chany_out_164_;
wire [0:0] cby_0__1__0_chany_out_165_;
wire [0:0] cby_0__1__0_chany_out_166_;
wire [0:0] cby_0__1__0_chany_out_167_;
wire [0:0] cby_0__1__0_chany_out_168_;
wire [0:0] cby_0__1__0_chany_out_169_;
wire [0:0] cby_0__1__0_chany_out_16_;
wire [0:0] cby_0__1__0_chany_out_170_;
wire [0:0] cby_0__1__0_chany_out_171_;
wire [0:0] cby_0__1__0_chany_out_172_;
wire [0:0] cby_0__1__0_chany_out_173_;
wire [0:0] cby_0__1__0_chany_out_174_;
wire [0:0] cby_0__1__0_chany_out_175_;
wire [0:0] cby_0__1__0_chany_out_176_;
wire [0:0] cby_0__1__0_chany_out_177_;
wire [0:0] cby_0__1__0_chany_out_178_;
wire [0:0] cby_0__1__0_chany_out_179_;
wire [0:0] cby_0__1__0_chany_out_17_;
wire [0:0] cby_0__1__0_chany_out_180_;
wire [0:0] cby_0__1__0_chany_out_181_;
wire [0:0] cby_0__1__0_chany_out_182_;
wire [0:0] cby_0__1__0_chany_out_183_;
wire [0:0] cby_0__1__0_chany_out_184_;
wire [0:0] cby_0__1__0_chany_out_185_;
wire [0:0] cby_0__1__0_chany_out_186_;
wire [0:0] cby_0__1__0_chany_out_187_;
wire [0:0] cby_0__1__0_chany_out_188_;
wire [0:0] cby_0__1__0_chany_out_189_;
wire [0:0] cby_0__1__0_chany_out_18_;
wire [0:0] cby_0__1__0_chany_out_190_;
wire [0:0] cby_0__1__0_chany_out_191_;
wire [0:0] cby_0__1__0_chany_out_192_;
wire [0:0] cby_0__1__0_chany_out_193_;
wire [0:0] cby_0__1__0_chany_out_194_;
wire [0:0] cby_0__1__0_chany_out_195_;
wire [0:0] cby_0__1__0_chany_out_196_;
wire [0:0] cby_0__1__0_chany_out_197_;
wire [0:0] cby_0__1__0_chany_out_198_;
wire [0:0] cby_0__1__0_chany_out_199_;
wire [0:0] cby_0__1__0_chany_out_19_;
wire [0:0] cby_0__1__0_chany_out_1_;
wire [0:0] cby_0__1__0_chany_out_20_;
wire [0:0] cby_0__1__0_chany_out_21_;
wire [0:0] cby_0__1__0_chany_out_22_;
wire [0:0] cby_0__1__0_chany_out_23_;
wire [0:0] cby_0__1__0_chany_out_24_;
wire [0:0] cby_0__1__0_chany_out_25_;
wire [0:0] cby_0__1__0_chany_out_26_;
wire [0:0] cby_0__1__0_chany_out_27_;
wire [0:0] cby_0__1__0_chany_out_28_;
wire [0:0] cby_0__1__0_chany_out_29_;
wire [0:0] cby_0__1__0_chany_out_2_;
wire [0:0] cby_0__1__0_chany_out_30_;
wire [0:0] cby_0__1__0_chany_out_31_;
wire [0:0] cby_0__1__0_chany_out_32_;
wire [0:0] cby_0__1__0_chany_out_33_;
wire [0:0] cby_0__1__0_chany_out_34_;
wire [0:0] cby_0__1__0_chany_out_35_;
wire [0:0] cby_0__1__0_chany_out_36_;
wire [0:0] cby_0__1__0_chany_out_37_;
wire [0:0] cby_0__1__0_chany_out_38_;
wire [0:0] cby_0__1__0_chany_out_39_;
wire [0:0] cby_0__1__0_chany_out_3_;
wire [0:0] cby_0__1__0_chany_out_40_;
wire [0:0] cby_0__1__0_chany_out_41_;
wire [0:0] cby_0__1__0_chany_out_42_;
wire [0:0] cby_0__1__0_chany_out_43_;
wire [0:0] cby_0__1__0_chany_out_44_;
wire [0:0] cby_0__1__0_chany_out_45_;
wire [0:0] cby_0__1__0_chany_out_46_;
wire [0:0] cby_0__1__0_chany_out_47_;
wire [0:0] cby_0__1__0_chany_out_48_;
wire [0:0] cby_0__1__0_chany_out_49_;
wire [0:0] cby_0__1__0_chany_out_4_;
wire [0:0] cby_0__1__0_chany_out_50_;
wire [0:0] cby_0__1__0_chany_out_51_;
wire [0:0] cby_0__1__0_chany_out_52_;
wire [0:0] cby_0__1__0_chany_out_53_;
wire [0:0] cby_0__1__0_chany_out_54_;
wire [0:0] cby_0__1__0_chany_out_55_;
wire [0:0] cby_0__1__0_chany_out_56_;
wire [0:0] cby_0__1__0_chany_out_57_;
wire [0:0] cby_0__1__0_chany_out_58_;
wire [0:0] cby_0__1__0_chany_out_59_;
wire [0:0] cby_0__1__0_chany_out_5_;
wire [0:0] cby_0__1__0_chany_out_60_;
wire [0:0] cby_0__1__0_chany_out_61_;
wire [0:0] cby_0__1__0_chany_out_62_;
wire [0:0] cby_0__1__0_chany_out_63_;
wire [0:0] cby_0__1__0_chany_out_64_;
wire [0:0] cby_0__1__0_chany_out_65_;
wire [0:0] cby_0__1__0_chany_out_66_;
wire [0:0] cby_0__1__0_chany_out_67_;
wire [0:0] cby_0__1__0_chany_out_68_;
wire [0:0] cby_0__1__0_chany_out_69_;
wire [0:0] cby_0__1__0_chany_out_6_;
wire [0:0] cby_0__1__0_chany_out_70_;
wire [0:0] cby_0__1__0_chany_out_71_;
wire [0:0] cby_0__1__0_chany_out_72_;
wire [0:0] cby_0__1__0_chany_out_73_;
wire [0:0] cby_0__1__0_chany_out_74_;
wire [0:0] cby_0__1__0_chany_out_75_;
wire [0:0] cby_0__1__0_chany_out_76_;
wire [0:0] cby_0__1__0_chany_out_77_;
wire [0:0] cby_0__1__0_chany_out_78_;
wire [0:0] cby_0__1__0_chany_out_79_;
wire [0:0] cby_0__1__0_chany_out_7_;
wire [0:0] cby_0__1__0_chany_out_80_;
wire [0:0] cby_0__1__0_chany_out_81_;
wire [0:0] cby_0__1__0_chany_out_82_;
wire [0:0] cby_0__1__0_chany_out_83_;
wire [0:0] cby_0__1__0_chany_out_84_;
wire [0:0] cby_0__1__0_chany_out_85_;
wire [0:0] cby_0__1__0_chany_out_86_;
wire [0:0] cby_0__1__0_chany_out_87_;
wire [0:0] cby_0__1__0_chany_out_88_;
wire [0:0] cby_0__1__0_chany_out_89_;
wire [0:0] cby_0__1__0_chany_out_8_;
wire [0:0] cby_0__1__0_chany_out_90_;
wire [0:0] cby_0__1__0_chany_out_91_;
wire [0:0] cby_0__1__0_chany_out_92_;
wire [0:0] cby_0__1__0_chany_out_93_;
wire [0:0] cby_0__1__0_chany_out_94_;
wire [0:0] cby_0__1__0_chany_out_95_;
wire [0:0] cby_0__1__0_chany_out_96_;
wire [0:0] cby_0__1__0_chany_out_97_;
wire [0:0] cby_0__1__0_chany_out_98_;
wire [0:0] cby_0__1__0_chany_out_99_;
wire [0:0] cby_0__1__0_chany_out_9_;
wire [0:0] cby_0__1__0_left_grid_pin_0_;
wire [0:0] cby_0__1__1_ccff_tail;
wire [0:0] cby_0__1__1_chany_out_0_;
wire [0:0] cby_0__1__1_chany_out_100_;
wire [0:0] cby_0__1__1_chany_out_101_;
wire [0:0] cby_0__1__1_chany_out_102_;
wire [0:0] cby_0__1__1_chany_out_103_;
wire [0:0] cby_0__1__1_chany_out_104_;
wire [0:0] cby_0__1__1_chany_out_105_;
wire [0:0] cby_0__1__1_chany_out_106_;
wire [0:0] cby_0__1__1_chany_out_107_;
wire [0:0] cby_0__1__1_chany_out_108_;
wire [0:0] cby_0__1__1_chany_out_109_;
wire [0:0] cby_0__1__1_chany_out_10_;
wire [0:0] cby_0__1__1_chany_out_110_;
wire [0:0] cby_0__1__1_chany_out_111_;
wire [0:0] cby_0__1__1_chany_out_112_;
wire [0:0] cby_0__1__1_chany_out_113_;
wire [0:0] cby_0__1__1_chany_out_114_;
wire [0:0] cby_0__1__1_chany_out_115_;
wire [0:0] cby_0__1__1_chany_out_116_;
wire [0:0] cby_0__1__1_chany_out_117_;
wire [0:0] cby_0__1__1_chany_out_118_;
wire [0:0] cby_0__1__1_chany_out_119_;
wire [0:0] cby_0__1__1_chany_out_11_;
wire [0:0] cby_0__1__1_chany_out_120_;
wire [0:0] cby_0__1__1_chany_out_121_;
wire [0:0] cby_0__1__1_chany_out_122_;
wire [0:0] cby_0__1__1_chany_out_123_;
wire [0:0] cby_0__1__1_chany_out_124_;
wire [0:0] cby_0__1__1_chany_out_125_;
wire [0:0] cby_0__1__1_chany_out_126_;
wire [0:0] cby_0__1__1_chany_out_127_;
wire [0:0] cby_0__1__1_chany_out_128_;
wire [0:0] cby_0__1__1_chany_out_129_;
wire [0:0] cby_0__1__1_chany_out_12_;
wire [0:0] cby_0__1__1_chany_out_130_;
wire [0:0] cby_0__1__1_chany_out_131_;
wire [0:0] cby_0__1__1_chany_out_132_;
wire [0:0] cby_0__1__1_chany_out_133_;
wire [0:0] cby_0__1__1_chany_out_134_;
wire [0:0] cby_0__1__1_chany_out_135_;
wire [0:0] cby_0__1__1_chany_out_136_;
wire [0:0] cby_0__1__1_chany_out_137_;
wire [0:0] cby_0__1__1_chany_out_138_;
wire [0:0] cby_0__1__1_chany_out_139_;
wire [0:0] cby_0__1__1_chany_out_13_;
wire [0:0] cby_0__1__1_chany_out_140_;
wire [0:0] cby_0__1__1_chany_out_141_;
wire [0:0] cby_0__1__1_chany_out_142_;
wire [0:0] cby_0__1__1_chany_out_143_;
wire [0:0] cby_0__1__1_chany_out_144_;
wire [0:0] cby_0__1__1_chany_out_145_;
wire [0:0] cby_0__1__1_chany_out_146_;
wire [0:0] cby_0__1__1_chany_out_147_;
wire [0:0] cby_0__1__1_chany_out_148_;
wire [0:0] cby_0__1__1_chany_out_149_;
wire [0:0] cby_0__1__1_chany_out_14_;
wire [0:0] cby_0__1__1_chany_out_150_;
wire [0:0] cby_0__1__1_chany_out_151_;
wire [0:0] cby_0__1__1_chany_out_152_;
wire [0:0] cby_0__1__1_chany_out_153_;
wire [0:0] cby_0__1__1_chany_out_154_;
wire [0:0] cby_0__1__1_chany_out_155_;
wire [0:0] cby_0__1__1_chany_out_156_;
wire [0:0] cby_0__1__1_chany_out_157_;
wire [0:0] cby_0__1__1_chany_out_158_;
wire [0:0] cby_0__1__1_chany_out_159_;
wire [0:0] cby_0__1__1_chany_out_15_;
wire [0:0] cby_0__1__1_chany_out_160_;
wire [0:0] cby_0__1__1_chany_out_161_;
wire [0:0] cby_0__1__1_chany_out_162_;
wire [0:0] cby_0__1__1_chany_out_163_;
wire [0:0] cby_0__1__1_chany_out_164_;
wire [0:0] cby_0__1__1_chany_out_165_;
wire [0:0] cby_0__1__1_chany_out_166_;
wire [0:0] cby_0__1__1_chany_out_167_;
wire [0:0] cby_0__1__1_chany_out_168_;
wire [0:0] cby_0__1__1_chany_out_169_;
wire [0:0] cby_0__1__1_chany_out_16_;
wire [0:0] cby_0__1__1_chany_out_170_;
wire [0:0] cby_0__1__1_chany_out_171_;
wire [0:0] cby_0__1__1_chany_out_172_;
wire [0:0] cby_0__1__1_chany_out_173_;
wire [0:0] cby_0__1__1_chany_out_174_;
wire [0:0] cby_0__1__1_chany_out_175_;
wire [0:0] cby_0__1__1_chany_out_176_;
wire [0:0] cby_0__1__1_chany_out_177_;
wire [0:0] cby_0__1__1_chany_out_178_;
wire [0:0] cby_0__1__1_chany_out_179_;
wire [0:0] cby_0__1__1_chany_out_17_;
wire [0:0] cby_0__1__1_chany_out_180_;
wire [0:0] cby_0__1__1_chany_out_181_;
wire [0:0] cby_0__1__1_chany_out_182_;
wire [0:0] cby_0__1__1_chany_out_183_;
wire [0:0] cby_0__1__1_chany_out_184_;
wire [0:0] cby_0__1__1_chany_out_185_;
wire [0:0] cby_0__1__1_chany_out_186_;
wire [0:0] cby_0__1__1_chany_out_187_;
wire [0:0] cby_0__1__1_chany_out_188_;
wire [0:0] cby_0__1__1_chany_out_189_;
wire [0:0] cby_0__1__1_chany_out_18_;
wire [0:0] cby_0__1__1_chany_out_190_;
wire [0:0] cby_0__1__1_chany_out_191_;
wire [0:0] cby_0__1__1_chany_out_192_;
wire [0:0] cby_0__1__1_chany_out_193_;
wire [0:0] cby_0__1__1_chany_out_194_;
wire [0:0] cby_0__1__1_chany_out_195_;
wire [0:0] cby_0__1__1_chany_out_196_;
wire [0:0] cby_0__1__1_chany_out_197_;
wire [0:0] cby_0__1__1_chany_out_198_;
wire [0:0] cby_0__1__1_chany_out_199_;
wire [0:0] cby_0__1__1_chany_out_19_;
wire [0:0] cby_0__1__1_chany_out_1_;
wire [0:0] cby_0__1__1_chany_out_20_;
wire [0:0] cby_0__1__1_chany_out_21_;
wire [0:0] cby_0__1__1_chany_out_22_;
wire [0:0] cby_0__1__1_chany_out_23_;
wire [0:0] cby_0__1__1_chany_out_24_;
wire [0:0] cby_0__1__1_chany_out_25_;
wire [0:0] cby_0__1__1_chany_out_26_;
wire [0:0] cby_0__1__1_chany_out_27_;
wire [0:0] cby_0__1__1_chany_out_28_;
wire [0:0] cby_0__1__1_chany_out_29_;
wire [0:0] cby_0__1__1_chany_out_2_;
wire [0:0] cby_0__1__1_chany_out_30_;
wire [0:0] cby_0__1__1_chany_out_31_;
wire [0:0] cby_0__1__1_chany_out_32_;
wire [0:0] cby_0__1__1_chany_out_33_;
wire [0:0] cby_0__1__1_chany_out_34_;
wire [0:0] cby_0__1__1_chany_out_35_;
wire [0:0] cby_0__1__1_chany_out_36_;
wire [0:0] cby_0__1__1_chany_out_37_;
wire [0:0] cby_0__1__1_chany_out_38_;
wire [0:0] cby_0__1__1_chany_out_39_;
wire [0:0] cby_0__1__1_chany_out_3_;
wire [0:0] cby_0__1__1_chany_out_40_;
wire [0:0] cby_0__1__1_chany_out_41_;
wire [0:0] cby_0__1__1_chany_out_42_;
wire [0:0] cby_0__1__1_chany_out_43_;
wire [0:0] cby_0__1__1_chany_out_44_;
wire [0:0] cby_0__1__1_chany_out_45_;
wire [0:0] cby_0__1__1_chany_out_46_;
wire [0:0] cby_0__1__1_chany_out_47_;
wire [0:0] cby_0__1__1_chany_out_48_;
wire [0:0] cby_0__1__1_chany_out_49_;
wire [0:0] cby_0__1__1_chany_out_4_;
wire [0:0] cby_0__1__1_chany_out_50_;
wire [0:0] cby_0__1__1_chany_out_51_;
wire [0:0] cby_0__1__1_chany_out_52_;
wire [0:0] cby_0__1__1_chany_out_53_;
wire [0:0] cby_0__1__1_chany_out_54_;
wire [0:0] cby_0__1__1_chany_out_55_;
wire [0:0] cby_0__1__1_chany_out_56_;
wire [0:0] cby_0__1__1_chany_out_57_;
wire [0:0] cby_0__1__1_chany_out_58_;
wire [0:0] cby_0__1__1_chany_out_59_;
wire [0:0] cby_0__1__1_chany_out_5_;
wire [0:0] cby_0__1__1_chany_out_60_;
wire [0:0] cby_0__1__1_chany_out_61_;
wire [0:0] cby_0__1__1_chany_out_62_;
wire [0:0] cby_0__1__1_chany_out_63_;
wire [0:0] cby_0__1__1_chany_out_64_;
wire [0:0] cby_0__1__1_chany_out_65_;
wire [0:0] cby_0__1__1_chany_out_66_;
wire [0:0] cby_0__1__1_chany_out_67_;
wire [0:0] cby_0__1__1_chany_out_68_;
wire [0:0] cby_0__1__1_chany_out_69_;
wire [0:0] cby_0__1__1_chany_out_6_;
wire [0:0] cby_0__1__1_chany_out_70_;
wire [0:0] cby_0__1__1_chany_out_71_;
wire [0:0] cby_0__1__1_chany_out_72_;
wire [0:0] cby_0__1__1_chany_out_73_;
wire [0:0] cby_0__1__1_chany_out_74_;
wire [0:0] cby_0__1__1_chany_out_75_;
wire [0:0] cby_0__1__1_chany_out_76_;
wire [0:0] cby_0__1__1_chany_out_77_;
wire [0:0] cby_0__1__1_chany_out_78_;
wire [0:0] cby_0__1__1_chany_out_79_;
wire [0:0] cby_0__1__1_chany_out_7_;
wire [0:0] cby_0__1__1_chany_out_80_;
wire [0:0] cby_0__1__1_chany_out_81_;
wire [0:0] cby_0__1__1_chany_out_82_;
wire [0:0] cby_0__1__1_chany_out_83_;
wire [0:0] cby_0__1__1_chany_out_84_;
wire [0:0] cby_0__1__1_chany_out_85_;
wire [0:0] cby_0__1__1_chany_out_86_;
wire [0:0] cby_0__1__1_chany_out_87_;
wire [0:0] cby_0__1__1_chany_out_88_;
wire [0:0] cby_0__1__1_chany_out_89_;
wire [0:0] cby_0__1__1_chany_out_8_;
wire [0:0] cby_0__1__1_chany_out_90_;
wire [0:0] cby_0__1__1_chany_out_91_;
wire [0:0] cby_0__1__1_chany_out_92_;
wire [0:0] cby_0__1__1_chany_out_93_;
wire [0:0] cby_0__1__1_chany_out_94_;
wire [0:0] cby_0__1__1_chany_out_95_;
wire [0:0] cby_0__1__1_chany_out_96_;
wire [0:0] cby_0__1__1_chany_out_97_;
wire [0:0] cby_0__1__1_chany_out_98_;
wire [0:0] cby_0__1__1_chany_out_99_;
wire [0:0] cby_0__1__1_chany_out_9_;
wire [0:0] cby_0__1__1_left_grid_pin_0_;
wire [0:0] cby_1__1__0_ccff_tail;
wire [0:0] cby_1__1__0_chany_out_0_;
wire [0:0] cby_1__1__0_chany_out_100_;
wire [0:0] cby_1__1__0_chany_out_101_;
wire [0:0] cby_1__1__0_chany_out_102_;
wire [0:0] cby_1__1__0_chany_out_103_;
wire [0:0] cby_1__1__0_chany_out_104_;
wire [0:0] cby_1__1__0_chany_out_105_;
wire [0:0] cby_1__1__0_chany_out_106_;
wire [0:0] cby_1__1__0_chany_out_107_;
wire [0:0] cby_1__1__0_chany_out_108_;
wire [0:0] cby_1__1__0_chany_out_109_;
wire [0:0] cby_1__1__0_chany_out_10_;
wire [0:0] cby_1__1__0_chany_out_110_;
wire [0:0] cby_1__1__0_chany_out_111_;
wire [0:0] cby_1__1__0_chany_out_112_;
wire [0:0] cby_1__1__0_chany_out_113_;
wire [0:0] cby_1__1__0_chany_out_114_;
wire [0:0] cby_1__1__0_chany_out_115_;
wire [0:0] cby_1__1__0_chany_out_116_;
wire [0:0] cby_1__1__0_chany_out_117_;
wire [0:0] cby_1__1__0_chany_out_118_;
wire [0:0] cby_1__1__0_chany_out_119_;
wire [0:0] cby_1__1__0_chany_out_11_;
wire [0:0] cby_1__1__0_chany_out_120_;
wire [0:0] cby_1__1__0_chany_out_121_;
wire [0:0] cby_1__1__0_chany_out_122_;
wire [0:0] cby_1__1__0_chany_out_123_;
wire [0:0] cby_1__1__0_chany_out_124_;
wire [0:0] cby_1__1__0_chany_out_125_;
wire [0:0] cby_1__1__0_chany_out_126_;
wire [0:0] cby_1__1__0_chany_out_127_;
wire [0:0] cby_1__1__0_chany_out_128_;
wire [0:0] cby_1__1__0_chany_out_129_;
wire [0:0] cby_1__1__0_chany_out_12_;
wire [0:0] cby_1__1__0_chany_out_130_;
wire [0:0] cby_1__1__0_chany_out_131_;
wire [0:0] cby_1__1__0_chany_out_132_;
wire [0:0] cby_1__1__0_chany_out_133_;
wire [0:0] cby_1__1__0_chany_out_134_;
wire [0:0] cby_1__1__0_chany_out_135_;
wire [0:0] cby_1__1__0_chany_out_136_;
wire [0:0] cby_1__1__0_chany_out_137_;
wire [0:0] cby_1__1__0_chany_out_138_;
wire [0:0] cby_1__1__0_chany_out_139_;
wire [0:0] cby_1__1__0_chany_out_13_;
wire [0:0] cby_1__1__0_chany_out_140_;
wire [0:0] cby_1__1__0_chany_out_141_;
wire [0:0] cby_1__1__0_chany_out_142_;
wire [0:0] cby_1__1__0_chany_out_143_;
wire [0:0] cby_1__1__0_chany_out_144_;
wire [0:0] cby_1__1__0_chany_out_145_;
wire [0:0] cby_1__1__0_chany_out_146_;
wire [0:0] cby_1__1__0_chany_out_147_;
wire [0:0] cby_1__1__0_chany_out_148_;
wire [0:0] cby_1__1__0_chany_out_149_;
wire [0:0] cby_1__1__0_chany_out_14_;
wire [0:0] cby_1__1__0_chany_out_150_;
wire [0:0] cby_1__1__0_chany_out_151_;
wire [0:0] cby_1__1__0_chany_out_152_;
wire [0:0] cby_1__1__0_chany_out_153_;
wire [0:0] cby_1__1__0_chany_out_154_;
wire [0:0] cby_1__1__0_chany_out_155_;
wire [0:0] cby_1__1__0_chany_out_156_;
wire [0:0] cby_1__1__0_chany_out_157_;
wire [0:0] cby_1__1__0_chany_out_158_;
wire [0:0] cby_1__1__0_chany_out_159_;
wire [0:0] cby_1__1__0_chany_out_15_;
wire [0:0] cby_1__1__0_chany_out_160_;
wire [0:0] cby_1__1__0_chany_out_161_;
wire [0:0] cby_1__1__0_chany_out_162_;
wire [0:0] cby_1__1__0_chany_out_163_;
wire [0:0] cby_1__1__0_chany_out_164_;
wire [0:0] cby_1__1__0_chany_out_165_;
wire [0:0] cby_1__1__0_chany_out_166_;
wire [0:0] cby_1__1__0_chany_out_167_;
wire [0:0] cby_1__1__0_chany_out_168_;
wire [0:0] cby_1__1__0_chany_out_169_;
wire [0:0] cby_1__1__0_chany_out_16_;
wire [0:0] cby_1__1__0_chany_out_170_;
wire [0:0] cby_1__1__0_chany_out_171_;
wire [0:0] cby_1__1__0_chany_out_172_;
wire [0:0] cby_1__1__0_chany_out_173_;
wire [0:0] cby_1__1__0_chany_out_174_;
wire [0:0] cby_1__1__0_chany_out_175_;
wire [0:0] cby_1__1__0_chany_out_176_;
wire [0:0] cby_1__1__0_chany_out_177_;
wire [0:0] cby_1__1__0_chany_out_178_;
wire [0:0] cby_1__1__0_chany_out_179_;
wire [0:0] cby_1__1__0_chany_out_17_;
wire [0:0] cby_1__1__0_chany_out_180_;
wire [0:0] cby_1__1__0_chany_out_181_;
wire [0:0] cby_1__1__0_chany_out_182_;
wire [0:0] cby_1__1__0_chany_out_183_;
wire [0:0] cby_1__1__0_chany_out_184_;
wire [0:0] cby_1__1__0_chany_out_185_;
wire [0:0] cby_1__1__0_chany_out_186_;
wire [0:0] cby_1__1__0_chany_out_187_;
wire [0:0] cby_1__1__0_chany_out_188_;
wire [0:0] cby_1__1__0_chany_out_189_;
wire [0:0] cby_1__1__0_chany_out_18_;
wire [0:0] cby_1__1__0_chany_out_190_;
wire [0:0] cby_1__1__0_chany_out_191_;
wire [0:0] cby_1__1__0_chany_out_192_;
wire [0:0] cby_1__1__0_chany_out_193_;
wire [0:0] cby_1__1__0_chany_out_194_;
wire [0:0] cby_1__1__0_chany_out_195_;
wire [0:0] cby_1__1__0_chany_out_196_;
wire [0:0] cby_1__1__0_chany_out_197_;
wire [0:0] cby_1__1__0_chany_out_198_;
wire [0:0] cby_1__1__0_chany_out_199_;
wire [0:0] cby_1__1__0_chany_out_19_;
wire [0:0] cby_1__1__0_chany_out_1_;
wire [0:0] cby_1__1__0_chany_out_20_;
wire [0:0] cby_1__1__0_chany_out_21_;
wire [0:0] cby_1__1__0_chany_out_22_;
wire [0:0] cby_1__1__0_chany_out_23_;
wire [0:0] cby_1__1__0_chany_out_24_;
wire [0:0] cby_1__1__0_chany_out_25_;
wire [0:0] cby_1__1__0_chany_out_26_;
wire [0:0] cby_1__1__0_chany_out_27_;
wire [0:0] cby_1__1__0_chany_out_28_;
wire [0:0] cby_1__1__0_chany_out_29_;
wire [0:0] cby_1__1__0_chany_out_2_;
wire [0:0] cby_1__1__0_chany_out_30_;
wire [0:0] cby_1__1__0_chany_out_31_;
wire [0:0] cby_1__1__0_chany_out_32_;
wire [0:0] cby_1__1__0_chany_out_33_;
wire [0:0] cby_1__1__0_chany_out_34_;
wire [0:0] cby_1__1__0_chany_out_35_;
wire [0:0] cby_1__1__0_chany_out_36_;
wire [0:0] cby_1__1__0_chany_out_37_;
wire [0:0] cby_1__1__0_chany_out_38_;
wire [0:0] cby_1__1__0_chany_out_39_;
wire [0:0] cby_1__1__0_chany_out_3_;
wire [0:0] cby_1__1__0_chany_out_40_;
wire [0:0] cby_1__1__0_chany_out_41_;
wire [0:0] cby_1__1__0_chany_out_42_;
wire [0:0] cby_1__1__0_chany_out_43_;
wire [0:0] cby_1__1__0_chany_out_44_;
wire [0:0] cby_1__1__0_chany_out_45_;
wire [0:0] cby_1__1__0_chany_out_46_;
wire [0:0] cby_1__1__0_chany_out_47_;
wire [0:0] cby_1__1__0_chany_out_48_;
wire [0:0] cby_1__1__0_chany_out_49_;
wire [0:0] cby_1__1__0_chany_out_4_;
wire [0:0] cby_1__1__0_chany_out_50_;
wire [0:0] cby_1__1__0_chany_out_51_;
wire [0:0] cby_1__1__0_chany_out_52_;
wire [0:0] cby_1__1__0_chany_out_53_;
wire [0:0] cby_1__1__0_chany_out_54_;
wire [0:0] cby_1__1__0_chany_out_55_;
wire [0:0] cby_1__1__0_chany_out_56_;
wire [0:0] cby_1__1__0_chany_out_57_;
wire [0:0] cby_1__1__0_chany_out_58_;
wire [0:0] cby_1__1__0_chany_out_59_;
wire [0:0] cby_1__1__0_chany_out_5_;
wire [0:0] cby_1__1__0_chany_out_60_;
wire [0:0] cby_1__1__0_chany_out_61_;
wire [0:0] cby_1__1__0_chany_out_62_;
wire [0:0] cby_1__1__0_chany_out_63_;
wire [0:0] cby_1__1__0_chany_out_64_;
wire [0:0] cby_1__1__0_chany_out_65_;
wire [0:0] cby_1__1__0_chany_out_66_;
wire [0:0] cby_1__1__0_chany_out_67_;
wire [0:0] cby_1__1__0_chany_out_68_;
wire [0:0] cby_1__1__0_chany_out_69_;
wire [0:0] cby_1__1__0_chany_out_6_;
wire [0:0] cby_1__1__0_chany_out_70_;
wire [0:0] cby_1__1__0_chany_out_71_;
wire [0:0] cby_1__1__0_chany_out_72_;
wire [0:0] cby_1__1__0_chany_out_73_;
wire [0:0] cby_1__1__0_chany_out_74_;
wire [0:0] cby_1__1__0_chany_out_75_;
wire [0:0] cby_1__1__0_chany_out_76_;
wire [0:0] cby_1__1__0_chany_out_77_;
wire [0:0] cby_1__1__0_chany_out_78_;
wire [0:0] cby_1__1__0_chany_out_79_;
wire [0:0] cby_1__1__0_chany_out_7_;
wire [0:0] cby_1__1__0_chany_out_80_;
wire [0:0] cby_1__1__0_chany_out_81_;
wire [0:0] cby_1__1__0_chany_out_82_;
wire [0:0] cby_1__1__0_chany_out_83_;
wire [0:0] cby_1__1__0_chany_out_84_;
wire [0:0] cby_1__1__0_chany_out_85_;
wire [0:0] cby_1__1__0_chany_out_86_;
wire [0:0] cby_1__1__0_chany_out_87_;
wire [0:0] cby_1__1__0_chany_out_88_;
wire [0:0] cby_1__1__0_chany_out_89_;
wire [0:0] cby_1__1__0_chany_out_8_;
wire [0:0] cby_1__1__0_chany_out_90_;
wire [0:0] cby_1__1__0_chany_out_91_;
wire [0:0] cby_1__1__0_chany_out_92_;
wire [0:0] cby_1__1__0_chany_out_93_;
wire [0:0] cby_1__1__0_chany_out_94_;
wire [0:0] cby_1__1__0_chany_out_95_;
wire [0:0] cby_1__1__0_chany_out_96_;
wire [0:0] cby_1__1__0_chany_out_97_;
wire [0:0] cby_1__1__0_chany_out_98_;
wire [0:0] cby_1__1__0_chany_out_99_;
wire [0:0] cby_1__1__0_chany_out_9_;
wire [0:0] cby_1__1__0_left_grid_pin_0_;
wire [0:0] cby_1__1__0_left_grid_pin_10_;
wire [0:0] cby_1__1__0_left_grid_pin_11_;
wire [0:0] cby_1__1__0_left_grid_pin_12_;
wire [0:0] cby_1__1__0_left_grid_pin_13_;
wire [0:0] cby_1__1__0_left_grid_pin_14_;
wire [0:0] cby_1__1__0_left_grid_pin_15_;
wire [0:0] cby_1__1__0_left_grid_pin_16_;
wire [0:0] cby_1__1__0_left_grid_pin_17_;
wire [0:0] cby_1__1__0_left_grid_pin_18_;
wire [0:0] cby_1__1__0_left_grid_pin_19_;
wire [0:0] cby_1__1__0_left_grid_pin_1_;
wire [0:0] cby_1__1__0_left_grid_pin_2_;
wire [0:0] cby_1__1__0_left_grid_pin_3_;
wire [0:0] cby_1__1__0_left_grid_pin_4_;
wire [0:0] cby_1__1__0_left_grid_pin_5_;
wire [0:0] cby_1__1__0_left_grid_pin_6_;
wire [0:0] cby_1__1__0_left_grid_pin_7_;
wire [0:0] cby_1__1__0_left_grid_pin_8_;
wire [0:0] cby_1__1__0_left_grid_pin_9_;
wire [0:0] cby_1__1__1_ccff_tail;
wire [0:0] cby_1__1__1_chany_out_0_;
wire [0:0] cby_1__1__1_chany_out_100_;
wire [0:0] cby_1__1__1_chany_out_101_;
wire [0:0] cby_1__1__1_chany_out_102_;
wire [0:0] cby_1__1__1_chany_out_103_;
wire [0:0] cby_1__1__1_chany_out_104_;
wire [0:0] cby_1__1__1_chany_out_105_;
wire [0:0] cby_1__1__1_chany_out_106_;
wire [0:0] cby_1__1__1_chany_out_107_;
wire [0:0] cby_1__1__1_chany_out_108_;
wire [0:0] cby_1__1__1_chany_out_109_;
wire [0:0] cby_1__1__1_chany_out_10_;
wire [0:0] cby_1__1__1_chany_out_110_;
wire [0:0] cby_1__1__1_chany_out_111_;
wire [0:0] cby_1__1__1_chany_out_112_;
wire [0:0] cby_1__1__1_chany_out_113_;
wire [0:0] cby_1__1__1_chany_out_114_;
wire [0:0] cby_1__1__1_chany_out_115_;
wire [0:0] cby_1__1__1_chany_out_116_;
wire [0:0] cby_1__1__1_chany_out_117_;
wire [0:0] cby_1__1__1_chany_out_118_;
wire [0:0] cby_1__1__1_chany_out_119_;
wire [0:0] cby_1__1__1_chany_out_11_;
wire [0:0] cby_1__1__1_chany_out_120_;
wire [0:0] cby_1__1__1_chany_out_121_;
wire [0:0] cby_1__1__1_chany_out_122_;
wire [0:0] cby_1__1__1_chany_out_123_;
wire [0:0] cby_1__1__1_chany_out_124_;
wire [0:0] cby_1__1__1_chany_out_125_;
wire [0:0] cby_1__1__1_chany_out_126_;
wire [0:0] cby_1__1__1_chany_out_127_;
wire [0:0] cby_1__1__1_chany_out_128_;
wire [0:0] cby_1__1__1_chany_out_129_;
wire [0:0] cby_1__1__1_chany_out_12_;
wire [0:0] cby_1__1__1_chany_out_130_;
wire [0:0] cby_1__1__1_chany_out_131_;
wire [0:0] cby_1__1__1_chany_out_132_;
wire [0:0] cby_1__1__1_chany_out_133_;
wire [0:0] cby_1__1__1_chany_out_134_;
wire [0:0] cby_1__1__1_chany_out_135_;
wire [0:0] cby_1__1__1_chany_out_136_;
wire [0:0] cby_1__1__1_chany_out_137_;
wire [0:0] cby_1__1__1_chany_out_138_;
wire [0:0] cby_1__1__1_chany_out_139_;
wire [0:0] cby_1__1__1_chany_out_13_;
wire [0:0] cby_1__1__1_chany_out_140_;
wire [0:0] cby_1__1__1_chany_out_141_;
wire [0:0] cby_1__1__1_chany_out_142_;
wire [0:0] cby_1__1__1_chany_out_143_;
wire [0:0] cby_1__1__1_chany_out_144_;
wire [0:0] cby_1__1__1_chany_out_145_;
wire [0:0] cby_1__1__1_chany_out_146_;
wire [0:0] cby_1__1__1_chany_out_147_;
wire [0:0] cby_1__1__1_chany_out_148_;
wire [0:0] cby_1__1__1_chany_out_149_;
wire [0:0] cby_1__1__1_chany_out_14_;
wire [0:0] cby_1__1__1_chany_out_150_;
wire [0:0] cby_1__1__1_chany_out_151_;
wire [0:0] cby_1__1__1_chany_out_152_;
wire [0:0] cby_1__1__1_chany_out_153_;
wire [0:0] cby_1__1__1_chany_out_154_;
wire [0:0] cby_1__1__1_chany_out_155_;
wire [0:0] cby_1__1__1_chany_out_156_;
wire [0:0] cby_1__1__1_chany_out_157_;
wire [0:0] cby_1__1__1_chany_out_158_;
wire [0:0] cby_1__1__1_chany_out_159_;
wire [0:0] cby_1__1__1_chany_out_15_;
wire [0:0] cby_1__1__1_chany_out_160_;
wire [0:0] cby_1__1__1_chany_out_161_;
wire [0:0] cby_1__1__1_chany_out_162_;
wire [0:0] cby_1__1__1_chany_out_163_;
wire [0:0] cby_1__1__1_chany_out_164_;
wire [0:0] cby_1__1__1_chany_out_165_;
wire [0:0] cby_1__1__1_chany_out_166_;
wire [0:0] cby_1__1__1_chany_out_167_;
wire [0:0] cby_1__1__1_chany_out_168_;
wire [0:0] cby_1__1__1_chany_out_169_;
wire [0:0] cby_1__1__1_chany_out_16_;
wire [0:0] cby_1__1__1_chany_out_170_;
wire [0:0] cby_1__1__1_chany_out_171_;
wire [0:0] cby_1__1__1_chany_out_172_;
wire [0:0] cby_1__1__1_chany_out_173_;
wire [0:0] cby_1__1__1_chany_out_174_;
wire [0:0] cby_1__1__1_chany_out_175_;
wire [0:0] cby_1__1__1_chany_out_176_;
wire [0:0] cby_1__1__1_chany_out_177_;
wire [0:0] cby_1__1__1_chany_out_178_;
wire [0:0] cby_1__1__1_chany_out_179_;
wire [0:0] cby_1__1__1_chany_out_17_;
wire [0:0] cby_1__1__1_chany_out_180_;
wire [0:0] cby_1__1__1_chany_out_181_;
wire [0:0] cby_1__1__1_chany_out_182_;
wire [0:0] cby_1__1__1_chany_out_183_;
wire [0:0] cby_1__1__1_chany_out_184_;
wire [0:0] cby_1__1__1_chany_out_185_;
wire [0:0] cby_1__1__1_chany_out_186_;
wire [0:0] cby_1__1__1_chany_out_187_;
wire [0:0] cby_1__1__1_chany_out_188_;
wire [0:0] cby_1__1__1_chany_out_189_;
wire [0:0] cby_1__1__1_chany_out_18_;
wire [0:0] cby_1__1__1_chany_out_190_;
wire [0:0] cby_1__1__1_chany_out_191_;
wire [0:0] cby_1__1__1_chany_out_192_;
wire [0:0] cby_1__1__1_chany_out_193_;
wire [0:0] cby_1__1__1_chany_out_194_;
wire [0:0] cby_1__1__1_chany_out_195_;
wire [0:0] cby_1__1__1_chany_out_196_;
wire [0:0] cby_1__1__1_chany_out_197_;
wire [0:0] cby_1__1__1_chany_out_198_;
wire [0:0] cby_1__1__1_chany_out_199_;
wire [0:0] cby_1__1__1_chany_out_19_;
wire [0:0] cby_1__1__1_chany_out_1_;
wire [0:0] cby_1__1__1_chany_out_20_;
wire [0:0] cby_1__1__1_chany_out_21_;
wire [0:0] cby_1__1__1_chany_out_22_;
wire [0:0] cby_1__1__1_chany_out_23_;
wire [0:0] cby_1__1__1_chany_out_24_;
wire [0:0] cby_1__1__1_chany_out_25_;
wire [0:0] cby_1__1__1_chany_out_26_;
wire [0:0] cby_1__1__1_chany_out_27_;
wire [0:0] cby_1__1__1_chany_out_28_;
wire [0:0] cby_1__1__1_chany_out_29_;
wire [0:0] cby_1__1__1_chany_out_2_;
wire [0:0] cby_1__1__1_chany_out_30_;
wire [0:0] cby_1__1__1_chany_out_31_;
wire [0:0] cby_1__1__1_chany_out_32_;
wire [0:0] cby_1__1__1_chany_out_33_;
wire [0:0] cby_1__1__1_chany_out_34_;
wire [0:0] cby_1__1__1_chany_out_35_;
wire [0:0] cby_1__1__1_chany_out_36_;
wire [0:0] cby_1__1__1_chany_out_37_;
wire [0:0] cby_1__1__1_chany_out_38_;
wire [0:0] cby_1__1__1_chany_out_39_;
wire [0:0] cby_1__1__1_chany_out_3_;
wire [0:0] cby_1__1__1_chany_out_40_;
wire [0:0] cby_1__1__1_chany_out_41_;
wire [0:0] cby_1__1__1_chany_out_42_;
wire [0:0] cby_1__1__1_chany_out_43_;
wire [0:0] cby_1__1__1_chany_out_44_;
wire [0:0] cby_1__1__1_chany_out_45_;
wire [0:0] cby_1__1__1_chany_out_46_;
wire [0:0] cby_1__1__1_chany_out_47_;
wire [0:0] cby_1__1__1_chany_out_48_;
wire [0:0] cby_1__1__1_chany_out_49_;
wire [0:0] cby_1__1__1_chany_out_4_;
wire [0:0] cby_1__1__1_chany_out_50_;
wire [0:0] cby_1__1__1_chany_out_51_;
wire [0:0] cby_1__1__1_chany_out_52_;
wire [0:0] cby_1__1__1_chany_out_53_;
wire [0:0] cby_1__1__1_chany_out_54_;
wire [0:0] cby_1__1__1_chany_out_55_;
wire [0:0] cby_1__1__1_chany_out_56_;
wire [0:0] cby_1__1__1_chany_out_57_;
wire [0:0] cby_1__1__1_chany_out_58_;
wire [0:0] cby_1__1__1_chany_out_59_;
wire [0:0] cby_1__1__1_chany_out_5_;
wire [0:0] cby_1__1__1_chany_out_60_;
wire [0:0] cby_1__1__1_chany_out_61_;
wire [0:0] cby_1__1__1_chany_out_62_;
wire [0:0] cby_1__1__1_chany_out_63_;
wire [0:0] cby_1__1__1_chany_out_64_;
wire [0:0] cby_1__1__1_chany_out_65_;
wire [0:0] cby_1__1__1_chany_out_66_;
wire [0:0] cby_1__1__1_chany_out_67_;
wire [0:0] cby_1__1__1_chany_out_68_;
wire [0:0] cby_1__1__1_chany_out_69_;
wire [0:0] cby_1__1__1_chany_out_6_;
wire [0:0] cby_1__1__1_chany_out_70_;
wire [0:0] cby_1__1__1_chany_out_71_;
wire [0:0] cby_1__1__1_chany_out_72_;
wire [0:0] cby_1__1__1_chany_out_73_;
wire [0:0] cby_1__1__1_chany_out_74_;
wire [0:0] cby_1__1__1_chany_out_75_;
wire [0:0] cby_1__1__1_chany_out_76_;
wire [0:0] cby_1__1__1_chany_out_77_;
wire [0:0] cby_1__1__1_chany_out_78_;
wire [0:0] cby_1__1__1_chany_out_79_;
wire [0:0] cby_1__1__1_chany_out_7_;
wire [0:0] cby_1__1__1_chany_out_80_;
wire [0:0] cby_1__1__1_chany_out_81_;
wire [0:0] cby_1__1__1_chany_out_82_;
wire [0:0] cby_1__1__1_chany_out_83_;
wire [0:0] cby_1__1__1_chany_out_84_;
wire [0:0] cby_1__1__1_chany_out_85_;
wire [0:0] cby_1__1__1_chany_out_86_;
wire [0:0] cby_1__1__1_chany_out_87_;
wire [0:0] cby_1__1__1_chany_out_88_;
wire [0:0] cby_1__1__1_chany_out_89_;
wire [0:0] cby_1__1__1_chany_out_8_;
wire [0:0] cby_1__1__1_chany_out_90_;
wire [0:0] cby_1__1__1_chany_out_91_;
wire [0:0] cby_1__1__1_chany_out_92_;
wire [0:0] cby_1__1__1_chany_out_93_;
wire [0:0] cby_1__1__1_chany_out_94_;
wire [0:0] cby_1__1__1_chany_out_95_;
wire [0:0] cby_1__1__1_chany_out_96_;
wire [0:0] cby_1__1__1_chany_out_97_;
wire [0:0] cby_1__1__1_chany_out_98_;
wire [0:0] cby_1__1__1_chany_out_99_;
wire [0:0] cby_1__1__1_chany_out_9_;
wire [0:0] cby_1__1__1_left_grid_pin_0_;
wire [0:0] cby_1__1__1_left_grid_pin_10_;
wire [0:0] cby_1__1__1_left_grid_pin_11_;
wire [0:0] cby_1__1__1_left_grid_pin_12_;
wire [0:0] cby_1__1__1_left_grid_pin_13_;
wire [0:0] cby_1__1__1_left_grid_pin_14_;
wire [0:0] cby_1__1__1_left_grid_pin_15_;
wire [0:0] cby_1__1__1_left_grid_pin_16_;
wire [0:0] cby_1__1__1_left_grid_pin_17_;
wire [0:0] cby_1__1__1_left_grid_pin_18_;
wire [0:0] cby_1__1__1_left_grid_pin_19_;
wire [0:0] cby_1__1__1_left_grid_pin_1_;
wire [0:0] cby_1__1__1_left_grid_pin_2_;
wire [0:0] cby_1__1__1_left_grid_pin_3_;
wire [0:0] cby_1__1__1_left_grid_pin_4_;
wire [0:0] cby_1__1__1_left_grid_pin_5_;
wire [0:0] cby_1__1__1_left_grid_pin_6_;
wire [0:0] cby_1__1__1_left_grid_pin_7_;
wire [0:0] cby_1__1__1_left_grid_pin_8_;
wire [0:0] cby_1__1__1_left_grid_pin_9_;
wire [0:0] cby_2__1__0_ccff_tail;
wire [0:0] cby_2__1__0_chany_out_0_;
wire [0:0] cby_2__1__0_chany_out_100_;
wire [0:0] cby_2__1__0_chany_out_101_;
wire [0:0] cby_2__1__0_chany_out_102_;
wire [0:0] cby_2__1__0_chany_out_103_;
wire [0:0] cby_2__1__0_chany_out_104_;
wire [0:0] cby_2__1__0_chany_out_105_;
wire [0:0] cby_2__1__0_chany_out_106_;
wire [0:0] cby_2__1__0_chany_out_107_;
wire [0:0] cby_2__1__0_chany_out_108_;
wire [0:0] cby_2__1__0_chany_out_109_;
wire [0:0] cby_2__1__0_chany_out_10_;
wire [0:0] cby_2__1__0_chany_out_110_;
wire [0:0] cby_2__1__0_chany_out_111_;
wire [0:0] cby_2__1__0_chany_out_112_;
wire [0:0] cby_2__1__0_chany_out_113_;
wire [0:0] cby_2__1__0_chany_out_114_;
wire [0:0] cby_2__1__0_chany_out_115_;
wire [0:0] cby_2__1__0_chany_out_116_;
wire [0:0] cby_2__1__0_chany_out_117_;
wire [0:0] cby_2__1__0_chany_out_118_;
wire [0:0] cby_2__1__0_chany_out_119_;
wire [0:0] cby_2__1__0_chany_out_11_;
wire [0:0] cby_2__1__0_chany_out_120_;
wire [0:0] cby_2__1__0_chany_out_121_;
wire [0:0] cby_2__1__0_chany_out_122_;
wire [0:0] cby_2__1__0_chany_out_123_;
wire [0:0] cby_2__1__0_chany_out_124_;
wire [0:0] cby_2__1__0_chany_out_125_;
wire [0:0] cby_2__1__0_chany_out_126_;
wire [0:0] cby_2__1__0_chany_out_127_;
wire [0:0] cby_2__1__0_chany_out_128_;
wire [0:0] cby_2__1__0_chany_out_129_;
wire [0:0] cby_2__1__0_chany_out_12_;
wire [0:0] cby_2__1__0_chany_out_130_;
wire [0:0] cby_2__1__0_chany_out_131_;
wire [0:0] cby_2__1__0_chany_out_132_;
wire [0:0] cby_2__1__0_chany_out_133_;
wire [0:0] cby_2__1__0_chany_out_134_;
wire [0:0] cby_2__1__0_chany_out_135_;
wire [0:0] cby_2__1__0_chany_out_136_;
wire [0:0] cby_2__1__0_chany_out_137_;
wire [0:0] cby_2__1__0_chany_out_138_;
wire [0:0] cby_2__1__0_chany_out_139_;
wire [0:0] cby_2__1__0_chany_out_13_;
wire [0:0] cby_2__1__0_chany_out_140_;
wire [0:0] cby_2__1__0_chany_out_141_;
wire [0:0] cby_2__1__0_chany_out_142_;
wire [0:0] cby_2__1__0_chany_out_143_;
wire [0:0] cby_2__1__0_chany_out_144_;
wire [0:0] cby_2__1__0_chany_out_145_;
wire [0:0] cby_2__1__0_chany_out_146_;
wire [0:0] cby_2__1__0_chany_out_147_;
wire [0:0] cby_2__1__0_chany_out_148_;
wire [0:0] cby_2__1__0_chany_out_149_;
wire [0:0] cby_2__1__0_chany_out_14_;
wire [0:0] cby_2__1__0_chany_out_150_;
wire [0:0] cby_2__1__0_chany_out_151_;
wire [0:0] cby_2__1__0_chany_out_152_;
wire [0:0] cby_2__1__0_chany_out_153_;
wire [0:0] cby_2__1__0_chany_out_154_;
wire [0:0] cby_2__1__0_chany_out_155_;
wire [0:0] cby_2__1__0_chany_out_156_;
wire [0:0] cby_2__1__0_chany_out_157_;
wire [0:0] cby_2__1__0_chany_out_158_;
wire [0:0] cby_2__1__0_chany_out_159_;
wire [0:0] cby_2__1__0_chany_out_15_;
wire [0:0] cby_2__1__0_chany_out_160_;
wire [0:0] cby_2__1__0_chany_out_161_;
wire [0:0] cby_2__1__0_chany_out_162_;
wire [0:0] cby_2__1__0_chany_out_163_;
wire [0:0] cby_2__1__0_chany_out_164_;
wire [0:0] cby_2__1__0_chany_out_165_;
wire [0:0] cby_2__1__0_chany_out_166_;
wire [0:0] cby_2__1__0_chany_out_167_;
wire [0:0] cby_2__1__0_chany_out_168_;
wire [0:0] cby_2__1__0_chany_out_169_;
wire [0:0] cby_2__1__0_chany_out_16_;
wire [0:0] cby_2__1__0_chany_out_170_;
wire [0:0] cby_2__1__0_chany_out_171_;
wire [0:0] cby_2__1__0_chany_out_172_;
wire [0:0] cby_2__1__0_chany_out_173_;
wire [0:0] cby_2__1__0_chany_out_174_;
wire [0:0] cby_2__1__0_chany_out_175_;
wire [0:0] cby_2__1__0_chany_out_176_;
wire [0:0] cby_2__1__0_chany_out_177_;
wire [0:0] cby_2__1__0_chany_out_178_;
wire [0:0] cby_2__1__0_chany_out_179_;
wire [0:0] cby_2__1__0_chany_out_17_;
wire [0:0] cby_2__1__0_chany_out_180_;
wire [0:0] cby_2__1__0_chany_out_181_;
wire [0:0] cby_2__1__0_chany_out_182_;
wire [0:0] cby_2__1__0_chany_out_183_;
wire [0:0] cby_2__1__0_chany_out_184_;
wire [0:0] cby_2__1__0_chany_out_185_;
wire [0:0] cby_2__1__0_chany_out_186_;
wire [0:0] cby_2__1__0_chany_out_187_;
wire [0:0] cby_2__1__0_chany_out_188_;
wire [0:0] cby_2__1__0_chany_out_189_;
wire [0:0] cby_2__1__0_chany_out_18_;
wire [0:0] cby_2__1__0_chany_out_190_;
wire [0:0] cby_2__1__0_chany_out_191_;
wire [0:0] cby_2__1__0_chany_out_192_;
wire [0:0] cby_2__1__0_chany_out_193_;
wire [0:0] cby_2__1__0_chany_out_194_;
wire [0:0] cby_2__1__0_chany_out_195_;
wire [0:0] cby_2__1__0_chany_out_196_;
wire [0:0] cby_2__1__0_chany_out_197_;
wire [0:0] cby_2__1__0_chany_out_198_;
wire [0:0] cby_2__1__0_chany_out_199_;
wire [0:0] cby_2__1__0_chany_out_19_;
wire [0:0] cby_2__1__0_chany_out_1_;
wire [0:0] cby_2__1__0_chany_out_20_;
wire [0:0] cby_2__1__0_chany_out_21_;
wire [0:0] cby_2__1__0_chany_out_22_;
wire [0:0] cby_2__1__0_chany_out_23_;
wire [0:0] cby_2__1__0_chany_out_24_;
wire [0:0] cby_2__1__0_chany_out_25_;
wire [0:0] cby_2__1__0_chany_out_26_;
wire [0:0] cby_2__1__0_chany_out_27_;
wire [0:0] cby_2__1__0_chany_out_28_;
wire [0:0] cby_2__1__0_chany_out_29_;
wire [0:0] cby_2__1__0_chany_out_2_;
wire [0:0] cby_2__1__0_chany_out_30_;
wire [0:0] cby_2__1__0_chany_out_31_;
wire [0:0] cby_2__1__0_chany_out_32_;
wire [0:0] cby_2__1__0_chany_out_33_;
wire [0:0] cby_2__1__0_chany_out_34_;
wire [0:0] cby_2__1__0_chany_out_35_;
wire [0:0] cby_2__1__0_chany_out_36_;
wire [0:0] cby_2__1__0_chany_out_37_;
wire [0:0] cby_2__1__0_chany_out_38_;
wire [0:0] cby_2__1__0_chany_out_39_;
wire [0:0] cby_2__1__0_chany_out_3_;
wire [0:0] cby_2__1__0_chany_out_40_;
wire [0:0] cby_2__1__0_chany_out_41_;
wire [0:0] cby_2__1__0_chany_out_42_;
wire [0:0] cby_2__1__0_chany_out_43_;
wire [0:0] cby_2__1__0_chany_out_44_;
wire [0:0] cby_2__1__0_chany_out_45_;
wire [0:0] cby_2__1__0_chany_out_46_;
wire [0:0] cby_2__1__0_chany_out_47_;
wire [0:0] cby_2__1__0_chany_out_48_;
wire [0:0] cby_2__1__0_chany_out_49_;
wire [0:0] cby_2__1__0_chany_out_4_;
wire [0:0] cby_2__1__0_chany_out_50_;
wire [0:0] cby_2__1__0_chany_out_51_;
wire [0:0] cby_2__1__0_chany_out_52_;
wire [0:0] cby_2__1__0_chany_out_53_;
wire [0:0] cby_2__1__0_chany_out_54_;
wire [0:0] cby_2__1__0_chany_out_55_;
wire [0:0] cby_2__1__0_chany_out_56_;
wire [0:0] cby_2__1__0_chany_out_57_;
wire [0:0] cby_2__1__0_chany_out_58_;
wire [0:0] cby_2__1__0_chany_out_59_;
wire [0:0] cby_2__1__0_chany_out_5_;
wire [0:0] cby_2__1__0_chany_out_60_;
wire [0:0] cby_2__1__0_chany_out_61_;
wire [0:0] cby_2__1__0_chany_out_62_;
wire [0:0] cby_2__1__0_chany_out_63_;
wire [0:0] cby_2__1__0_chany_out_64_;
wire [0:0] cby_2__1__0_chany_out_65_;
wire [0:0] cby_2__1__0_chany_out_66_;
wire [0:0] cby_2__1__0_chany_out_67_;
wire [0:0] cby_2__1__0_chany_out_68_;
wire [0:0] cby_2__1__0_chany_out_69_;
wire [0:0] cby_2__1__0_chany_out_6_;
wire [0:0] cby_2__1__0_chany_out_70_;
wire [0:0] cby_2__1__0_chany_out_71_;
wire [0:0] cby_2__1__0_chany_out_72_;
wire [0:0] cby_2__1__0_chany_out_73_;
wire [0:0] cby_2__1__0_chany_out_74_;
wire [0:0] cby_2__1__0_chany_out_75_;
wire [0:0] cby_2__1__0_chany_out_76_;
wire [0:0] cby_2__1__0_chany_out_77_;
wire [0:0] cby_2__1__0_chany_out_78_;
wire [0:0] cby_2__1__0_chany_out_79_;
wire [0:0] cby_2__1__0_chany_out_7_;
wire [0:0] cby_2__1__0_chany_out_80_;
wire [0:0] cby_2__1__0_chany_out_81_;
wire [0:0] cby_2__1__0_chany_out_82_;
wire [0:0] cby_2__1__0_chany_out_83_;
wire [0:0] cby_2__1__0_chany_out_84_;
wire [0:0] cby_2__1__0_chany_out_85_;
wire [0:0] cby_2__1__0_chany_out_86_;
wire [0:0] cby_2__1__0_chany_out_87_;
wire [0:0] cby_2__1__0_chany_out_88_;
wire [0:0] cby_2__1__0_chany_out_89_;
wire [0:0] cby_2__1__0_chany_out_8_;
wire [0:0] cby_2__1__0_chany_out_90_;
wire [0:0] cby_2__1__0_chany_out_91_;
wire [0:0] cby_2__1__0_chany_out_92_;
wire [0:0] cby_2__1__0_chany_out_93_;
wire [0:0] cby_2__1__0_chany_out_94_;
wire [0:0] cby_2__1__0_chany_out_95_;
wire [0:0] cby_2__1__0_chany_out_96_;
wire [0:0] cby_2__1__0_chany_out_97_;
wire [0:0] cby_2__1__0_chany_out_98_;
wire [0:0] cby_2__1__0_chany_out_99_;
wire [0:0] cby_2__1__0_chany_out_9_;
wire [0:0] cby_2__1__0_left_grid_pin_0_;
wire [0:0] cby_2__1__0_left_grid_pin_10_;
wire [0:0] cby_2__1__0_left_grid_pin_11_;
wire [0:0] cby_2__1__0_left_grid_pin_12_;
wire [0:0] cby_2__1__0_left_grid_pin_13_;
wire [0:0] cby_2__1__0_left_grid_pin_14_;
wire [0:0] cby_2__1__0_left_grid_pin_15_;
wire [0:0] cby_2__1__0_left_grid_pin_16_;
wire [0:0] cby_2__1__0_left_grid_pin_17_;
wire [0:0] cby_2__1__0_left_grid_pin_18_;
wire [0:0] cby_2__1__0_left_grid_pin_19_;
wire [0:0] cby_2__1__0_left_grid_pin_1_;
wire [0:0] cby_2__1__0_left_grid_pin_2_;
wire [0:0] cby_2__1__0_left_grid_pin_3_;
wire [0:0] cby_2__1__0_left_grid_pin_4_;
wire [0:0] cby_2__1__0_left_grid_pin_5_;
wire [0:0] cby_2__1__0_left_grid_pin_6_;
wire [0:0] cby_2__1__0_left_grid_pin_7_;
wire [0:0] cby_2__1__0_left_grid_pin_8_;
wire [0:0] cby_2__1__0_left_grid_pin_9_;
wire [0:0] cby_2__1__0_right_grid_pin_0_;
wire [0:0] cby_2__1__1_ccff_tail;
wire [0:0] cby_2__1__1_chany_out_0_;
wire [0:0] cby_2__1__1_chany_out_100_;
wire [0:0] cby_2__1__1_chany_out_101_;
wire [0:0] cby_2__1__1_chany_out_102_;
wire [0:0] cby_2__1__1_chany_out_103_;
wire [0:0] cby_2__1__1_chany_out_104_;
wire [0:0] cby_2__1__1_chany_out_105_;
wire [0:0] cby_2__1__1_chany_out_106_;
wire [0:0] cby_2__1__1_chany_out_107_;
wire [0:0] cby_2__1__1_chany_out_108_;
wire [0:0] cby_2__1__1_chany_out_109_;
wire [0:0] cby_2__1__1_chany_out_10_;
wire [0:0] cby_2__1__1_chany_out_110_;
wire [0:0] cby_2__1__1_chany_out_111_;
wire [0:0] cby_2__1__1_chany_out_112_;
wire [0:0] cby_2__1__1_chany_out_113_;
wire [0:0] cby_2__1__1_chany_out_114_;
wire [0:0] cby_2__1__1_chany_out_115_;
wire [0:0] cby_2__1__1_chany_out_116_;
wire [0:0] cby_2__1__1_chany_out_117_;
wire [0:0] cby_2__1__1_chany_out_118_;
wire [0:0] cby_2__1__1_chany_out_119_;
wire [0:0] cby_2__1__1_chany_out_11_;
wire [0:0] cby_2__1__1_chany_out_120_;
wire [0:0] cby_2__1__1_chany_out_121_;
wire [0:0] cby_2__1__1_chany_out_122_;
wire [0:0] cby_2__1__1_chany_out_123_;
wire [0:0] cby_2__1__1_chany_out_124_;
wire [0:0] cby_2__1__1_chany_out_125_;
wire [0:0] cby_2__1__1_chany_out_126_;
wire [0:0] cby_2__1__1_chany_out_127_;
wire [0:0] cby_2__1__1_chany_out_128_;
wire [0:0] cby_2__1__1_chany_out_129_;
wire [0:0] cby_2__1__1_chany_out_12_;
wire [0:0] cby_2__1__1_chany_out_130_;
wire [0:0] cby_2__1__1_chany_out_131_;
wire [0:0] cby_2__1__1_chany_out_132_;
wire [0:0] cby_2__1__1_chany_out_133_;
wire [0:0] cby_2__1__1_chany_out_134_;
wire [0:0] cby_2__1__1_chany_out_135_;
wire [0:0] cby_2__1__1_chany_out_136_;
wire [0:0] cby_2__1__1_chany_out_137_;
wire [0:0] cby_2__1__1_chany_out_138_;
wire [0:0] cby_2__1__1_chany_out_139_;
wire [0:0] cby_2__1__1_chany_out_13_;
wire [0:0] cby_2__1__1_chany_out_140_;
wire [0:0] cby_2__1__1_chany_out_141_;
wire [0:0] cby_2__1__1_chany_out_142_;
wire [0:0] cby_2__1__1_chany_out_143_;
wire [0:0] cby_2__1__1_chany_out_144_;
wire [0:0] cby_2__1__1_chany_out_145_;
wire [0:0] cby_2__1__1_chany_out_146_;
wire [0:0] cby_2__1__1_chany_out_147_;
wire [0:0] cby_2__1__1_chany_out_148_;
wire [0:0] cby_2__1__1_chany_out_149_;
wire [0:0] cby_2__1__1_chany_out_14_;
wire [0:0] cby_2__1__1_chany_out_150_;
wire [0:0] cby_2__1__1_chany_out_151_;
wire [0:0] cby_2__1__1_chany_out_152_;
wire [0:0] cby_2__1__1_chany_out_153_;
wire [0:0] cby_2__1__1_chany_out_154_;
wire [0:0] cby_2__1__1_chany_out_155_;
wire [0:0] cby_2__1__1_chany_out_156_;
wire [0:0] cby_2__1__1_chany_out_157_;
wire [0:0] cby_2__1__1_chany_out_158_;
wire [0:0] cby_2__1__1_chany_out_159_;
wire [0:0] cby_2__1__1_chany_out_15_;
wire [0:0] cby_2__1__1_chany_out_160_;
wire [0:0] cby_2__1__1_chany_out_161_;
wire [0:0] cby_2__1__1_chany_out_162_;
wire [0:0] cby_2__1__1_chany_out_163_;
wire [0:0] cby_2__1__1_chany_out_164_;
wire [0:0] cby_2__1__1_chany_out_165_;
wire [0:0] cby_2__1__1_chany_out_166_;
wire [0:0] cby_2__1__1_chany_out_167_;
wire [0:0] cby_2__1__1_chany_out_168_;
wire [0:0] cby_2__1__1_chany_out_169_;
wire [0:0] cby_2__1__1_chany_out_16_;
wire [0:0] cby_2__1__1_chany_out_170_;
wire [0:0] cby_2__1__1_chany_out_171_;
wire [0:0] cby_2__1__1_chany_out_172_;
wire [0:0] cby_2__1__1_chany_out_173_;
wire [0:0] cby_2__1__1_chany_out_174_;
wire [0:0] cby_2__1__1_chany_out_175_;
wire [0:0] cby_2__1__1_chany_out_176_;
wire [0:0] cby_2__1__1_chany_out_177_;
wire [0:0] cby_2__1__1_chany_out_178_;
wire [0:0] cby_2__1__1_chany_out_179_;
wire [0:0] cby_2__1__1_chany_out_17_;
wire [0:0] cby_2__1__1_chany_out_180_;
wire [0:0] cby_2__1__1_chany_out_181_;
wire [0:0] cby_2__1__1_chany_out_182_;
wire [0:0] cby_2__1__1_chany_out_183_;
wire [0:0] cby_2__1__1_chany_out_184_;
wire [0:0] cby_2__1__1_chany_out_185_;
wire [0:0] cby_2__1__1_chany_out_186_;
wire [0:0] cby_2__1__1_chany_out_187_;
wire [0:0] cby_2__1__1_chany_out_188_;
wire [0:0] cby_2__1__1_chany_out_189_;
wire [0:0] cby_2__1__1_chany_out_18_;
wire [0:0] cby_2__1__1_chany_out_190_;
wire [0:0] cby_2__1__1_chany_out_191_;
wire [0:0] cby_2__1__1_chany_out_192_;
wire [0:0] cby_2__1__1_chany_out_193_;
wire [0:0] cby_2__1__1_chany_out_194_;
wire [0:0] cby_2__1__1_chany_out_195_;
wire [0:0] cby_2__1__1_chany_out_196_;
wire [0:0] cby_2__1__1_chany_out_197_;
wire [0:0] cby_2__1__1_chany_out_198_;
wire [0:0] cby_2__1__1_chany_out_199_;
wire [0:0] cby_2__1__1_chany_out_19_;
wire [0:0] cby_2__1__1_chany_out_1_;
wire [0:0] cby_2__1__1_chany_out_20_;
wire [0:0] cby_2__1__1_chany_out_21_;
wire [0:0] cby_2__1__1_chany_out_22_;
wire [0:0] cby_2__1__1_chany_out_23_;
wire [0:0] cby_2__1__1_chany_out_24_;
wire [0:0] cby_2__1__1_chany_out_25_;
wire [0:0] cby_2__1__1_chany_out_26_;
wire [0:0] cby_2__1__1_chany_out_27_;
wire [0:0] cby_2__1__1_chany_out_28_;
wire [0:0] cby_2__1__1_chany_out_29_;
wire [0:0] cby_2__1__1_chany_out_2_;
wire [0:0] cby_2__1__1_chany_out_30_;
wire [0:0] cby_2__1__1_chany_out_31_;
wire [0:0] cby_2__1__1_chany_out_32_;
wire [0:0] cby_2__1__1_chany_out_33_;
wire [0:0] cby_2__1__1_chany_out_34_;
wire [0:0] cby_2__1__1_chany_out_35_;
wire [0:0] cby_2__1__1_chany_out_36_;
wire [0:0] cby_2__1__1_chany_out_37_;
wire [0:0] cby_2__1__1_chany_out_38_;
wire [0:0] cby_2__1__1_chany_out_39_;
wire [0:0] cby_2__1__1_chany_out_3_;
wire [0:0] cby_2__1__1_chany_out_40_;
wire [0:0] cby_2__1__1_chany_out_41_;
wire [0:0] cby_2__1__1_chany_out_42_;
wire [0:0] cby_2__1__1_chany_out_43_;
wire [0:0] cby_2__1__1_chany_out_44_;
wire [0:0] cby_2__1__1_chany_out_45_;
wire [0:0] cby_2__1__1_chany_out_46_;
wire [0:0] cby_2__1__1_chany_out_47_;
wire [0:0] cby_2__1__1_chany_out_48_;
wire [0:0] cby_2__1__1_chany_out_49_;
wire [0:0] cby_2__1__1_chany_out_4_;
wire [0:0] cby_2__1__1_chany_out_50_;
wire [0:0] cby_2__1__1_chany_out_51_;
wire [0:0] cby_2__1__1_chany_out_52_;
wire [0:0] cby_2__1__1_chany_out_53_;
wire [0:0] cby_2__1__1_chany_out_54_;
wire [0:0] cby_2__1__1_chany_out_55_;
wire [0:0] cby_2__1__1_chany_out_56_;
wire [0:0] cby_2__1__1_chany_out_57_;
wire [0:0] cby_2__1__1_chany_out_58_;
wire [0:0] cby_2__1__1_chany_out_59_;
wire [0:0] cby_2__1__1_chany_out_5_;
wire [0:0] cby_2__1__1_chany_out_60_;
wire [0:0] cby_2__1__1_chany_out_61_;
wire [0:0] cby_2__1__1_chany_out_62_;
wire [0:0] cby_2__1__1_chany_out_63_;
wire [0:0] cby_2__1__1_chany_out_64_;
wire [0:0] cby_2__1__1_chany_out_65_;
wire [0:0] cby_2__1__1_chany_out_66_;
wire [0:0] cby_2__1__1_chany_out_67_;
wire [0:0] cby_2__1__1_chany_out_68_;
wire [0:0] cby_2__1__1_chany_out_69_;
wire [0:0] cby_2__1__1_chany_out_6_;
wire [0:0] cby_2__1__1_chany_out_70_;
wire [0:0] cby_2__1__1_chany_out_71_;
wire [0:0] cby_2__1__1_chany_out_72_;
wire [0:0] cby_2__1__1_chany_out_73_;
wire [0:0] cby_2__1__1_chany_out_74_;
wire [0:0] cby_2__1__1_chany_out_75_;
wire [0:0] cby_2__1__1_chany_out_76_;
wire [0:0] cby_2__1__1_chany_out_77_;
wire [0:0] cby_2__1__1_chany_out_78_;
wire [0:0] cby_2__1__1_chany_out_79_;
wire [0:0] cby_2__1__1_chany_out_7_;
wire [0:0] cby_2__1__1_chany_out_80_;
wire [0:0] cby_2__1__1_chany_out_81_;
wire [0:0] cby_2__1__1_chany_out_82_;
wire [0:0] cby_2__1__1_chany_out_83_;
wire [0:0] cby_2__1__1_chany_out_84_;
wire [0:0] cby_2__1__1_chany_out_85_;
wire [0:0] cby_2__1__1_chany_out_86_;
wire [0:0] cby_2__1__1_chany_out_87_;
wire [0:0] cby_2__1__1_chany_out_88_;
wire [0:0] cby_2__1__1_chany_out_89_;
wire [0:0] cby_2__1__1_chany_out_8_;
wire [0:0] cby_2__1__1_chany_out_90_;
wire [0:0] cby_2__1__1_chany_out_91_;
wire [0:0] cby_2__1__1_chany_out_92_;
wire [0:0] cby_2__1__1_chany_out_93_;
wire [0:0] cby_2__1__1_chany_out_94_;
wire [0:0] cby_2__1__1_chany_out_95_;
wire [0:0] cby_2__1__1_chany_out_96_;
wire [0:0] cby_2__1__1_chany_out_97_;
wire [0:0] cby_2__1__1_chany_out_98_;
wire [0:0] cby_2__1__1_chany_out_99_;
wire [0:0] cby_2__1__1_chany_out_9_;
wire [0:0] cby_2__1__1_left_grid_pin_0_;
wire [0:0] cby_2__1__1_left_grid_pin_10_;
wire [0:0] cby_2__1__1_left_grid_pin_11_;
wire [0:0] cby_2__1__1_left_grid_pin_12_;
wire [0:0] cby_2__1__1_left_grid_pin_13_;
wire [0:0] cby_2__1__1_left_grid_pin_14_;
wire [0:0] cby_2__1__1_left_grid_pin_15_;
wire [0:0] cby_2__1__1_left_grid_pin_16_;
wire [0:0] cby_2__1__1_left_grid_pin_17_;
wire [0:0] cby_2__1__1_left_grid_pin_18_;
wire [0:0] cby_2__1__1_left_grid_pin_19_;
wire [0:0] cby_2__1__1_left_grid_pin_1_;
wire [0:0] cby_2__1__1_left_grid_pin_2_;
wire [0:0] cby_2__1__1_left_grid_pin_3_;
wire [0:0] cby_2__1__1_left_grid_pin_4_;
wire [0:0] cby_2__1__1_left_grid_pin_5_;
wire [0:0] cby_2__1__1_left_grid_pin_6_;
wire [0:0] cby_2__1__1_left_grid_pin_7_;
wire [0:0] cby_2__1__1_left_grid_pin_8_;
wire [0:0] cby_2__1__1_left_grid_pin_9_;
wire [0:0] cby_2__1__1_right_grid_pin_0_;
wire [0:0] direct_interc_0_out;
wire [0:0] direct_interc_1_out;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_54_lower;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_54_upper;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_55_lower;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_55_upper;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_56_lower;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_56_upper;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_57_lower;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_57_upper;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_58_lower;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_58_upper;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_59_lower;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_59_upper;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_60_lower;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_60_upper;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_61_lower;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_61_upper;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_62_lower;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_62_upper;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_63_lower;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_63_upper;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_66_lower;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_66_upper;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_67_lower;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_67_upper;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_50_lower;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_50_upper;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_51_lower;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_51_upper;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_52_lower;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_52_upper;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_53_lower;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_53_upper;
wire [0:0] grid_clb_1_2_undriven_bottom_width_0_height_0__pin_64_;
wire [0:0] grid_clb_1_2_undriven_bottom_width_0_height_0__pin_65_;
wire [0:0] grid_clb_1_2_undriven_top_width_0_height_0__pin_40_;
wire [0:0] grid_clb_1_2_undriven_top_width_0_height_0__pin_41_;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_54_lower;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_54_upper;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_55_lower;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_55_upper;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_56_lower;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_56_upper;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_57_lower;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_57_upper;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_58_lower;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_58_upper;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_59_lower;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_59_upper;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_60_lower;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_60_upper;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_61_lower;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_61_upper;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_62_lower;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_62_upper;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_63_lower;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_63_upper;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_66_lower;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_66_upper;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_67_lower;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_67_upper;
wire [0:0] grid_clb_1_ccff_tail;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_50_lower;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_50_upper;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_51_lower;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_51_upper;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_52_lower;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_52_upper;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_53_lower;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_53_upper;
wire [0:0] grid_clb_2_1_undriven_bottom_width_0_height_0__pin_64_;
wire [0:0] grid_clb_2_1_undriven_bottom_width_0_height_0__pin_65_;
wire [0:0] grid_clb_2_2_undriven_top_width_0_height_0__pin_40_;
wire [0:0] grid_clb_2_2_undriven_top_width_0_height_0__pin_41_;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_54_lower;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_54_upper;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_55_lower;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_55_upper;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_56_lower;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_56_upper;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_57_lower;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_57_upper;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_58_lower;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_58_upper;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_59_lower;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_59_upper;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_60_lower;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_60_upper;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_61_lower;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_61_upper;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_62_lower;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_62_upper;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_63_lower;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_63_upper;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_64_;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_65_;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_66_lower;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_66_upper;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_67_lower;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_67_upper;
wire [0:0] grid_clb_2_ccff_tail;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_50_lower;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_50_upper;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_51_lower;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_51_upper;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_52_lower;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_52_upper;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_53_lower;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_53_upper;
wire [0:0] grid_clb_spypad_0_bottom_width_0_height_0__pin_54_lower;
wire [0:0] grid_clb_spypad_0_bottom_width_0_height_0__pin_54_upper;
wire [0:0] grid_clb_spypad_0_bottom_width_0_height_0__pin_55_lower;
wire [0:0] grid_clb_spypad_0_bottom_width_0_height_0__pin_55_upper;
wire [0:0] grid_clb_spypad_0_bottom_width_0_height_0__pin_56_lower;
wire [0:0] grid_clb_spypad_0_bottom_width_0_height_0__pin_56_upper;
wire [0:0] grid_clb_spypad_0_bottom_width_0_height_0__pin_57_lower;
wire [0:0] grid_clb_spypad_0_bottom_width_0_height_0__pin_57_upper;
wire [0:0] grid_clb_spypad_0_bottom_width_0_height_0__pin_58_lower;
wire [0:0] grid_clb_spypad_0_bottom_width_0_height_0__pin_58_upper;
wire [0:0] grid_clb_spypad_0_bottom_width_0_height_0__pin_59_lower;
wire [0:0] grid_clb_spypad_0_bottom_width_0_height_0__pin_59_upper;
wire [0:0] grid_clb_spypad_0_bottom_width_0_height_0__pin_60_lower;
wire [0:0] grid_clb_spypad_0_bottom_width_0_height_0__pin_60_upper;
wire [0:0] grid_clb_spypad_0_bottom_width_0_height_0__pin_61_lower;
wire [0:0] grid_clb_spypad_0_bottom_width_0_height_0__pin_61_upper;
wire [0:0] grid_clb_spypad_0_bottom_width_0_height_0__pin_62_lower;
wire [0:0] grid_clb_spypad_0_bottom_width_0_height_0__pin_62_upper;
wire [0:0] grid_clb_spypad_0_bottom_width_0_height_0__pin_63_lower;
wire [0:0] grid_clb_spypad_0_bottom_width_0_height_0__pin_63_upper;
wire [0:0] grid_clb_spypad_0_bottom_width_0_height_0__pin_66_lower;
wire [0:0] grid_clb_spypad_0_bottom_width_0_height_0__pin_66_upper;
wire [0:0] grid_clb_spypad_0_bottom_width_0_height_0__pin_67_lower;
wire [0:0] grid_clb_spypad_0_bottom_width_0_height_0__pin_67_upper;
wire [0:0] grid_clb_spypad_0_ccff_tail;
wire [0:0] grid_clb_spypad_0_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_spypad_0_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_spypad_0_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_spypad_0_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_spypad_0_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_spypad_0_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_spypad_0_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_spypad_0_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_spypad_0_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_spypad_0_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_spypad_0_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_spypad_0_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_spypad_0_right_width_0_height_0__pin_50_lower;
wire [0:0] grid_clb_spypad_0_right_width_0_height_0__pin_50_upper;
wire [0:0] grid_clb_spypad_0_right_width_0_height_0__pin_51_lower;
wire [0:0] grid_clb_spypad_0_right_width_0_height_0__pin_51_upper;
wire [0:0] grid_clb_spypad_0_right_width_0_height_0__pin_52_lower;
wire [0:0] grid_clb_spypad_0_right_width_0_height_0__pin_52_upper;
wire [0:0] grid_clb_spypad_0_right_width_0_height_0__pin_53_lower;
wire [0:0] grid_clb_spypad_0_right_width_0_height_0__pin_53_upper;
wire [0:0] grid_clb_1_1_undriven_bottom_width_0_height_0__pin_64_;
wire [0:0] grid_clb_1_1_undriven_bottom_width_0_height_0__pin_65_;
wire [0:0] grid_clb_1_1_undriven_top_width_0_height_0__pin_40_;
wire [0:0] grid_clb_1_1_undriven_top_width_0_height_0__pin_41_;
wire [0:0] grid_clb_1_1_undriven_top_width_0_height_0__pin_68_;
wire [0:0] grid_io_bottom_0_ccff_tail;
wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_bottom_1_ccff_tail;
wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_left_0_ccff_tail;
wire [0:0] grid_io_left_0_right_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_left_0_right_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_left_1_ccff_tail;
wire [0:0] grid_io_left_1_right_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_left_1_right_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_right_0_ccff_tail;
wire [0:0] grid_io_right_0_left_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_right_0_left_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_right_1_ccff_tail;
wire [0:0] grid_io_right_1_left_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_right_1_left_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_top_0_bottom_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_top_0_bottom_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_top_0_ccff_tail;
wire [0:0] grid_io_top_1_bottom_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_top_1_bottom_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_top_1_ccff_tail;
wire [0:0] sb_0__0__0_ccff_tail;
wire [0:0] sb_0__0__0_chanx_right_out_0_;
wire [0:0] sb_0__0__0_chanx_right_out_100_;
wire [0:0] sb_0__0__0_chanx_right_out_102_;
wire [0:0] sb_0__0__0_chanx_right_out_104_;
wire [0:0] sb_0__0__0_chanx_right_out_106_;
wire [0:0] sb_0__0__0_chanx_right_out_108_;
wire [0:0] sb_0__0__0_chanx_right_out_10_;
wire [0:0] sb_0__0__0_chanx_right_out_110_;
wire [0:0] sb_0__0__0_chanx_right_out_112_;
wire [0:0] sb_0__0__0_chanx_right_out_114_;
wire [0:0] sb_0__0__0_chanx_right_out_116_;
wire [0:0] sb_0__0__0_chanx_right_out_118_;
wire [0:0] sb_0__0__0_chanx_right_out_120_;
wire [0:0] sb_0__0__0_chanx_right_out_122_;
wire [0:0] sb_0__0__0_chanx_right_out_124_;
wire [0:0] sb_0__0__0_chanx_right_out_126_;
wire [0:0] sb_0__0__0_chanx_right_out_128_;
wire [0:0] sb_0__0__0_chanx_right_out_12_;
wire [0:0] sb_0__0__0_chanx_right_out_130_;
wire [0:0] sb_0__0__0_chanx_right_out_132_;
wire [0:0] sb_0__0__0_chanx_right_out_134_;
wire [0:0] sb_0__0__0_chanx_right_out_136_;
wire [0:0] sb_0__0__0_chanx_right_out_138_;
wire [0:0] sb_0__0__0_chanx_right_out_140_;
wire [0:0] sb_0__0__0_chanx_right_out_142_;
wire [0:0] sb_0__0__0_chanx_right_out_144_;
wire [0:0] sb_0__0__0_chanx_right_out_146_;
wire [0:0] sb_0__0__0_chanx_right_out_148_;
wire [0:0] sb_0__0__0_chanx_right_out_14_;
wire [0:0] sb_0__0__0_chanx_right_out_150_;
wire [0:0] sb_0__0__0_chanx_right_out_152_;
wire [0:0] sb_0__0__0_chanx_right_out_154_;
wire [0:0] sb_0__0__0_chanx_right_out_156_;
wire [0:0] sb_0__0__0_chanx_right_out_158_;
wire [0:0] sb_0__0__0_chanx_right_out_160_;
wire [0:0] sb_0__0__0_chanx_right_out_162_;
wire [0:0] sb_0__0__0_chanx_right_out_164_;
wire [0:0] sb_0__0__0_chanx_right_out_166_;
wire [0:0] sb_0__0__0_chanx_right_out_168_;
wire [0:0] sb_0__0__0_chanx_right_out_16_;
wire [0:0] sb_0__0__0_chanx_right_out_170_;
wire [0:0] sb_0__0__0_chanx_right_out_172_;
wire [0:0] sb_0__0__0_chanx_right_out_174_;
wire [0:0] sb_0__0__0_chanx_right_out_176_;
wire [0:0] sb_0__0__0_chanx_right_out_178_;
wire [0:0] sb_0__0__0_chanx_right_out_180_;
wire [0:0] sb_0__0__0_chanx_right_out_182_;
wire [0:0] sb_0__0__0_chanx_right_out_184_;
wire [0:0] sb_0__0__0_chanx_right_out_186_;
wire [0:0] sb_0__0__0_chanx_right_out_188_;
wire [0:0] sb_0__0__0_chanx_right_out_18_;
wire [0:0] sb_0__0__0_chanx_right_out_190_;
wire [0:0] sb_0__0__0_chanx_right_out_192_;
wire [0:0] sb_0__0__0_chanx_right_out_194_;
wire [0:0] sb_0__0__0_chanx_right_out_196_;
wire [0:0] sb_0__0__0_chanx_right_out_198_;
wire [0:0] sb_0__0__0_chanx_right_out_20_;
wire [0:0] sb_0__0__0_chanx_right_out_22_;
wire [0:0] sb_0__0__0_chanx_right_out_24_;
wire [0:0] sb_0__0__0_chanx_right_out_26_;
wire [0:0] sb_0__0__0_chanx_right_out_28_;
wire [0:0] sb_0__0__0_chanx_right_out_2_;
wire [0:0] sb_0__0__0_chanx_right_out_30_;
wire [0:0] sb_0__0__0_chanx_right_out_32_;
wire [0:0] sb_0__0__0_chanx_right_out_34_;
wire [0:0] sb_0__0__0_chanx_right_out_36_;
wire [0:0] sb_0__0__0_chanx_right_out_38_;
wire [0:0] sb_0__0__0_chanx_right_out_40_;
wire [0:0] sb_0__0__0_chanx_right_out_42_;
wire [0:0] sb_0__0__0_chanx_right_out_44_;
wire [0:0] sb_0__0__0_chanx_right_out_46_;
wire [0:0] sb_0__0__0_chanx_right_out_48_;
wire [0:0] sb_0__0__0_chanx_right_out_4_;
wire [0:0] sb_0__0__0_chanx_right_out_50_;
wire [0:0] sb_0__0__0_chanx_right_out_52_;
wire [0:0] sb_0__0__0_chanx_right_out_54_;
wire [0:0] sb_0__0__0_chanx_right_out_56_;
wire [0:0] sb_0__0__0_chanx_right_out_58_;
wire [0:0] sb_0__0__0_chanx_right_out_60_;
wire [0:0] sb_0__0__0_chanx_right_out_62_;
wire [0:0] sb_0__0__0_chanx_right_out_64_;
wire [0:0] sb_0__0__0_chanx_right_out_66_;
wire [0:0] sb_0__0__0_chanx_right_out_68_;
wire [0:0] sb_0__0__0_chanx_right_out_6_;
wire [0:0] sb_0__0__0_chanx_right_out_70_;
wire [0:0] sb_0__0__0_chanx_right_out_72_;
wire [0:0] sb_0__0__0_chanx_right_out_74_;
wire [0:0] sb_0__0__0_chanx_right_out_76_;
wire [0:0] sb_0__0__0_chanx_right_out_78_;
wire [0:0] sb_0__0__0_chanx_right_out_80_;
wire [0:0] sb_0__0__0_chanx_right_out_82_;
wire [0:0] sb_0__0__0_chanx_right_out_84_;
wire [0:0] sb_0__0__0_chanx_right_out_86_;
wire [0:0] sb_0__0__0_chanx_right_out_88_;
wire [0:0] sb_0__0__0_chanx_right_out_8_;
wire [0:0] sb_0__0__0_chanx_right_out_90_;
wire [0:0] sb_0__0__0_chanx_right_out_92_;
wire [0:0] sb_0__0__0_chanx_right_out_94_;
wire [0:0] sb_0__0__0_chanx_right_out_96_;
wire [0:0] sb_0__0__0_chanx_right_out_98_;
wire [0:0] sb_0__0__0_chany_top_out_0_;
wire [0:0] sb_0__0__0_chany_top_out_100_;
wire [0:0] sb_0__0__0_chany_top_out_102_;
wire [0:0] sb_0__0__0_chany_top_out_104_;
wire [0:0] sb_0__0__0_chany_top_out_106_;
wire [0:0] sb_0__0__0_chany_top_out_108_;
wire [0:0] sb_0__0__0_chany_top_out_10_;
wire [0:0] sb_0__0__0_chany_top_out_110_;
wire [0:0] sb_0__0__0_chany_top_out_112_;
wire [0:0] sb_0__0__0_chany_top_out_114_;
wire [0:0] sb_0__0__0_chany_top_out_116_;
wire [0:0] sb_0__0__0_chany_top_out_118_;
wire [0:0] sb_0__0__0_chany_top_out_120_;
wire [0:0] sb_0__0__0_chany_top_out_122_;
wire [0:0] sb_0__0__0_chany_top_out_124_;
wire [0:0] sb_0__0__0_chany_top_out_126_;
wire [0:0] sb_0__0__0_chany_top_out_128_;
wire [0:0] sb_0__0__0_chany_top_out_12_;
wire [0:0] sb_0__0__0_chany_top_out_130_;
wire [0:0] sb_0__0__0_chany_top_out_132_;
wire [0:0] sb_0__0__0_chany_top_out_134_;
wire [0:0] sb_0__0__0_chany_top_out_136_;
wire [0:0] sb_0__0__0_chany_top_out_138_;
wire [0:0] sb_0__0__0_chany_top_out_140_;
wire [0:0] sb_0__0__0_chany_top_out_142_;
wire [0:0] sb_0__0__0_chany_top_out_144_;
wire [0:0] sb_0__0__0_chany_top_out_146_;
wire [0:0] sb_0__0__0_chany_top_out_148_;
wire [0:0] sb_0__0__0_chany_top_out_14_;
wire [0:0] sb_0__0__0_chany_top_out_150_;
wire [0:0] sb_0__0__0_chany_top_out_152_;
wire [0:0] sb_0__0__0_chany_top_out_154_;
wire [0:0] sb_0__0__0_chany_top_out_156_;
wire [0:0] sb_0__0__0_chany_top_out_158_;
wire [0:0] sb_0__0__0_chany_top_out_160_;
wire [0:0] sb_0__0__0_chany_top_out_162_;
wire [0:0] sb_0__0__0_chany_top_out_164_;
wire [0:0] sb_0__0__0_chany_top_out_166_;
wire [0:0] sb_0__0__0_chany_top_out_168_;
wire [0:0] sb_0__0__0_chany_top_out_16_;
wire [0:0] sb_0__0__0_chany_top_out_170_;
wire [0:0] sb_0__0__0_chany_top_out_172_;
wire [0:0] sb_0__0__0_chany_top_out_174_;
wire [0:0] sb_0__0__0_chany_top_out_176_;
wire [0:0] sb_0__0__0_chany_top_out_178_;
wire [0:0] sb_0__0__0_chany_top_out_180_;
wire [0:0] sb_0__0__0_chany_top_out_182_;
wire [0:0] sb_0__0__0_chany_top_out_184_;
wire [0:0] sb_0__0__0_chany_top_out_186_;
wire [0:0] sb_0__0__0_chany_top_out_188_;
wire [0:0] sb_0__0__0_chany_top_out_18_;
wire [0:0] sb_0__0__0_chany_top_out_190_;
wire [0:0] sb_0__0__0_chany_top_out_192_;
wire [0:0] sb_0__0__0_chany_top_out_194_;
wire [0:0] sb_0__0__0_chany_top_out_196_;
wire [0:0] sb_0__0__0_chany_top_out_198_;
wire [0:0] sb_0__0__0_chany_top_out_20_;
wire [0:0] sb_0__0__0_chany_top_out_22_;
wire [0:0] sb_0__0__0_chany_top_out_24_;
wire [0:0] sb_0__0__0_chany_top_out_26_;
wire [0:0] sb_0__0__0_chany_top_out_28_;
wire [0:0] sb_0__0__0_chany_top_out_2_;
wire [0:0] sb_0__0__0_chany_top_out_30_;
wire [0:0] sb_0__0__0_chany_top_out_32_;
wire [0:0] sb_0__0__0_chany_top_out_34_;
wire [0:0] sb_0__0__0_chany_top_out_36_;
wire [0:0] sb_0__0__0_chany_top_out_38_;
wire [0:0] sb_0__0__0_chany_top_out_40_;
wire [0:0] sb_0__0__0_chany_top_out_42_;
wire [0:0] sb_0__0__0_chany_top_out_44_;
wire [0:0] sb_0__0__0_chany_top_out_46_;
wire [0:0] sb_0__0__0_chany_top_out_48_;
wire [0:0] sb_0__0__0_chany_top_out_4_;
wire [0:0] sb_0__0__0_chany_top_out_50_;
wire [0:0] sb_0__0__0_chany_top_out_52_;
wire [0:0] sb_0__0__0_chany_top_out_54_;
wire [0:0] sb_0__0__0_chany_top_out_56_;
wire [0:0] sb_0__0__0_chany_top_out_58_;
wire [0:0] sb_0__0__0_chany_top_out_60_;
wire [0:0] sb_0__0__0_chany_top_out_62_;
wire [0:0] sb_0__0__0_chany_top_out_64_;
wire [0:0] sb_0__0__0_chany_top_out_66_;
wire [0:0] sb_0__0__0_chany_top_out_68_;
wire [0:0] sb_0__0__0_chany_top_out_6_;
wire [0:0] sb_0__0__0_chany_top_out_70_;
wire [0:0] sb_0__0__0_chany_top_out_72_;
wire [0:0] sb_0__0__0_chany_top_out_74_;
wire [0:0] sb_0__0__0_chany_top_out_76_;
wire [0:0] sb_0__0__0_chany_top_out_78_;
wire [0:0] sb_0__0__0_chany_top_out_80_;
wire [0:0] sb_0__0__0_chany_top_out_82_;
wire [0:0] sb_0__0__0_chany_top_out_84_;
wire [0:0] sb_0__0__0_chany_top_out_86_;
wire [0:0] sb_0__0__0_chany_top_out_88_;
wire [0:0] sb_0__0__0_chany_top_out_8_;
wire [0:0] sb_0__0__0_chany_top_out_90_;
wire [0:0] sb_0__0__0_chany_top_out_92_;
wire [0:0] sb_0__0__0_chany_top_out_94_;
wire [0:0] sb_0__0__0_chany_top_out_96_;
wire [0:0] sb_0__0__0_chany_top_out_98_;
wire [0:0] sb_0__1__0_ccff_tail;
wire [0:0] sb_0__1__0_chanx_right_out_0_;
wire [0:0] sb_0__1__0_chanx_right_out_100_;
wire [0:0] sb_0__1__0_chanx_right_out_102_;
wire [0:0] sb_0__1__0_chanx_right_out_104_;
wire [0:0] sb_0__1__0_chanx_right_out_106_;
wire [0:0] sb_0__1__0_chanx_right_out_108_;
wire [0:0] sb_0__1__0_chanx_right_out_10_;
wire [0:0] sb_0__1__0_chanx_right_out_110_;
wire [0:0] sb_0__1__0_chanx_right_out_112_;
wire [0:0] sb_0__1__0_chanx_right_out_114_;
wire [0:0] sb_0__1__0_chanx_right_out_116_;
wire [0:0] sb_0__1__0_chanx_right_out_118_;
wire [0:0] sb_0__1__0_chanx_right_out_120_;
wire [0:0] sb_0__1__0_chanx_right_out_122_;
wire [0:0] sb_0__1__0_chanx_right_out_124_;
wire [0:0] sb_0__1__0_chanx_right_out_126_;
wire [0:0] sb_0__1__0_chanx_right_out_128_;
wire [0:0] sb_0__1__0_chanx_right_out_12_;
wire [0:0] sb_0__1__0_chanx_right_out_130_;
wire [0:0] sb_0__1__0_chanx_right_out_132_;
wire [0:0] sb_0__1__0_chanx_right_out_134_;
wire [0:0] sb_0__1__0_chanx_right_out_136_;
wire [0:0] sb_0__1__0_chanx_right_out_138_;
wire [0:0] sb_0__1__0_chanx_right_out_140_;
wire [0:0] sb_0__1__0_chanx_right_out_142_;
wire [0:0] sb_0__1__0_chanx_right_out_144_;
wire [0:0] sb_0__1__0_chanx_right_out_146_;
wire [0:0] sb_0__1__0_chanx_right_out_148_;
wire [0:0] sb_0__1__0_chanx_right_out_14_;
wire [0:0] sb_0__1__0_chanx_right_out_150_;
wire [0:0] sb_0__1__0_chanx_right_out_152_;
wire [0:0] sb_0__1__0_chanx_right_out_154_;
wire [0:0] sb_0__1__0_chanx_right_out_156_;
wire [0:0] sb_0__1__0_chanx_right_out_158_;
wire [0:0] sb_0__1__0_chanx_right_out_160_;
wire [0:0] sb_0__1__0_chanx_right_out_162_;
wire [0:0] sb_0__1__0_chanx_right_out_164_;
wire [0:0] sb_0__1__0_chanx_right_out_166_;
wire [0:0] sb_0__1__0_chanx_right_out_168_;
wire [0:0] sb_0__1__0_chanx_right_out_16_;
wire [0:0] sb_0__1__0_chanx_right_out_170_;
wire [0:0] sb_0__1__0_chanx_right_out_172_;
wire [0:0] sb_0__1__0_chanx_right_out_174_;
wire [0:0] sb_0__1__0_chanx_right_out_176_;
wire [0:0] sb_0__1__0_chanx_right_out_178_;
wire [0:0] sb_0__1__0_chanx_right_out_180_;
wire [0:0] sb_0__1__0_chanx_right_out_182_;
wire [0:0] sb_0__1__0_chanx_right_out_184_;
wire [0:0] sb_0__1__0_chanx_right_out_186_;
wire [0:0] sb_0__1__0_chanx_right_out_188_;
wire [0:0] sb_0__1__0_chanx_right_out_18_;
wire [0:0] sb_0__1__0_chanx_right_out_190_;
wire [0:0] sb_0__1__0_chanx_right_out_192_;
wire [0:0] sb_0__1__0_chanx_right_out_194_;
wire [0:0] sb_0__1__0_chanx_right_out_196_;
wire [0:0] sb_0__1__0_chanx_right_out_198_;
wire [0:0] sb_0__1__0_chanx_right_out_20_;
wire [0:0] sb_0__1__0_chanx_right_out_22_;
wire [0:0] sb_0__1__0_chanx_right_out_24_;
wire [0:0] sb_0__1__0_chanx_right_out_26_;
wire [0:0] sb_0__1__0_chanx_right_out_28_;
wire [0:0] sb_0__1__0_chanx_right_out_2_;
wire [0:0] sb_0__1__0_chanx_right_out_30_;
wire [0:0] sb_0__1__0_chanx_right_out_32_;
wire [0:0] sb_0__1__0_chanx_right_out_34_;
wire [0:0] sb_0__1__0_chanx_right_out_36_;
wire [0:0] sb_0__1__0_chanx_right_out_38_;
wire [0:0] sb_0__1__0_chanx_right_out_40_;
wire [0:0] sb_0__1__0_chanx_right_out_42_;
wire [0:0] sb_0__1__0_chanx_right_out_44_;
wire [0:0] sb_0__1__0_chanx_right_out_46_;
wire [0:0] sb_0__1__0_chanx_right_out_48_;
wire [0:0] sb_0__1__0_chanx_right_out_4_;
wire [0:0] sb_0__1__0_chanx_right_out_50_;
wire [0:0] sb_0__1__0_chanx_right_out_52_;
wire [0:0] sb_0__1__0_chanx_right_out_54_;
wire [0:0] sb_0__1__0_chanx_right_out_56_;
wire [0:0] sb_0__1__0_chanx_right_out_58_;
wire [0:0] sb_0__1__0_chanx_right_out_60_;
wire [0:0] sb_0__1__0_chanx_right_out_62_;
wire [0:0] sb_0__1__0_chanx_right_out_64_;
wire [0:0] sb_0__1__0_chanx_right_out_66_;
wire [0:0] sb_0__1__0_chanx_right_out_68_;
wire [0:0] sb_0__1__0_chanx_right_out_6_;
wire [0:0] sb_0__1__0_chanx_right_out_70_;
wire [0:0] sb_0__1__0_chanx_right_out_72_;
wire [0:0] sb_0__1__0_chanx_right_out_74_;
wire [0:0] sb_0__1__0_chanx_right_out_76_;
wire [0:0] sb_0__1__0_chanx_right_out_78_;
wire [0:0] sb_0__1__0_chanx_right_out_80_;
wire [0:0] sb_0__1__0_chanx_right_out_82_;
wire [0:0] sb_0__1__0_chanx_right_out_84_;
wire [0:0] sb_0__1__0_chanx_right_out_86_;
wire [0:0] sb_0__1__0_chanx_right_out_88_;
wire [0:0] sb_0__1__0_chanx_right_out_8_;
wire [0:0] sb_0__1__0_chanx_right_out_90_;
wire [0:0] sb_0__1__0_chanx_right_out_92_;
wire [0:0] sb_0__1__0_chanx_right_out_94_;
wire [0:0] sb_0__1__0_chanx_right_out_96_;
wire [0:0] sb_0__1__0_chanx_right_out_98_;
wire [0:0] sb_0__1__0_chany_bottom_out_101_;
wire [0:0] sb_0__1__0_chany_bottom_out_103_;
wire [0:0] sb_0__1__0_chany_bottom_out_105_;
wire [0:0] sb_0__1__0_chany_bottom_out_107_;
wire [0:0] sb_0__1__0_chany_bottom_out_109_;
wire [0:0] sb_0__1__0_chany_bottom_out_111_;
wire [0:0] sb_0__1__0_chany_bottom_out_113_;
wire [0:0] sb_0__1__0_chany_bottom_out_115_;
wire [0:0] sb_0__1__0_chany_bottom_out_117_;
wire [0:0] sb_0__1__0_chany_bottom_out_119_;
wire [0:0] sb_0__1__0_chany_bottom_out_11_;
wire [0:0] sb_0__1__0_chany_bottom_out_121_;
wire [0:0] sb_0__1__0_chany_bottom_out_123_;
wire [0:0] sb_0__1__0_chany_bottom_out_125_;
wire [0:0] sb_0__1__0_chany_bottom_out_127_;
wire [0:0] sb_0__1__0_chany_bottom_out_129_;
wire [0:0] sb_0__1__0_chany_bottom_out_131_;
wire [0:0] sb_0__1__0_chany_bottom_out_133_;
wire [0:0] sb_0__1__0_chany_bottom_out_135_;
wire [0:0] sb_0__1__0_chany_bottom_out_137_;
wire [0:0] sb_0__1__0_chany_bottom_out_139_;
wire [0:0] sb_0__1__0_chany_bottom_out_13_;
wire [0:0] sb_0__1__0_chany_bottom_out_141_;
wire [0:0] sb_0__1__0_chany_bottom_out_143_;
wire [0:0] sb_0__1__0_chany_bottom_out_145_;
wire [0:0] sb_0__1__0_chany_bottom_out_147_;
wire [0:0] sb_0__1__0_chany_bottom_out_149_;
wire [0:0] sb_0__1__0_chany_bottom_out_151_;
wire [0:0] sb_0__1__0_chany_bottom_out_153_;
wire [0:0] sb_0__1__0_chany_bottom_out_155_;
wire [0:0] sb_0__1__0_chany_bottom_out_157_;
wire [0:0] sb_0__1__0_chany_bottom_out_159_;
wire [0:0] sb_0__1__0_chany_bottom_out_15_;
wire [0:0] sb_0__1__0_chany_bottom_out_161_;
wire [0:0] sb_0__1__0_chany_bottom_out_163_;
wire [0:0] sb_0__1__0_chany_bottom_out_165_;
wire [0:0] sb_0__1__0_chany_bottom_out_167_;
wire [0:0] sb_0__1__0_chany_bottom_out_169_;
wire [0:0] sb_0__1__0_chany_bottom_out_171_;
wire [0:0] sb_0__1__0_chany_bottom_out_173_;
wire [0:0] sb_0__1__0_chany_bottom_out_175_;
wire [0:0] sb_0__1__0_chany_bottom_out_177_;
wire [0:0] sb_0__1__0_chany_bottom_out_179_;
wire [0:0] sb_0__1__0_chany_bottom_out_17_;
wire [0:0] sb_0__1__0_chany_bottom_out_181_;
wire [0:0] sb_0__1__0_chany_bottom_out_183_;
wire [0:0] sb_0__1__0_chany_bottom_out_185_;
wire [0:0] sb_0__1__0_chany_bottom_out_187_;
wire [0:0] sb_0__1__0_chany_bottom_out_189_;
wire [0:0] sb_0__1__0_chany_bottom_out_191_;
wire [0:0] sb_0__1__0_chany_bottom_out_193_;
wire [0:0] sb_0__1__0_chany_bottom_out_195_;
wire [0:0] sb_0__1__0_chany_bottom_out_197_;
wire [0:0] sb_0__1__0_chany_bottom_out_199_;
wire [0:0] sb_0__1__0_chany_bottom_out_19_;
wire [0:0] sb_0__1__0_chany_bottom_out_1_;
wire [0:0] sb_0__1__0_chany_bottom_out_21_;
wire [0:0] sb_0__1__0_chany_bottom_out_23_;
wire [0:0] sb_0__1__0_chany_bottom_out_25_;
wire [0:0] sb_0__1__0_chany_bottom_out_27_;
wire [0:0] sb_0__1__0_chany_bottom_out_29_;
wire [0:0] sb_0__1__0_chany_bottom_out_31_;
wire [0:0] sb_0__1__0_chany_bottom_out_33_;
wire [0:0] sb_0__1__0_chany_bottom_out_35_;
wire [0:0] sb_0__1__0_chany_bottom_out_37_;
wire [0:0] sb_0__1__0_chany_bottom_out_39_;
wire [0:0] sb_0__1__0_chany_bottom_out_3_;
wire [0:0] sb_0__1__0_chany_bottom_out_41_;
wire [0:0] sb_0__1__0_chany_bottom_out_43_;
wire [0:0] sb_0__1__0_chany_bottom_out_45_;
wire [0:0] sb_0__1__0_chany_bottom_out_47_;
wire [0:0] sb_0__1__0_chany_bottom_out_49_;
wire [0:0] sb_0__1__0_chany_bottom_out_51_;
wire [0:0] sb_0__1__0_chany_bottom_out_53_;
wire [0:0] sb_0__1__0_chany_bottom_out_55_;
wire [0:0] sb_0__1__0_chany_bottom_out_57_;
wire [0:0] sb_0__1__0_chany_bottom_out_59_;
wire [0:0] sb_0__1__0_chany_bottom_out_5_;
wire [0:0] sb_0__1__0_chany_bottom_out_61_;
wire [0:0] sb_0__1__0_chany_bottom_out_63_;
wire [0:0] sb_0__1__0_chany_bottom_out_65_;
wire [0:0] sb_0__1__0_chany_bottom_out_67_;
wire [0:0] sb_0__1__0_chany_bottom_out_69_;
wire [0:0] sb_0__1__0_chany_bottom_out_71_;
wire [0:0] sb_0__1__0_chany_bottom_out_73_;
wire [0:0] sb_0__1__0_chany_bottom_out_75_;
wire [0:0] sb_0__1__0_chany_bottom_out_77_;
wire [0:0] sb_0__1__0_chany_bottom_out_79_;
wire [0:0] sb_0__1__0_chany_bottom_out_7_;
wire [0:0] sb_0__1__0_chany_bottom_out_81_;
wire [0:0] sb_0__1__0_chany_bottom_out_83_;
wire [0:0] sb_0__1__0_chany_bottom_out_85_;
wire [0:0] sb_0__1__0_chany_bottom_out_87_;
wire [0:0] sb_0__1__0_chany_bottom_out_89_;
wire [0:0] sb_0__1__0_chany_bottom_out_91_;
wire [0:0] sb_0__1__0_chany_bottom_out_93_;
wire [0:0] sb_0__1__0_chany_bottom_out_95_;
wire [0:0] sb_0__1__0_chany_bottom_out_97_;
wire [0:0] sb_0__1__0_chany_bottom_out_99_;
wire [0:0] sb_0__1__0_chany_bottom_out_9_;
wire [0:0] sb_0__1__0_chany_top_out_0_;
wire [0:0] sb_0__1__0_chany_top_out_100_;
wire [0:0] sb_0__1__0_chany_top_out_102_;
wire [0:0] sb_0__1__0_chany_top_out_104_;
wire [0:0] sb_0__1__0_chany_top_out_106_;
wire [0:0] sb_0__1__0_chany_top_out_108_;
wire [0:0] sb_0__1__0_chany_top_out_10_;
wire [0:0] sb_0__1__0_chany_top_out_110_;
wire [0:0] sb_0__1__0_chany_top_out_112_;
wire [0:0] sb_0__1__0_chany_top_out_114_;
wire [0:0] sb_0__1__0_chany_top_out_116_;
wire [0:0] sb_0__1__0_chany_top_out_118_;
wire [0:0] sb_0__1__0_chany_top_out_120_;
wire [0:0] sb_0__1__0_chany_top_out_122_;
wire [0:0] sb_0__1__0_chany_top_out_124_;
wire [0:0] sb_0__1__0_chany_top_out_126_;
wire [0:0] sb_0__1__0_chany_top_out_128_;
wire [0:0] sb_0__1__0_chany_top_out_12_;
wire [0:0] sb_0__1__0_chany_top_out_130_;
wire [0:0] sb_0__1__0_chany_top_out_132_;
wire [0:0] sb_0__1__0_chany_top_out_134_;
wire [0:0] sb_0__1__0_chany_top_out_136_;
wire [0:0] sb_0__1__0_chany_top_out_138_;
wire [0:0] sb_0__1__0_chany_top_out_140_;
wire [0:0] sb_0__1__0_chany_top_out_142_;
wire [0:0] sb_0__1__0_chany_top_out_144_;
wire [0:0] sb_0__1__0_chany_top_out_146_;
wire [0:0] sb_0__1__0_chany_top_out_148_;
wire [0:0] sb_0__1__0_chany_top_out_14_;
wire [0:0] sb_0__1__0_chany_top_out_150_;
wire [0:0] sb_0__1__0_chany_top_out_152_;
wire [0:0] sb_0__1__0_chany_top_out_154_;
wire [0:0] sb_0__1__0_chany_top_out_156_;
wire [0:0] sb_0__1__0_chany_top_out_158_;
wire [0:0] sb_0__1__0_chany_top_out_160_;
wire [0:0] sb_0__1__0_chany_top_out_162_;
wire [0:0] sb_0__1__0_chany_top_out_164_;
wire [0:0] sb_0__1__0_chany_top_out_166_;
wire [0:0] sb_0__1__0_chany_top_out_168_;
wire [0:0] sb_0__1__0_chany_top_out_16_;
wire [0:0] sb_0__1__0_chany_top_out_170_;
wire [0:0] sb_0__1__0_chany_top_out_172_;
wire [0:0] sb_0__1__0_chany_top_out_174_;
wire [0:0] sb_0__1__0_chany_top_out_176_;
wire [0:0] sb_0__1__0_chany_top_out_178_;
wire [0:0] sb_0__1__0_chany_top_out_180_;
wire [0:0] sb_0__1__0_chany_top_out_182_;
wire [0:0] sb_0__1__0_chany_top_out_184_;
wire [0:0] sb_0__1__0_chany_top_out_186_;
wire [0:0] sb_0__1__0_chany_top_out_188_;
wire [0:0] sb_0__1__0_chany_top_out_18_;
wire [0:0] sb_0__1__0_chany_top_out_190_;
wire [0:0] sb_0__1__0_chany_top_out_192_;
wire [0:0] sb_0__1__0_chany_top_out_194_;
wire [0:0] sb_0__1__0_chany_top_out_196_;
wire [0:0] sb_0__1__0_chany_top_out_198_;
wire [0:0] sb_0__1__0_chany_top_out_20_;
wire [0:0] sb_0__1__0_chany_top_out_22_;
wire [0:0] sb_0__1__0_chany_top_out_24_;
wire [0:0] sb_0__1__0_chany_top_out_26_;
wire [0:0] sb_0__1__0_chany_top_out_28_;
wire [0:0] sb_0__1__0_chany_top_out_2_;
wire [0:0] sb_0__1__0_chany_top_out_30_;
wire [0:0] sb_0__1__0_chany_top_out_32_;
wire [0:0] sb_0__1__0_chany_top_out_34_;
wire [0:0] sb_0__1__0_chany_top_out_36_;
wire [0:0] sb_0__1__0_chany_top_out_38_;
wire [0:0] sb_0__1__0_chany_top_out_40_;
wire [0:0] sb_0__1__0_chany_top_out_42_;
wire [0:0] sb_0__1__0_chany_top_out_44_;
wire [0:0] sb_0__1__0_chany_top_out_46_;
wire [0:0] sb_0__1__0_chany_top_out_48_;
wire [0:0] sb_0__1__0_chany_top_out_4_;
wire [0:0] sb_0__1__0_chany_top_out_50_;
wire [0:0] sb_0__1__0_chany_top_out_52_;
wire [0:0] sb_0__1__0_chany_top_out_54_;
wire [0:0] sb_0__1__0_chany_top_out_56_;
wire [0:0] sb_0__1__0_chany_top_out_58_;
wire [0:0] sb_0__1__0_chany_top_out_60_;
wire [0:0] sb_0__1__0_chany_top_out_62_;
wire [0:0] sb_0__1__0_chany_top_out_64_;
wire [0:0] sb_0__1__0_chany_top_out_66_;
wire [0:0] sb_0__1__0_chany_top_out_68_;
wire [0:0] sb_0__1__0_chany_top_out_6_;
wire [0:0] sb_0__1__0_chany_top_out_70_;
wire [0:0] sb_0__1__0_chany_top_out_72_;
wire [0:0] sb_0__1__0_chany_top_out_74_;
wire [0:0] sb_0__1__0_chany_top_out_76_;
wire [0:0] sb_0__1__0_chany_top_out_78_;
wire [0:0] sb_0__1__0_chany_top_out_80_;
wire [0:0] sb_0__1__0_chany_top_out_82_;
wire [0:0] sb_0__1__0_chany_top_out_84_;
wire [0:0] sb_0__1__0_chany_top_out_86_;
wire [0:0] sb_0__1__0_chany_top_out_88_;
wire [0:0] sb_0__1__0_chany_top_out_8_;
wire [0:0] sb_0__1__0_chany_top_out_90_;
wire [0:0] sb_0__1__0_chany_top_out_92_;
wire [0:0] sb_0__1__0_chany_top_out_94_;
wire [0:0] sb_0__1__0_chany_top_out_96_;
wire [0:0] sb_0__1__0_chany_top_out_98_;
wire [0:0] sb_0__2__0_ccff_tail;
wire [0:0] sb_0__2__0_chanx_right_out_0_;
wire [0:0] sb_0__2__0_chanx_right_out_100_;
wire [0:0] sb_0__2__0_chanx_right_out_102_;
wire [0:0] sb_0__2__0_chanx_right_out_104_;
wire [0:0] sb_0__2__0_chanx_right_out_106_;
wire [0:0] sb_0__2__0_chanx_right_out_108_;
wire [0:0] sb_0__2__0_chanx_right_out_10_;
wire [0:0] sb_0__2__0_chanx_right_out_110_;
wire [0:0] sb_0__2__0_chanx_right_out_112_;
wire [0:0] sb_0__2__0_chanx_right_out_114_;
wire [0:0] sb_0__2__0_chanx_right_out_116_;
wire [0:0] sb_0__2__0_chanx_right_out_118_;
wire [0:0] sb_0__2__0_chanx_right_out_120_;
wire [0:0] sb_0__2__0_chanx_right_out_122_;
wire [0:0] sb_0__2__0_chanx_right_out_124_;
wire [0:0] sb_0__2__0_chanx_right_out_126_;
wire [0:0] sb_0__2__0_chanx_right_out_128_;
wire [0:0] sb_0__2__0_chanx_right_out_12_;
wire [0:0] sb_0__2__0_chanx_right_out_130_;
wire [0:0] sb_0__2__0_chanx_right_out_132_;
wire [0:0] sb_0__2__0_chanx_right_out_134_;
wire [0:0] sb_0__2__0_chanx_right_out_136_;
wire [0:0] sb_0__2__0_chanx_right_out_138_;
wire [0:0] sb_0__2__0_chanx_right_out_140_;
wire [0:0] sb_0__2__0_chanx_right_out_142_;
wire [0:0] sb_0__2__0_chanx_right_out_144_;
wire [0:0] sb_0__2__0_chanx_right_out_146_;
wire [0:0] sb_0__2__0_chanx_right_out_148_;
wire [0:0] sb_0__2__0_chanx_right_out_14_;
wire [0:0] sb_0__2__0_chanx_right_out_150_;
wire [0:0] sb_0__2__0_chanx_right_out_152_;
wire [0:0] sb_0__2__0_chanx_right_out_154_;
wire [0:0] sb_0__2__0_chanx_right_out_156_;
wire [0:0] sb_0__2__0_chanx_right_out_158_;
wire [0:0] sb_0__2__0_chanx_right_out_160_;
wire [0:0] sb_0__2__0_chanx_right_out_162_;
wire [0:0] sb_0__2__0_chanx_right_out_164_;
wire [0:0] sb_0__2__0_chanx_right_out_166_;
wire [0:0] sb_0__2__0_chanx_right_out_168_;
wire [0:0] sb_0__2__0_chanx_right_out_16_;
wire [0:0] sb_0__2__0_chanx_right_out_170_;
wire [0:0] sb_0__2__0_chanx_right_out_172_;
wire [0:0] sb_0__2__0_chanx_right_out_174_;
wire [0:0] sb_0__2__0_chanx_right_out_176_;
wire [0:0] sb_0__2__0_chanx_right_out_178_;
wire [0:0] sb_0__2__0_chanx_right_out_180_;
wire [0:0] sb_0__2__0_chanx_right_out_182_;
wire [0:0] sb_0__2__0_chanx_right_out_184_;
wire [0:0] sb_0__2__0_chanx_right_out_186_;
wire [0:0] sb_0__2__0_chanx_right_out_188_;
wire [0:0] sb_0__2__0_chanx_right_out_18_;
wire [0:0] sb_0__2__0_chanx_right_out_190_;
wire [0:0] sb_0__2__0_chanx_right_out_192_;
wire [0:0] sb_0__2__0_chanx_right_out_194_;
wire [0:0] sb_0__2__0_chanx_right_out_196_;
wire [0:0] sb_0__2__0_chanx_right_out_198_;
wire [0:0] sb_0__2__0_chanx_right_out_20_;
wire [0:0] sb_0__2__0_chanx_right_out_22_;
wire [0:0] sb_0__2__0_chanx_right_out_24_;
wire [0:0] sb_0__2__0_chanx_right_out_26_;
wire [0:0] sb_0__2__0_chanx_right_out_28_;
wire [0:0] sb_0__2__0_chanx_right_out_2_;
wire [0:0] sb_0__2__0_chanx_right_out_30_;
wire [0:0] sb_0__2__0_chanx_right_out_32_;
wire [0:0] sb_0__2__0_chanx_right_out_34_;
wire [0:0] sb_0__2__0_chanx_right_out_36_;
wire [0:0] sb_0__2__0_chanx_right_out_38_;
wire [0:0] sb_0__2__0_chanx_right_out_40_;
wire [0:0] sb_0__2__0_chanx_right_out_42_;
wire [0:0] sb_0__2__0_chanx_right_out_44_;
wire [0:0] sb_0__2__0_chanx_right_out_46_;
wire [0:0] sb_0__2__0_chanx_right_out_48_;
wire [0:0] sb_0__2__0_chanx_right_out_4_;
wire [0:0] sb_0__2__0_chanx_right_out_50_;
wire [0:0] sb_0__2__0_chanx_right_out_52_;
wire [0:0] sb_0__2__0_chanx_right_out_54_;
wire [0:0] sb_0__2__0_chanx_right_out_56_;
wire [0:0] sb_0__2__0_chanx_right_out_58_;
wire [0:0] sb_0__2__0_chanx_right_out_60_;
wire [0:0] sb_0__2__0_chanx_right_out_62_;
wire [0:0] sb_0__2__0_chanx_right_out_64_;
wire [0:0] sb_0__2__0_chanx_right_out_66_;
wire [0:0] sb_0__2__0_chanx_right_out_68_;
wire [0:0] sb_0__2__0_chanx_right_out_6_;
wire [0:0] sb_0__2__0_chanx_right_out_70_;
wire [0:0] sb_0__2__0_chanx_right_out_72_;
wire [0:0] sb_0__2__0_chanx_right_out_74_;
wire [0:0] sb_0__2__0_chanx_right_out_76_;
wire [0:0] sb_0__2__0_chanx_right_out_78_;
wire [0:0] sb_0__2__0_chanx_right_out_80_;
wire [0:0] sb_0__2__0_chanx_right_out_82_;
wire [0:0] sb_0__2__0_chanx_right_out_84_;
wire [0:0] sb_0__2__0_chanx_right_out_86_;
wire [0:0] sb_0__2__0_chanx_right_out_88_;
wire [0:0] sb_0__2__0_chanx_right_out_8_;
wire [0:0] sb_0__2__0_chanx_right_out_90_;
wire [0:0] sb_0__2__0_chanx_right_out_92_;
wire [0:0] sb_0__2__0_chanx_right_out_94_;
wire [0:0] sb_0__2__0_chanx_right_out_96_;
wire [0:0] sb_0__2__0_chanx_right_out_98_;
wire [0:0] sb_0__2__0_chany_bottom_out_101_;
wire [0:0] sb_0__2__0_chany_bottom_out_103_;
wire [0:0] sb_0__2__0_chany_bottom_out_105_;
wire [0:0] sb_0__2__0_chany_bottom_out_107_;
wire [0:0] sb_0__2__0_chany_bottom_out_109_;
wire [0:0] sb_0__2__0_chany_bottom_out_111_;
wire [0:0] sb_0__2__0_chany_bottom_out_113_;
wire [0:0] sb_0__2__0_chany_bottom_out_115_;
wire [0:0] sb_0__2__0_chany_bottom_out_117_;
wire [0:0] sb_0__2__0_chany_bottom_out_119_;
wire [0:0] sb_0__2__0_chany_bottom_out_11_;
wire [0:0] sb_0__2__0_chany_bottom_out_121_;
wire [0:0] sb_0__2__0_chany_bottom_out_123_;
wire [0:0] sb_0__2__0_chany_bottom_out_125_;
wire [0:0] sb_0__2__0_chany_bottom_out_127_;
wire [0:0] sb_0__2__0_chany_bottom_out_129_;
wire [0:0] sb_0__2__0_chany_bottom_out_131_;
wire [0:0] sb_0__2__0_chany_bottom_out_133_;
wire [0:0] sb_0__2__0_chany_bottom_out_135_;
wire [0:0] sb_0__2__0_chany_bottom_out_137_;
wire [0:0] sb_0__2__0_chany_bottom_out_139_;
wire [0:0] sb_0__2__0_chany_bottom_out_13_;
wire [0:0] sb_0__2__0_chany_bottom_out_141_;
wire [0:0] sb_0__2__0_chany_bottom_out_143_;
wire [0:0] sb_0__2__0_chany_bottom_out_145_;
wire [0:0] sb_0__2__0_chany_bottom_out_147_;
wire [0:0] sb_0__2__0_chany_bottom_out_149_;
wire [0:0] sb_0__2__0_chany_bottom_out_151_;
wire [0:0] sb_0__2__0_chany_bottom_out_153_;
wire [0:0] sb_0__2__0_chany_bottom_out_155_;
wire [0:0] sb_0__2__0_chany_bottom_out_157_;
wire [0:0] sb_0__2__0_chany_bottom_out_159_;
wire [0:0] sb_0__2__0_chany_bottom_out_15_;
wire [0:0] sb_0__2__0_chany_bottom_out_161_;
wire [0:0] sb_0__2__0_chany_bottom_out_163_;
wire [0:0] sb_0__2__0_chany_bottom_out_165_;
wire [0:0] sb_0__2__0_chany_bottom_out_167_;
wire [0:0] sb_0__2__0_chany_bottom_out_169_;
wire [0:0] sb_0__2__0_chany_bottom_out_171_;
wire [0:0] sb_0__2__0_chany_bottom_out_173_;
wire [0:0] sb_0__2__0_chany_bottom_out_175_;
wire [0:0] sb_0__2__0_chany_bottom_out_177_;
wire [0:0] sb_0__2__0_chany_bottom_out_179_;
wire [0:0] sb_0__2__0_chany_bottom_out_17_;
wire [0:0] sb_0__2__0_chany_bottom_out_181_;
wire [0:0] sb_0__2__0_chany_bottom_out_183_;
wire [0:0] sb_0__2__0_chany_bottom_out_185_;
wire [0:0] sb_0__2__0_chany_bottom_out_187_;
wire [0:0] sb_0__2__0_chany_bottom_out_189_;
wire [0:0] sb_0__2__0_chany_bottom_out_191_;
wire [0:0] sb_0__2__0_chany_bottom_out_193_;
wire [0:0] sb_0__2__0_chany_bottom_out_195_;
wire [0:0] sb_0__2__0_chany_bottom_out_197_;
wire [0:0] sb_0__2__0_chany_bottom_out_199_;
wire [0:0] sb_0__2__0_chany_bottom_out_19_;
wire [0:0] sb_0__2__0_chany_bottom_out_1_;
wire [0:0] sb_0__2__0_chany_bottom_out_21_;
wire [0:0] sb_0__2__0_chany_bottom_out_23_;
wire [0:0] sb_0__2__0_chany_bottom_out_25_;
wire [0:0] sb_0__2__0_chany_bottom_out_27_;
wire [0:0] sb_0__2__0_chany_bottom_out_29_;
wire [0:0] sb_0__2__0_chany_bottom_out_31_;
wire [0:0] sb_0__2__0_chany_bottom_out_33_;
wire [0:0] sb_0__2__0_chany_bottom_out_35_;
wire [0:0] sb_0__2__0_chany_bottom_out_37_;
wire [0:0] sb_0__2__0_chany_bottom_out_39_;
wire [0:0] sb_0__2__0_chany_bottom_out_3_;
wire [0:0] sb_0__2__0_chany_bottom_out_41_;
wire [0:0] sb_0__2__0_chany_bottom_out_43_;
wire [0:0] sb_0__2__0_chany_bottom_out_45_;
wire [0:0] sb_0__2__0_chany_bottom_out_47_;
wire [0:0] sb_0__2__0_chany_bottom_out_49_;
wire [0:0] sb_0__2__0_chany_bottom_out_51_;
wire [0:0] sb_0__2__0_chany_bottom_out_53_;
wire [0:0] sb_0__2__0_chany_bottom_out_55_;
wire [0:0] sb_0__2__0_chany_bottom_out_57_;
wire [0:0] sb_0__2__0_chany_bottom_out_59_;
wire [0:0] sb_0__2__0_chany_bottom_out_5_;
wire [0:0] sb_0__2__0_chany_bottom_out_61_;
wire [0:0] sb_0__2__0_chany_bottom_out_63_;
wire [0:0] sb_0__2__0_chany_bottom_out_65_;
wire [0:0] sb_0__2__0_chany_bottom_out_67_;
wire [0:0] sb_0__2__0_chany_bottom_out_69_;
wire [0:0] sb_0__2__0_chany_bottom_out_71_;
wire [0:0] sb_0__2__0_chany_bottom_out_73_;
wire [0:0] sb_0__2__0_chany_bottom_out_75_;
wire [0:0] sb_0__2__0_chany_bottom_out_77_;
wire [0:0] sb_0__2__0_chany_bottom_out_79_;
wire [0:0] sb_0__2__0_chany_bottom_out_7_;
wire [0:0] sb_0__2__0_chany_bottom_out_81_;
wire [0:0] sb_0__2__0_chany_bottom_out_83_;
wire [0:0] sb_0__2__0_chany_bottom_out_85_;
wire [0:0] sb_0__2__0_chany_bottom_out_87_;
wire [0:0] sb_0__2__0_chany_bottom_out_89_;
wire [0:0] sb_0__2__0_chany_bottom_out_91_;
wire [0:0] sb_0__2__0_chany_bottom_out_93_;
wire [0:0] sb_0__2__0_chany_bottom_out_95_;
wire [0:0] sb_0__2__0_chany_bottom_out_97_;
wire [0:0] sb_0__2__0_chany_bottom_out_99_;
wire [0:0] sb_0__2__0_chany_bottom_out_9_;
wire [0:0] sb_1__0__0_ccff_tail;
wire [0:0] sb_1__0__0_chanx_left_out_101_;
wire [0:0] sb_1__0__0_chanx_left_out_103_;
wire [0:0] sb_1__0__0_chanx_left_out_105_;
wire [0:0] sb_1__0__0_chanx_left_out_107_;
wire [0:0] sb_1__0__0_chanx_left_out_109_;
wire [0:0] sb_1__0__0_chanx_left_out_111_;
wire [0:0] sb_1__0__0_chanx_left_out_113_;
wire [0:0] sb_1__0__0_chanx_left_out_115_;
wire [0:0] sb_1__0__0_chanx_left_out_117_;
wire [0:0] sb_1__0__0_chanx_left_out_119_;
wire [0:0] sb_1__0__0_chanx_left_out_11_;
wire [0:0] sb_1__0__0_chanx_left_out_121_;
wire [0:0] sb_1__0__0_chanx_left_out_123_;
wire [0:0] sb_1__0__0_chanx_left_out_125_;
wire [0:0] sb_1__0__0_chanx_left_out_127_;
wire [0:0] sb_1__0__0_chanx_left_out_129_;
wire [0:0] sb_1__0__0_chanx_left_out_131_;
wire [0:0] sb_1__0__0_chanx_left_out_133_;
wire [0:0] sb_1__0__0_chanx_left_out_135_;
wire [0:0] sb_1__0__0_chanx_left_out_137_;
wire [0:0] sb_1__0__0_chanx_left_out_139_;
wire [0:0] sb_1__0__0_chanx_left_out_13_;
wire [0:0] sb_1__0__0_chanx_left_out_141_;
wire [0:0] sb_1__0__0_chanx_left_out_143_;
wire [0:0] sb_1__0__0_chanx_left_out_145_;
wire [0:0] sb_1__0__0_chanx_left_out_147_;
wire [0:0] sb_1__0__0_chanx_left_out_149_;
wire [0:0] sb_1__0__0_chanx_left_out_151_;
wire [0:0] sb_1__0__0_chanx_left_out_153_;
wire [0:0] sb_1__0__0_chanx_left_out_155_;
wire [0:0] sb_1__0__0_chanx_left_out_157_;
wire [0:0] sb_1__0__0_chanx_left_out_159_;
wire [0:0] sb_1__0__0_chanx_left_out_15_;
wire [0:0] sb_1__0__0_chanx_left_out_161_;
wire [0:0] sb_1__0__0_chanx_left_out_163_;
wire [0:0] sb_1__0__0_chanx_left_out_165_;
wire [0:0] sb_1__0__0_chanx_left_out_167_;
wire [0:0] sb_1__0__0_chanx_left_out_169_;
wire [0:0] sb_1__0__0_chanx_left_out_171_;
wire [0:0] sb_1__0__0_chanx_left_out_173_;
wire [0:0] sb_1__0__0_chanx_left_out_175_;
wire [0:0] sb_1__0__0_chanx_left_out_177_;
wire [0:0] sb_1__0__0_chanx_left_out_179_;
wire [0:0] sb_1__0__0_chanx_left_out_17_;
wire [0:0] sb_1__0__0_chanx_left_out_181_;
wire [0:0] sb_1__0__0_chanx_left_out_183_;
wire [0:0] sb_1__0__0_chanx_left_out_185_;
wire [0:0] sb_1__0__0_chanx_left_out_187_;
wire [0:0] sb_1__0__0_chanx_left_out_189_;
wire [0:0] sb_1__0__0_chanx_left_out_191_;
wire [0:0] sb_1__0__0_chanx_left_out_193_;
wire [0:0] sb_1__0__0_chanx_left_out_195_;
wire [0:0] sb_1__0__0_chanx_left_out_197_;
wire [0:0] sb_1__0__0_chanx_left_out_199_;
wire [0:0] sb_1__0__0_chanx_left_out_19_;
wire [0:0] sb_1__0__0_chanx_left_out_1_;
wire [0:0] sb_1__0__0_chanx_left_out_21_;
wire [0:0] sb_1__0__0_chanx_left_out_23_;
wire [0:0] sb_1__0__0_chanx_left_out_25_;
wire [0:0] sb_1__0__0_chanx_left_out_27_;
wire [0:0] sb_1__0__0_chanx_left_out_29_;
wire [0:0] sb_1__0__0_chanx_left_out_31_;
wire [0:0] sb_1__0__0_chanx_left_out_33_;
wire [0:0] sb_1__0__0_chanx_left_out_35_;
wire [0:0] sb_1__0__0_chanx_left_out_37_;
wire [0:0] sb_1__0__0_chanx_left_out_39_;
wire [0:0] sb_1__0__0_chanx_left_out_3_;
wire [0:0] sb_1__0__0_chanx_left_out_41_;
wire [0:0] sb_1__0__0_chanx_left_out_43_;
wire [0:0] sb_1__0__0_chanx_left_out_45_;
wire [0:0] sb_1__0__0_chanx_left_out_47_;
wire [0:0] sb_1__0__0_chanx_left_out_49_;
wire [0:0] sb_1__0__0_chanx_left_out_51_;
wire [0:0] sb_1__0__0_chanx_left_out_53_;
wire [0:0] sb_1__0__0_chanx_left_out_55_;
wire [0:0] sb_1__0__0_chanx_left_out_57_;
wire [0:0] sb_1__0__0_chanx_left_out_59_;
wire [0:0] sb_1__0__0_chanx_left_out_5_;
wire [0:0] sb_1__0__0_chanx_left_out_61_;
wire [0:0] sb_1__0__0_chanx_left_out_63_;
wire [0:0] sb_1__0__0_chanx_left_out_65_;
wire [0:0] sb_1__0__0_chanx_left_out_67_;
wire [0:0] sb_1__0__0_chanx_left_out_69_;
wire [0:0] sb_1__0__0_chanx_left_out_71_;
wire [0:0] sb_1__0__0_chanx_left_out_73_;
wire [0:0] sb_1__0__0_chanx_left_out_75_;
wire [0:0] sb_1__0__0_chanx_left_out_77_;
wire [0:0] sb_1__0__0_chanx_left_out_79_;
wire [0:0] sb_1__0__0_chanx_left_out_7_;
wire [0:0] sb_1__0__0_chanx_left_out_81_;
wire [0:0] sb_1__0__0_chanx_left_out_83_;
wire [0:0] sb_1__0__0_chanx_left_out_85_;
wire [0:0] sb_1__0__0_chanx_left_out_87_;
wire [0:0] sb_1__0__0_chanx_left_out_89_;
wire [0:0] sb_1__0__0_chanx_left_out_91_;
wire [0:0] sb_1__0__0_chanx_left_out_93_;
wire [0:0] sb_1__0__0_chanx_left_out_95_;
wire [0:0] sb_1__0__0_chanx_left_out_97_;
wire [0:0] sb_1__0__0_chanx_left_out_99_;
wire [0:0] sb_1__0__0_chanx_left_out_9_;
wire [0:0] sb_1__0__0_chanx_right_out_0_;
wire [0:0] sb_1__0__0_chanx_right_out_100_;
wire [0:0] sb_1__0__0_chanx_right_out_102_;
wire [0:0] sb_1__0__0_chanx_right_out_104_;
wire [0:0] sb_1__0__0_chanx_right_out_106_;
wire [0:0] sb_1__0__0_chanx_right_out_108_;
wire [0:0] sb_1__0__0_chanx_right_out_10_;
wire [0:0] sb_1__0__0_chanx_right_out_110_;
wire [0:0] sb_1__0__0_chanx_right_out_112_;
wire [0:0] sb_1__0__0_chanx_right_out_114_;
wire [0:0] sb_1__0__0_chanx_right_out_116_;
wire [0:0] sb_1__0__0_chanx_right_out_118_;
wire [0:0] sb_1__0__0_chanx_right_out_120_;
wire [0:0] sb_1__0__0_chanx_right_out_122_;
wire [0:0] sb_1__0__0_chanx_right_out_124_;
wire [0:0] sb_1__0__0_chanx_right_out_126_;
wire [0:0] sb_1__0__0_chanx_right_out_128_;
wire [0:0] sb_1__0__0_chanx_right_out_12_;
wire [0:0] sb_1__0__0_chanx_right_out_130_;
wire [0:0] sb_1__0__0_chanx_right_out_132_;
wire [0:0] sb_1__0__0_chanx_right_out_134_;
wire [0:0] sb_1__0__0_chanx_right_out_136_;
wire [0:0] sb_1__0__0_chanx_right_out_138_;
wire [0:0] sb_1__0__0_chanx_right_out_140_;
wire [0:0] sb_1__0__0_chanx_right_out_142_;
wire [0:0] sb_1__0__0_chanx_right_out_144_;
wire [0:0] sb_1__0__0_chanx_right_out_146_;
wire [0:0] sb_1__0__0_chanx_right_out_148_;
wire [0:0] sb_1__0__0_chanx_right_out_14_;
wire [0:0] sb_1__0__0_chanx_right_out_150_;
wire [0:0] sb_1__0__0_chanx_right_out_152_;
wire [0:0] sb_1__0__0_chanx_right_out_154_;
wire [0:0] sb_1__0__0_chanx_right_out_156_;
wire [0:0] sb_1__0__0_chanx_right_out_158_;
wire [0:0] sb_1__0__0_chanx_right_out_160_;
wire [0:0] sb_1__0__0_chanx_right_out_162_;
wire [0:0] sb_1__0__0_chanx_right_out_164_;
wire [0:0] sb_1__0__0_chanx_right_out_166_;
wire [0:0] sb_1__0__0_chanx_right_out_168_;
wire [0:0] sb_1__0__0_chanx_right_out_16_;
wire [0:0] sb_1__0__0_chanx_right_out_170_;
wire [0:0] sb_1__0__0_chanx_right_out_172_;
wire [0:0] sb_1__0__0_chanx_right_out_174_;
wire [0:0] sb_1__0__0_chanx_right_out_176_;
wire [0:0] sb_1__0__0_chanx_right_out_178_;
wire [0:0] sb_1__0__0_chanx_right_out_180_;
wire [0:0] sb_1__0__0_chanx_right_out_182_;
wire [0:0] sb_1__0__0_chanx_right_out_184_;
wire [0:0] sb_1__0__0_chanx_right_out_186_;
wire [0:0] sb_1__0__0_chanx_right_out_188_;
wire [0:0] sb_1__0__0_chanx_right_out_18_;
wire [0:0] sb_1__0__0_chanx_right_out_190_;
wire [0:0] sb_1__0__0_chanx_right_out_192_;
wire [0:0] sb_1__0__0_chanx_right_out_194_;
wire [0:0] sb_1__0__0_chanx_right_out_196_;
wire [0:0] sb_1__0__0_chanx_right_out_198_;
wire [0:0] sb_1__0__0_chanx_right_out_20_;
wire [0:0] sb_1__0__0_chanx_right_out_22_;
wire [0:0] sb_1__0__0_chanx_right_out_24_;
wire [0:0] sb_1__0__0_chanx_right_out_26_;
wire [0:0] sb_1__0__0_chanx_right_out_28_;
wire [0:0] sb_1__0__0_chanx_right_out_2_;
wire [0:0] sb_1__0__0_chanx_right_out_30_;
wire [0:0] sb_1__0__0_chanx_right_out_32_;
wire [0:0] sb_1__0__0_chanx_right_out_34_;
wire [0:0] sb_1__0__0_chanx_right_out_36_;
wire [0:0] sb_1__0__0_chanx_right_out_38_;
wire [0:0] sb_1__0__0_chanx_right_out_40_;
wire [0:0] sb_1__0__0_chanx_right_out_42_;
wire [0:0] sb_1__0__0_chanx_right_out_44_;
wire [0:0] sb_1__0__0_chanx_right_out_46_;
wire [0:0] sb_1__0__0_chanx_right_out_48_;
wire [0:0] sb_1__0__0_chanx_right_out_4_;
wire [0:0] sb_1__0__0_chanx_right_out_50_;
wire [0:0] sb_1__0__0_chanx_right_out_52_;
wire [0:0] sb_1__0__0_chanx_right_out_54_;
wire [0:0] sb_1__0__0_chanx_right_out_56_;
wire [0:0] sb_1__0__0_chanx_right_out_58_;
wire [0:0] sb_1__0__0_chanx_right_out_60_;
wire [0:0] sb_1__0__0_chanx_right_out_62_;
wire [0:0] sb_1__0__0_chanx_right_out_64_;
wire [0:0] sb_1__0__0_chanx_right_out_66_;
wire [0:0] sb_1__0__0_chanx_right_out_68_;
wire [0:0] sb_1__0__0_chanx_right_out_6_;
wire [0:0] sb_1__0__0_chanx_right_out_70_;
wire [0:0] sb_1__0__0_chanx_right_out_72_;
wire [0:0] sb_1__0__0_chanx_right_out_74_;
wire [0:0] sb_1__0__0_chanx_right_out_76_;
wire [0:0] sb_1__0__0_chanx_right_out_78_;
wire [0:0] sb_1__0__0_chanx_right_out_80_;
wire [0:0] sb_1__0__0_chanx_right_out_82_;
wire [0:0] sb_1__0__0_chanx_right_out_84_;
wire [0:0] sb_1__0__0_chanx_right_out_86_;
wire [0:0] sb_1__0__0_chanx_right_out_88_;
wire [0:0] sb_1__0__0_chanx_right_out_8_;
wire [0:0] sb_1__0__0_chanx_right_out_90_;
wire [0:0] sb_1__0__0_chanx_right_out_92_;
wire [0:0] sb_1__0__0_chanx_right_out_94_;
wire [0:0] sb_1__0__0_chanx_right_out_96_;
wire [0:0] sb_1__0__0_chanx_right_out_98_;
wire [0:0] sb_1__0__0_chany_top_out_0_;
wire [0:0] sb_1__0__0_chany_top_out_100_;
wire [0:0] sb_1__0__0_chany_top_out_102_;
wire [0:0] sb_1__0__0_chany_top_out_104_;
wire [0:0] sb_1__0__0_chany_top_out_106_;
wire [0:0] sb_1__0__0_chany_top_out_108_;
wire [0:0] sb_1__0__0_chany_top_out_10_;
wire [0:0] sb_1__0__0_chany_top_out_110_;
wire [0:0] sb_1__0__0_chany_top_out_112_;
wire [0:0] sb_1__0__0_chany_top_out_114_;
wire [0:0] sb_1__0__0_chany_top_out_116_;
wire [0:0] sb_1__0__0_chany_top_out_118_;
wire [0:0] sb_1__0__0_chany_top_out_120_;
wire [0:0] sb_1__0__0_chany_top_out_122_;
wire [0:0] sb_1__0__0_chany_top_out_124_;
wire [0:0] sb_1__0__0_chany_top_out_126_;
wire [0:0] sb_1__0__0_chany_top_out_128_;
wire [0:0] sb_1__0__0_chany_top_out_12_;
wire [0:0] sb_1__0__0_chany_top_out_130_;
wire [0:0] sb_1__0__0_chany_top_out_132_;
wire [0:0] sb_1__0__0_chany_top_out_134_;
wire [0:0] sb_1__0__0_chany_top_out_136_;
wire [0:0] sb_1__0__0_chany_top_out_138_;
wire [0:0] sb_1__0__0_chany_top_out_140_;
wire [0:0] sb_1__0__0_chany_top_out_142_;
wire [0:0] sb_1__0__0_chany_top_out_144_;
wire [0:0] sb_1__0__0_chany_top_out_146_;
wire [0:0] sb_1__0__0_chany_top_out_148_;
wire [0:0] sb_1__0__0_chany_top_out_14_;
wire [0:0] sb_1__0__0_chany_top_out_150_;
wire [0:0] sb_1__0__0_chany_top_out_152_;
wire [0:0] sb_1__0__0_chany_top_out_154_;
wire [0:0] sb_1__0__0_chany_top_out_156_;
wire [0:0] sb_1__0__0_chany_top_out_158_;
wire [0:0] sb_1__0__0_chany_top_out_160_;
wire [0:0] sb_1__0__0_chany_top_out_162_;
wire [0:0] sb_1__0__0_chany_top_out_164_;
wire [0:0] sb_1__0__0_chany_top_out_166_;
wire [0:0] sb_1__0__0_chany_top_out_168_;
wire [0:0] sb_1__0__0_chany_top_out_16_;
wire [0:0] sb_1__0__0_chany_top_out_170_;
wire [0:0] sb_1__0__0_chany_top_out_172_;
wire [0:0] sb_1__0__0_chany_top_out_174_;
wire [0:0] sb_1__0__0_chany_top_out_176_;
wire [0:0] sb_1__0__0_chany_top_out_178_;
wire [0:0] sb_1__0__0_chany_top_out_180_;
wire [0:0] sb_1__0__0_chany_top_out_182_;
wire [0:0] sb_1__0__0_chany_top_out_184_;
wire [0:0] sb_1__0__0_chany_top_out_186_;
wire [0:0] sb_1__0__0_chany_top_out_188_;
wire [0:0] sb_1__0__0_chany_top_out_18_;
wire [0:0] sb_1__0__0_chany_top_out_190_;
wire [0:0] sb_1__0__0_chany_top_out_192_;
wire [0:0] sb_1__0__0_chany_top_out_194_;
wire [0:0] sb_1__0__0_chany_top_out_196_;
wire [0:0] sb_1__0__0_chany_top_out_198_;
wire [0:0] sb_1__0__0_chany_top_out_20_;
wire [0:0] sb_1__0__0_chany_top_out_22_;
wire [0:0] sb_1__0__0_chany_top_out_24_;
wire [0:0] sb_1__0__0_chany_top_out_26_;
wire [0:0] sb_1__0__0_chany_top_out_28_;
wire [0:0] sb_1__0__0_chany_top_out_2_;
wire [0:0] sb_1__0__0_chany_top_out_30_;
wire [0:0] sb_1__0__0_chany_top_out_32_;
wire [0:0] sb_1__0__0_chany_top_out_34_;
wire [0:0] sb_1__0__0_chany_top_out_36_;
wire [0:0] sb_1__0__0_chany_top_out_38_;
wire [0:0] sb_1__0__0_chany_top_out_40_;
wire [0:0] sb_1__0__0_chany_top_out_42_;
wire [0:0] sb_1__0__0_chany_top_out_44_;
wire [0:0] sb_1__0__0_chany_top_out_46_;
wire [0:0] sb_1__0__0_chany_top_out_48_;
wire [0:0] sb_1__0__0_chany_top_out_4_;
wire [0:0] sb_1__0__0_chany_top_out_50_;
wire [0:0] sb_1__0__0_chany_top_out_52_;
wire [0:0] sb_1__0__0_chany_top_out_54_;
wire [0:0] sb_1__0__0_chany_top_out_56_;
wire [0:0] sb_1__0__0_chany_top_out_58_;
wire [0:0] sb_1__0__0_chany_top_out_60_;
wire [0:0] sb_1__0__0_chany_top_out_62_;
wire [0:0] sb_1__0__0_chany_top_out_64_;
wire [0:0] sb_1__0__0_chany_top_out_66_;
wire [0:0] sb_1__0__0_chany_top_out_68_;
wire [0:0] sb_1__0__0_chany_top_out_6_;
wire [0:0] sb_1__0__0_chany_top_out_70_;
wire [0:0] sb_1__0__0_chany_top_out_72_;
wire [0:0] sb_1__0__0_chany_top_out_74_;
wire [0:0] sb_1__0__0_chany_top_out_76_;
wire [0:0] sb_1__0__0_chany_top_out_78_;
wire [0:0] sb_1__0__0_chany_top_out_80_;
wire [0:0] sb_1__0__0_chany_top_out_82_;
wire [0:0] sb_1__0__0_chany_top_out_84_;
wire [0:0] sb_1__0__0_chany_top_out_86_;
wire [0:0] sb_1__0__0_chany_top_out_88_;
wire [0:0] sb_1__0__0_chany_top_out_8_;
wire [0:0] sb_1__0__0_chany_top_out_90_;
wire [0:0] sb_1__0__0_chany_top_out_92_;
wire [0:0] sb_1__0__0_chany_top_out_94_;
wire [0:0] sb_1__0__0_chany_top_out_96_;
wire [0:0] sb_1__0__0_chany_top_out_98_;
wire [0:0] sb_1__1__0_ccff_tail;
wire [0:0] sb_1__1__0_chanx_left_out_101_;
wire [0:0] sb_1__1__0_chanx_left_out_103_;
wire [0:0] sb_1__1__0_chanx_left_out_105_;
wire [0:0] sb_1__1__0_chanx_left_out_107_;
wire [0:0] sb_1__1__0_chanx_left_out_109_;
wire [0:0] sb_1__1__0_chanx_left_out_111_;
wire [0:0] sb_1__1__0_chanx_left_out_113_;
wire [0:0] sb_1__1__0_chanx_left_out_115_;
wire [0:0] sb_1__1__0_chanx_left_out_117_;
wire [0:0] sb_1__1__0_chanx_left_out_119_;
wire [0:0] sb_1__1__0_chanx_left_out_11_;
wire [0:0] sb_1__1__0_chanx_left_out_121_;
wire [0:0] sb_1__1__0_chanx_left_out_123_;
wire [0:0] sb_1__1__0_chanx_left_out_125_;
wire [0:0] sb_1__1__0_chanx_left_out_127_;
wire [0:0] sb_1__1__0_chanx_left_out_129_;
wire [0:0] sb_1__1__0_chanx_left_out_131_;
wire [0:0] sb_1__1__0_chanx_left_out_133_;
wire [0:0] sb_1__1__0_chanx_left_out_135_;
wire [0:0] sb_1__1__0_chanx_left_out_137_;
wire [0:0] sb_1__1__0_chanx_left_out_139_;
wire [0:0] sb_1__1__0_chanx_left_out_13_;
wire [0:0] sb_1__1__0_chanx_left_out_141_;
wire [0:0] sb_1__1__0_chanx_left_out_143_;
wire [0:0] sb_1__1__0_chanx_left_out_145_;
wire [0:0] sb_1__1__0_chanx_left_out_147_;
wire [0:0] sb_1__1__0_chanx_left_out_149_;
wire [0:0] sb_1__1__0_chanx_left_out_151_;
wire [0:0] sb_1__1__0_chanx_left_out_153_;
wire [0:0] sb_1__1__0_chanx_left_out_155_;
wire [0:0] sb_1__1__0_chanx_left_out_157_;
wire [0:0] sb_1__1__0_chanx_left_out_159_;
wire [0:0] sb_1__1__0_chanx_left_out_15_;
wire [0:0] sb_1__1__0_chanx_left_out_161_;
wire [0:0] sb_1__1__0_chanx_left_out_163_;
wire [0:0] sb_1__1__0_chanx_left_out_165_;
wire [0:0] sb_1__1__0_chanx_left_out_167_;
wire [0:0] sb_1__1__0_chanx_left_out_169_;
wire [0:0] sb_1__1__0_chanx_left_out_171_;
wire [0:0] sb_1__1__0_chanx_left_out_173_;
wire [0:0] sb_1__1__0_chanx_left_out_175_;
wire [0:0] sb_1__1__0_chanx_left_out_177_;
wire [0:0] sb_1__1__0_chanx_left_out_179_;
wire [0:0] sb_1__1__0_chanx_left_out_17_;
wire [0:0] sb_1__1__0_chanx_left_out_181_;
wire [0:0] sb_1__1__0_chanx_left_out_183_;
wire [0:0] sb_1__1__0_chanx_left_out_185_;
wire [0:0] sb_1__1__0_chanx_left_out_187_;
wire [0:0] sb_1__1__0_chanx_left_out_189_;
wire [0:0] sb_1__1__0_chanx_left_out_191_;
wire [0:0] sb_1__1__0_chanx_left_out_193_;
wire [0:0] sb_1__1__0_chanx_left_out_195_;
wire [0:0] sb_1__1__0_chanx_left_out_197_;
wire [0:0] sb_1__1__0_chanx_left_out_199_;
wire [0:0] sb_1__1__0_chanx_left_out_19_;
wire [0:0] sb_1__1__0_chanx_left_out_1_;
wire [0:0] sb_1__1__0_chanx_left_out_21_;
wire [0:0] sb_1__1__0_chanx_left_out_23_;
wire [0:0] sb_1__1__0_chanx_left_out_25_;
wire [0:0] sb_1__1__0_chanx_left_out_27_;
wire [0:0] sb_1__1__0_chanx_left_out_29_;
wire [0:0] sb_1__1__0_chanx_left_out_31_;
wire [0:0] sb_1__1__0_chanx_left_out_33_;
wire [0:0] sb_1__1__0_chanx_left_out_35_;
wire [0:0] sb_1__1__0_chanx_left_out_37_;
wire [0:0] sb_1__1__0_chanx_left_out_39_;
wire [0:0] sb_1__1__0_chanx_left_out_3_;
wire [0:0] sb_1__1__0_chanx_left_out_41_;
wire [0:0] sb_1__1__0_chanx_left_out_43_;
wire [0:0] sb_1__1__0_chanx_left_out_45_;
wire [0:0] sb_1__1__0_chanx_left_out_47_;
wire [0:0] sb_1__1__0_chanx_left_out_49_;
wire [0:0] sb_1__1__0_chanx_left_out_51_;
wire [0:0] sb_1__1__0_chanx_left_out_53_;
wire [0:0] sb_1__1__0_chanx_left_out_55_;
wire [0:0] sb_1__1__0_chanx_left_out_57_;
wire [0:0] sb_1__1__0_chanx_left_out_59_;
wire [0:0] sb_1__1__0_chanx_left_out_5_;
wire [0:0] sb_1__1__0_chanx_left_out_61_;
wire [0:0] sb_1__1__0_chanx_left_out_63_;
wire [0:0] sb_1__1__0_chanx_left_out_65_;
wire [0:0] sb_1__1__0_chanx_left_out_67_;
wire [0:0] sb_1__1__0_chanx_left_out_69_;
wire [0:0] sb_1__1__0_chanx_left_out_71_;
wire [0:0] sb_1__1__0_chanx_left_out_73_;
wire [0:0] sb_1__1__0_chanx_left_out_75_;
wire [0:0] sb_1__1__0_chanx_left_out_77_;
wire [0:0] sb_1__1__0_chanx_left_out_79_;
wire [0:0] sb_1__1__0_chanx_left_out_7_;
wire [0:0] sb_1__1__0_chanx_left_out_81_;
wire [0:0] sb_1__1__0_chanx_left_out_83_;
wire [0:0] sb_1__1__0_chanx_left_out_85_;
wire [0:0] sb_1__1__0_chanx_left_out_87_;
wire [0:0] sb_1__1__0_chanx_left_out_89_;
wire [0:0] sb_1__1__0_chanx_left_out_91_;
wire [0:0] sb_1__1__0_chanx_left_out_93_;
wire [0:0] sb_1__1__0_chanx_left_out_95_;
wire [0:0] sb_1__1__0_chanx_left_out_97_;
wire [0:0] sb_1__1__0_chanx_left_out_99_;
wire [0:0] sb_1__1__0_chanx_left_out_9_;
wire [0:0] sb_1__1__0_chanx_right_out_0_;
wire [0:0] sb_1__1__0_chanx_right_out_100_;
wire [0:0] sb_1__1__0_chanx_right_out_102_;
wire [0:0] sb_1__1__0_chanx_right_out_104_;
wire [0:0] sb_1__1__0_chanx_right_out_106_;
wire [0:0] sb_1__1__0_chanx_right_out_108_;
wire [0:0] sb_1__1__0_chanx_right_out_10_;
wire [0:0] sb_1__1__0_chanx_right_out_110_;
wire [0:0] sb_1__1__0_chanx_right_out_112_;
wire [0:0] sb_1__1__0_chanx_right_out_114_;
wire [0:0] sb_1__1__0_chanx_right_out_116_;
wire [0:0] sb_1__1__0_chanx_right_out_118_;
wire [0:0] sb_1__1__0_chanx_right_out_120_;
wire [0:0] sb_1__1__0_chanx_right_out_122_;
wire [0:0] sb_1__1__0_chanx_right_out_124_;
wire [0:0] sb_1__1__0_chanx_right_out_126_;
wire [0:0] sb_1__1__0_chanx_right_out_128_;
wire [0:0] sb_1__1__0_chanx_right_out_12_;
wire [0:0] sb_1__1__0_chanx_right_out_130_;
wire [0:0] sb_1__1__0_chanx_right_out_132_;
wire [0:0] sb_1__1__0_chanx_right_out_134_;
wire [0:0] sb_1__1__0_chanx_right_out_136_;
wire [0:0] sb_1__1__0_chanx_right_out_138_;
wire [0:0] sb_1__1__0_chanx_right_out_140_;
wire [0:0] sb_1__1__0_chanx_right_out_142_;
wire [0:0] sb_1__1__0_chanx_right_out_144_;
wire [0:0] sb_1__1__0_chanx_right_out_146_;
wire [0:0] sb_1__1__0_chanx_right_out_148_;
wire [0:0] sb_1__1__0_chanx_right_out_14_;
wire [0:0] sb_1__1__0_chanx_right_out_150_;
wire [0:0] sb_1__1__0_chanx_right_out_152_;
wire [0:0] sb_1__1__0_chanx_right_out_154_;
wire [0:0] sb_1__1__0_chanx_right_out_156_;
wire [0:0] sb_1__1__0_chanx_right_out_158_;
wire [0:0] sb_1__1__0_chanx_right_out_160_;
wire [0:0] sb_1__1__0_chanx_right_out_162_;
wire [0:0] sb_1__1__0_chanx_right_out_164_;
wire [0:0] sb_1__1__0_chanx_right_out_166_;
wire [0:0] sb_1__1__0_chanx_right_out_168_;
wire [0:0] sb_1__1__0_chanx_right_out_16_;
wire [0:0] sb_1__1__0_chanx_right_out_170_;
wire [0:0] sb_1__1__0_chanx_right_out_172_;
wire [0:0] sb_1__1__0_chanx_right_out_174_;
wire [0:0] sb_1__1__0_chanx_right_out_176_;
wire [0:0] sb_1__1__0_chanx_right_out_178_;
wire [0:0] sb_1__1__0_chanx_right_out_180_;
wire [0:0] sb_1__1__0_chanx_right_out_182_;
wire [0:0] sb_1__1__0_chanx_right_out_184_;
wire [0:0] sb_1__1__0_chanx_right_out_186_;
wire [0:0] sb_1__1__0_chanx_right_out_188_;
wire [0:0] sb_1__1__0_chanx_right_out_18_;
wire [0:0] sb_1__1__0_chanx_right_out_190_;
wire [0:0] sb_1__1__0_chanx_right_out_192_;
wire [0:0] sb_1__1__0_chanx_right_out_194_;
wire [0:0] sb_1__1__0_chanx_right_out_196_;
wire [0:0] sb_1__1__0_chanx_right_out_198_;
wire [0:0] sb_1__1__0_chanx_right_out_20_;
wire [0:0] sb_1__1__0_chanx_right_out_22_;
wire [0:0] sb_1__1__0_chanx_right_out_24_;
wire [0:0] sb_1__1__0_chanx_right_out_26_;
wire [0:0] sb_1__1__0_chanx_right_out_28_;
wire [0:0] sb_1__1__0_chanx_right_out_2_;
wire [0:0] sb_1__1__0_chanx_right_out_30_;
wire [0:0] sb_1__1__0_chanx_right_out_32_;
wire [0:0] sb_1__1__0_chanx_right_out_34_;
wire [0:0] sb_1__1__0_chanx_right_out_36_;
wire [0:0] sb_1__1__0_chanx_right_out_38_;
wire [0:0] sb_1__1__0_chanx_right_out_40_;
wire [0:0] sb_1__1__0_chanx_right_out_42_;
wire [0:0] sb_1__1__0_chanx_right_out_44_;
wire [0:0] sb_1__1__0_chanx_right_out_46_;
wire [0:0] sb_1__1__0_chanx_right_out_48_;
wire [0:0] sb_1__1__0_chanx_right_out_4_;
wire [0:0] sb_1__1__0_chanx_right_out_50_;
wire [0:0] sb_1__1__0_chanx_right_out_52_;
wire [0:0] sb_1__1__0_chanx_right_out_54_;
wire [0:0] sb_1__1__0_chanx_right_out_56_;
wire [0:0] sb_1__1__0_chanx_right_out_58_;
wire [0:0] sb_1__1__0_chanx_right_out_60_;
wire [0:0] sb_1__1__0_chanx_right_out_62_;
wire [0:0] sb_1__1__0_chanx_right_out_64_;
wire [0:0] sb_1__1__0_chanx_right_out_66_;
wire [0:0] sb_1__1__0_chanx_right_out_68_;
wire [0:0] sb_1__1__0_chanx_right_out_6_;
wire [0:0] sb_1__1__0_chanx_right_out_70_;
wire [0:0] sb_1__1__0_chanx_right_out_72_;
wire [0:0] sb_1__1__0_chanx_right_out_74_;
wire [0:0] sb_1__1__0_chanx_right_out_76_;
wire [0:0] sb_1__1__0_chanx_right_out_78_;
wire [0:0] sb_1__1__0_chanx_right_out_80_;
wire [0:0] sb_1__1__0_chanx_right_out_82_;
wire [0:0] sb_1__1__0_chanx_right_out_84_;
wire [0:0] sb_1__1__0_chanx_right_out_86_;
wire [0:0] sb_1__1__0_chanx_right_out_88_;
wire [0:0] sb_1__1__0_chanx_right_out_8_;
wire [0:0] sb_1__1__0_chanx_right_out_90_;
wire [0:0] sb_1__1__0_chanx_right_out_92_;
wire [0:0] sb_1__1__0_chanx_right_out_94_;
wire [0:0] sb_1__1__0_chanx_right_out_96_;
wire [0:0] sb_1__1__0_chanx_right_out_98_;
wire [0:0] sb_1__1__0_chany_bottom_out_101_;
wire [0:0] sb_1__1__0_chany_bottom_out_103_;
wire [0:0] sb_1__1__0_chany_bottom_out_105_;
wire [0:0] sb_1__1__0_chany_bottom_out_107_;
wire [0:0] sb_1__1__0_chany_bottom_out_109_;
wire [0:0] sb_1__1__0_chany_bottom_out_111_;
wire [0:0] sb_1__1__0_chany_bottom_out_113_;
wire [0:0] sb_1__1__0_chany_bottom_out_115_;
wire [0:0] sb_1__1__0_chany_bottom_out_117_;
wire [0:0] sb_1__1__0_chany_bottom_out_119_;
wire [0:0] sb_1__1__0_chany_bottom_out_11_;
wire [0:0] sb_1__1__0_chany_bottom_out_121_;
wire [0:0] sb_1__1__0_chany_bottom_out_123_;
wire [0:0] sb_1__1__0_chany_bottom_out_125_;
wire [0:0] sb_1__1__0_chany_bottom_out_127_;
wire [0:0] sb_1__1__0_chany_bottom_out_129_;
wire [0:0] sb_1__1__0_chany_bottom_out_131_;
wire [0:0] sb_1__1__0_chany_bottom_out_133_;
wire [0:0] sb_1__1__0_chany_bottom_out_135_;
wire [0:0] sb_1__1__0_chany_bottom_out_137_;
wire [0:0] sb_1__1__0_chany_bottom_out_139_;
wire [0:0] sb_1__1__0_chany_bottom_out_13_;
wire [0:0] sb_1__1__0_chany_bottom_out_141_;
wire [0:0] sb_1__1__0_chany_bottom_out_143_;
wire [0:0] sb_1__1__0_chany_bottom_out_145_;
wire [0:0] sb_1__1__0_chany_bottom_out_147_;
wire [0:0] sb_1__1__0_chany_bottom_out_149_;
wire [0:0] sb_1__1__0_chany_bottom_out_151_;
wire [0:0] sb_1__1__0_chany_bottom_out_153_;
wire [0:0] sb_1__1__0_chany_bottom_out_155_;
wire [0:0] sb_1__1__0_chany_bottom_out_157_;
wire [0:0] sb_1__1__0_chany_bottom_out_159_;
wire [0:0] sb_1__1__0_chany_bottom_out_15_;
wire [0:0] sb_1__1__0_chany_bottom_out_161_;
wire [0:0] sb_1__1__0_chany_bottom_out_163_;
wire [0:0] sb_1__1__0_chany_bottom_out_165_;
wire [0:0] sb_1__1__0_chany_bottom_out_167_;
wire [0:0] sb_1__1__0_chany_bottom_out_169_;
wire [0:0] sb_1__1__0_chany_bottom_out_171_;
wire [0:0] sb_1__1__0_chany_bottom_out_173_;
wire [0:0] sb_1__1__0_chany_bottom_out_175_;
wire [0:0] sb_1__1__0_chany_bottom_out_177_;
wire [0:0] sb_1__1__0_chany_bottom_out_179_;
wire [0:0] sb_1__1__0_chany_bottom_out_17_;
wire [0:0] sb_1__1__0_chany_bottom_out_181_;
wire [0:0] sb_1__1__0_chany_bottom_out_183_;
wire [0:0] sb_1__1__0_chany_bottom_out_185_;
wire [0:0] sb_1__1__0_chany_bottom_out_187_;
wire [0:0] sb_1__1__0_chany_bottom_out_189_;
wire [0:0] sb_1__1__0_chany_bottom_out_191_;
wire [0:0] sb_1__1__0_chany_bottom_out_193_;
wire [0:0] sb_1__1__0_chany_bottom_out_195_;
wire [0:0] sb_1__1__0_chany_bottom_out_197_;
wire [0:0] sb_1__1__0_chany_bottom_out_199_;
wire [0:0] sb_1__1__0_chany_bottom_out_19_;
wire [0:0] sb_1__1__0_chany_bottom_out_1_;
wire [0:0] sb_1__1__0_chany_bottom_out_21_;
wire [0:0] sb_1__1__0_chany_bottom_out_23_;
wire [0:0] sb_1__1__0_chany_bottom_out_25_;
wire [0:0] sb_1__1__0_chany_bottom_out_27_;
wire [0:0] sb_1__1__0_chany_bottom_out_29_;
wire [0:0] sb_1__1__0_chany_bottom_out_31_;
wire [0:0] sb_1__1__0_chany_bottom_out_33_;
wire [0:0] sb_1__1__0_chany_bottom_out_35_;
wire [0:0] sb_1__1__0_chany_bottom_out_37_;
wire [0:0] sb_1__1__0_chany_bottom_out_39_;
wire [0:0] sb_1__1__0_chany_bottom_out_3_;
wire [0:0] sb_1__1__0_chany_bottom_out_41_;
wire [0:0] sb_1__1__0_chany_bottom_out_43_;
wire [0:0] sb_1__1__0_chany_bottom_out_45_;
wire [0:0] sb_1__1__0_chany_bottom_out_47_;
wire [0:0] sb_1__1__0_chany_bottom_out_49_;
wire [0:0] sb_1__1__0_chany_bottom_out_51_;
wire [0:0] sb_1__1__0_chany_bottom_out_53_;
wire [0:0] sb_1__1__0_chany_bottom_out_55_;
wire [0:0] sb_1__1__0_chany_bottom_out_57_;
wire [0:0] sb_1__1__0_chany_bottom_out_59_;
wire [0:0] sb_1__1__0_chany_bottom_out_5_;
wire [0:0] sb_1__1__0_chany_bottom_out_61_;
wire [0:0] sb_1__1__0_chany_bottom_out_63_;
wire [0:0] sb_1__1__0_chany_bottom_out_65_;
wire [0:0] sb_1__1__0_chany_bottom_out_67_;
wire [0:0] sb_1__1__0_chany_bottom_out_69_;
wire [0:0] sb_1__1__0_chany_bottom_out_71_;
wire [0:0] sb_1__1__0_chany_bottom_out_73_;
wire [0:0] sb_1__1__0_chany_bottom_out_75_;
wire [0:0] sb_1__1__0_chany_bottom_out_77_;
wire [0:0] sb_1__1__0_chany_bottom_out_79_;
wire [0:0] sb_1__1__0_chany_bottom_out_7_;
wire [0:0] sb_1__1__0_chany_bottom_out_81_;
wire [0:0] sb_1__1__0_chany_bottom_out_83_;
wire [0:0] sb_1__1__0_chany_bottom_out_85_;
wire [0:0] sb_1__1__0_chany_bottom_out_87_;
wire [0:0] sb_1__1__0_chany_bottom_out_89_;
wire [0:0] sb_1__1__0_chany_bottom_out_91_;
wire [0:0] sb_1__1__0_chany_bottom_out_93_;
wire [0:0] sb_1__1__0_chany_bottom_out_95_;
wire [0:0] sb_1__1__0_chany_bottom_out_97_;
wire [0:0] sb_1__1__0_chany_bottom_out_99_;
wire [0:0] sb_1__1__0_chany_bottom_out_9_;
wire [0:0] sb_1__1__0_chany_top_out_0_;
wire [0:0] sb_1__1__0_chany_top_out_100_;
wire [0:0] sb_1__1__0_chany_top_out_102_;
wire [0:0] sb_1__1__0_chany_top_out_104_;
wire [0:0] sb_1__1__0_chany_top_out_106_;
wire [0:0] sb_1__1__0_chany_top_out_108_;
wire [0:0] sb_1__1__0_chany_top_out_10_;
wire [0:0] sb_1__1__0_chany_top_out_110_;
wire [0:0] sb_1__1__0_chany_top_out_112_;
wire [0:0] sb_1__1__0_chany_top_out_114_;
wire [0:0] sb_1__1__0_chany_top_out_116_;
wire [0:0] sb_1__1__0_chany_top_out_118_;
wire [0:0] sb_1__1__0_chany_top_out_120_;
wire [0:0] sb_1__1__0_chany_top_out_122_;
wire [0:0] sb_1__1__0_chany_top_out_124_;
wire [0:0] sb_1__1__0_chany_top_out_126_;
wire [0:0] sb_1__1__0_chany_top_out_128_;
wire [0:0] sb_1__1__0_chany_top_out_12_;
wire [0:0] sb_1__1__0_chany_top_out_130_;
wire [0:0] sb_1__1__0_chany_top_out_132_;
wire [0:0] sb_1__1__0_chany_top_out_134_;
wire [0:0] sb_1__1__0_chany_top_out_136_;
wire [0:0] sb_1__1__0_chany_top_out_138_;
wire [0:0] sb_1__1__0_chany_top_out_140_;
wire [0:0] sb_1__1__0_chany_top_out_142_;
wire [0:0] sb_1__1__0_chany_top_out_144_;
wire [0:0] sb_1__1__0_chany_top_out_146_;
wire [0:0] sb_1__1__0_chany_top_out_148_;
wire [0:0] sb_1__1__0_chany_top_out_14_;
wire [0:0] sb_1__1__0_chany_top_out_150_;
wire [0:0] sb_1__1__0_chany_top_out_152_;
wire [0:0] sb_1__1__0_chany_top_out_154_;
wire [0:0] sb_1__1__0_chany_top_out_156_;
wire [0:0] sb_1__1__0_chany_top_out_158_;
wire [0:0] sb_1__1__0_chany_top_out_160_;
wire [0:0] sb_1__1__0_chany_top_out_162_;
wire [0:0] sb_1__1__0_chany_top_out_164_;
wire [0:0] sb_1__1__0_chany_top_out_166_;
wire [0:0] sb_1__1__0_chany_top_out_168_;
wire [0:0] sb_1__1__0_chany_top_out_16_;
wire [0:0] sb_1__1__0_chany_top_out_170_;
wire [0:0] sb_1__1__0_chany_top_out_172_;
wire [0:0] sb_1__1__0_chany_top_out_174_;
wire [0:0] sb_1__1__0_chany_top_out_176_;
wire [0:0] sb_1__1__0_chany_top_out_178_;
wire [0:0] sb_1__1__0_chany_top_out_180_;
wire [0:0] sb_1__1__0_chany_top_out_182_;
wire [0:0] sb_1__1__0_chany_top_out_184_;
wire [0:0] sb_1__1__0_chany_top_out_186_;
wire [0:0] sb_1__1__0_chany_top_out_188_;
wire [0:0] sb_1__1__0_chany_top_out_18_;
wire [0:0] sb_1__1__0_chany_top_out_190_;
wire [0:0] sb_1__1__0_chany_top_out_192_;
wire [0:0] sb_1__1__0_chany_top_out_194_;
wire [0:0] sb_1__1__0_chany_top_out_196_;
wire [0:0] sb_1__1__0_chany_top_out_198_;
wire [0:0] sb_1__1__0_chany_top_out_20_;
wire [0:0] sb_1__1__0_chany_top_out_22_;
wire [0:0] sb_1__1__0_chany_top_out_24_;
wire [0:0] sb_1__1__0_chany_top_out_26_;
wire [0:0] sb_1__1__0_chany_top_out_28_;
wire [0:0] sb_1__1__0_chany_top_out_2_;
wire [0:0] sb_1__1__0_chany_top_out_30_;
wire [0:0] sb_1__1__0_chany_top_out_32_;
wire [0:0] sb_1__1__0_chany_top_out_34_;
wire [0:0] sb_1__1__0_chany_top_out_36_;
wire [0:0] sb_1__1__0_chany_top_out_38_;
wire [0:0] sb_1__1__0_chany_top_out_40_;
wire [0:0] sb_1__1__0_chany_top_out_42_;
wire [0:0] sb_1__1__0_chany_top_out_44_;
wire [0:0] sb_1__1__0_chany_top_out_46_;
wire [0:0] sb_1__1__0_chany_top_out_48_;
wire [0:0] sb_1__1__0_chany_top_out_4_;
wire [0:0] sb_1__1__0_chany_top_out_50_;
wire [0:0] sb_1__1__0_chany_top_out_52_;
wire [0:0] sb_1__1__0_chany_top_out_54_;
wire [0:0] sb_1__1__0_chany_top_out_56_;
wire [0:0] sb_1__1__0_chany_top_out_58_;
wire [0:0] sb_1__1__0_chany_top_out_60_;
wire [0:0] sb_1__1__0_chany_top_out_62_;
wire [0:0] sb_1__1__0_chany_top_out_64_;
wire [0:0] sb_1__1__0_chany_top_out_66_;
wire [0:0] sb_1__1__0_chany_top_out_68_;
wire [0:0] sb_1__1__0_chany_top_out_6_;
wire [0:0] sb_1__1__0_chany_top_out_70_;
wire [0:0] sb_1__1__0_chany_top_out_72_;
wire [0:0] sb_1__1__0_chany_top_out_74_;
wire [0:0] sb_1__1__0_chany_top_out_76_;
wire [0:0] sb_1__1__0_chany_top_out_78_;
wire [0:0] sb_1__1__0_chany_top_out_80_;
wire [0:0] sb_1__1__0_chany_top_out_82_;
wire [0:0] sb_1__1__0_chany_top_out_84_;
wire [0:0] sb_1__1__0_chany_top_out_86_;
wire [0:0] sb_1__1__0_chany_top_out_88_;
wire [0:0] sb_1__1__0_chany_top_out_8_;
wire [0:0] sb_1__1__0_chany_top_out_90_;
wire [0:0] sb_1__1__0_chany_top_out_92_;
wire [0:0] sb_1__1__0_chany_top_out_94_;
wire [0:0] sb_1__1__0_chany_top_out_96_;
wire [0:0] sb_1__1__0_chany_top_out_98_;
wire [0:0] sb_1__2__0_ccff_tail;
wire [0:0] sb_1__2__0_chanx_left_out_101_;
wire [0:0] sb_1__2__0_chanx_left_out_103_;
wire [0:0] sb_1__2__0_chanx_left_out_105_;
wire [0:0] sb_1__2__0_chanx_left_out_107_;
wire [0:0] sb_1__2__0_chanx_left_out_109_;
wire [0:0] sb_1__2__0_chanx_left_out_111_;
wire [0:0] sb_1__2__0_chanx_left_out_113_;
wire [0:0] sb_1__2__0_chanx_left_out_115_;
wire [0:0] sb_1__2__0_chanx_left_out_117_;
wire [0:0] sb_1__2__0_chanx_left_out_119_;
wire [0:0] sb_1__2__0_chanx_left_out_11_;
wire [0:0] sb_1__2__0_chanx_left_out_121_;
wire [0:0] sb_1__2__0_chanx_left_out_123_;
wire [0:0] sb_1__2__0_chanx_left_out_125_;
wire [0:0] sb_1__2__0_chanx_left_out_127_;
wire [0:0] sb_1__2__0_chanx_left_out_129_;
wire [0:0] sb_1__2__0_chanx_left_out_131_;
wire [0:0] sb_1__2__0_chanx_left_out_133_;
wire [0:0] sb_1__2__0_chanx_left_out_135_;
wire [0:0] sb_1__2__0_chanx_left_out_137_;
wire [0:0] sb_1__2__0_chanx_left_out_139_;
wire [0:0] sb_1__2__0_chanx_left_out_13_;
wire [0:0] sb_1__2__0_chanx_left_out_141_;
wire [0:0] sb_1__2__0_chanx_left_out_143_;
wire [0:0] sb_1__2__0_chanx_left_out_145_;
wire [0:0] sb_1__2__0_chanx_left_out_147_;
wire [0:0] sb_1__2__0_chanx_left_out_149_;
wire [0:0] sb_1__2__0_chanx_left_out_151_;
wire [0:0] sb_1__2__0_chanx_left_out_153_;
wire [0:0] sb_1__2__0_chanx_left_out_155_;
wire [0:0] sb_1__2__0_chanx_left_out_157_;
wire [0:0] sb_1__2__0_chanx_left_out_159_;
wire [0:0] sb_1__2__0_chanx_left_out_15_;
wire [0:0] sb_1__2__0_chanx_left_out_161_;
wire [0:0] sb_1__2__0_chanx_left_out_163_;
wire [0:0] sb_1__2__0_chanx_left_out_165_;
wire [0:0] sb_1__2__0_chanx_left_out_167_;
wire [0:0] sb_1__2__0_chanx_left_out_169_;
wire [0:0] sb_1__2__0_chanx_left_out_171_;
wire [0:0] sb_1__2__0_chanx_left_out_173_;
wire [0:0] sb_1__2__0_chanx_left_out_175_;
wire [0:0] sb_1__2__0_chanx_left_out_177_;
wire [0:0] sb_1__2__0_chanx_left_out_179_;
wire [0:0] sb_1__2__0_chanx_left_out_17_;
wire [0:0] sb_1__2__0_chanx_left_out_181_;
wire [0:0] sb_1__2__0_chanx_left_out_183_;
wire [0:0] sb_1__2__0_chanx_left_out_185_;
wire [0:0] sb_1__2__0_chanx_left_out_187_;
wire [0:0] sb_1__2__0_chanx_left_out_189_;
wire [0:0] sb_1__2__0_chanx_left_out_191_;
wire [0:0] sb_1__2__0_chanx_left_out_193_;
wire [0:0] sb_1__2__0_chanx_left_out_195_;
wire [0:0] sb_1__2__0_chanx_left_out_197_;
wire [0:0] sb_1__2__0_chanx_left_out_199_;
wire [0:0] sb_1__2__0_chanx_left_out_19_;
wire [0:0] sb_1__2__0_chanx_left_out_1_;
wire [0:0] sb_1__2__0_chanx_left_out_21_;
wire [0:0] sb_1__2__0_chanx_left_out_23_;
wire [0:0] sb_1__2__0_chanx_left_out_25_;
wire [0:0] sb_1__2__0_chanx_left_out_27_;
wire [0:0] sb_1__2__0_chanx_left_out_29_;
wire [0:0] sb_1__2__0_chanx_left_out_31_;
wire [0:0] sb_1__2__0_chanx_left_out_33_;
wire [0:0] sb_1__2__0_chanx_left_out_35_;
wire [0:0] sb_1__2__0_chanx_left_out_37_;
wire [0:0] sb_1__2__0_chanx_left_out_39_;
wire [0:0] sb_1__2__0_chanx_left_out_3_;
wire [0:0] sb_1__2__0_chanx_left_out_41_;
wire [0:0] sb_1__2__0_chanx_left_out_43_;
wire [0:0] sb_1__2__0_chanx_left_out_45_;
wire [0:0] sb_1__2__0_chanx_left_out_47_;
wire [0:0] sb_1__2__0_chanx_left_out_49_;
wire [0:0] sb_1__2__0_chanx_left_out_51_;
wire [0:0] sb_1__2__0_chanx_left_out_53_;
wire [0:0] sb_1__2__0_chanx_left_out_55_;
wire [0:0] sb_1__2__0_chanx_left_out_57_;
wire [0:0] sb_1__2__0_chanx_left_out_59_;
wire [0:0] sb_1__2__0_chanx_left_out_5_;
wire [0:0] sb_1__2__0_chanx_left_out_61_;
wire [0:0] sb_1__2__0_chanx_left_out_63_;
wire [0:0] sb_1__2__0_chanx_left_out_65_;
wire [0:0] sb_1__2__0_chanx_left_out_67_;
wire [0:0] sb_1__2__0_chanx_left_out_69_;
wire [0:0] sb_1__2__0_chanx_left_out_71_;
wire [0:0] sb_1__2__0_chanx_left_out_73_;
wire [0:0] sb_1__2__0_chanx_left_out_75_;
wire [0:0] sb_1__2__0_chanx_left_out_77_;
wire [0:0] sb_1__2__0_chanx_left_out_79_;
wire [0:0] sb_1__2__0_chanx_left_out_7_;
wire [0:0] sb_1__2__0_chanx_left_out_81_;
wire [0:0] sb_1__2__0_chanx_left_out_83_;
wire [0:0] sb_1__2__0_chanx_left_out_85_;
wire [0:0] sb_1__2__0_chanx_left_out_87_;
wire [0:0] sb_1__2__0_chanx_left_out_89_;
wire [0:0] sb_1__2__0_chanx_left_out_91_;
wire [0:0] sb_1__2__0_chanx_left_out_93_;
wire [0:0] sb_1__2__0_chanx_left_out_95_;
wire [0:0] sb_1__2__0_chanx_left_out_97_;
wire [0:0] sb_1__2__0_chanx_left_out_99_;
wire [0:0] sb_1__2__0_chanx_left_out_9_;
wire [0:0] sb_1__2__0_chanx_right_out_0_;
wire [0:0] sb_1__2__0_chanx_right_out_100_;
wire [0:0] sb_1__2__0_chanx_right_out_102_;
wire [0:0] sb_1__2__0_chanx_right_out_104_;
wire [0:0] sb_1__2__0_chanx_right_out_106_;
wire [0:0] sb_1__2__0_chanx_right_out_108_;
wire [0:0] sb_1__2__0_chanx_right_out_10_;
wire [0:0] sb_1__2__0_chanx_right_out_110_;
wire [0:0] sb_1__2__0_chanx_right_out_112_;
wire [0:0] sb_1__2__0_chanx_right_out_114_;
wire [0:0] sb_1__2__0_chanx_right_out_116_;
wire [0:0] sb_1__2__0_chanx_right_out_118_;
wire [0:0] sb_1__2__0_chanx_right_out_120_;
wire [0:0] sb_1__2__0_chanx_right_out_122_;
wire [0:0] sb_1__2__0_chanx_right_out_124_;
wire [0:0] sb_1__2__0_chanx_right_out_126_;
wire [0:0] sb_1__2__0_chanx_right_out_128_;
wire [0:0] sb_1__2__0_chanx_right_out_12_;
wire [0:0] sb_1__2__0_chanx_right_out_130_;
wire [0:0] sb_1__2__0_chanx_right_out_132_;
wire [0:0] sb_1__2__0_chanx_right_out_134_;
wire [0:0] sb_1__2__0_chanx_right_out_136_;
wire [0:0] sb_1__2__0_chanx_right_out_138_;
wire [0:0] sb_1__2__0_chanx_right_out_140_;
wire [0:0] sb_1__2__0_chanx_right_out_142_;
wire [0:0] sb_1__2__0_chanx_right_out_144_;
wire [0:0] sb_1__2__0_chanx_right_out_146_;
wire [0:0] sb_1__2__0_chanx_right_out_148_;
wire [0:0] sb_1__2__0_chanx_right_out_14_;
wire [0:0] sb_1__2__0_chanx_right_out_150_;
wire [0:0] sb_1__2__0_chanx_right_out_152_;
wire [0:0] sb_1__2__0_chanx_right_out_154_;
wire [0:0] sb_1__2__0_chanx_right_out_156_;
wire [0:0] sb_1__2__0_chanx_right_out_158_;
wire [0:0] sb_1__2__0_chanx_right_out_160_;
wire [0:0] sb_1__2__0_chanx_right_out_162_;
wire [0:0] sb_1__2__0_chanx_right_out_164_;
wire [0:0] sb_1__2__0_chanx_right_out_166_;
wire [0:0] sb_1__2__0_chanx_right_out_168_;
wire [0:0] sb_1__2__0_chanx_right_out_16_;
wire [0:0] sb_1__2__0_chanx_right_out_170_;
wire [0:0] sb_1__2__0_chanx_right_out_172_;
wire [0:0] sb_1__2__0_chanx_right_out_174_;
wire [0:0] sb_1__2__0_chanx_right_out_176_;
wire [0:0] sb_1__2__0_chanx_right_out_178_;
wire [0:0] sb_1__2__0_chanx_right_out_180_;
wire [0:0] sb_1__2__0_chanx_right_out_182_;
wire [0:0] sb_1__2__0_chanx_right_out_184_;
wire [0:0] sb_1__2__0_chanx_right_out_186_;
wire [0:0] sb_1__2__0_chanx_right_out_188_;
wire [0:0] sb_1__2__0_chanx_right_out_18_;
wire [0:0] sb_1__2__0_chanx_right_out_190_;
wire [0:0] sb_1__2__0_chanx_right_out_192_;
wire [0:0] sb_1__2__0_chanx_right_out_194_;
wire [0:0] sb_1__2__0_chanx_right_out_196_;
wire [0:0] sb_1__2__0_chanx_right_out_198_;
wire [0:0] sb_1__2__0_chanx_right_out_20_;
wire [0:0] sb_1__2__0_chanx_right_out_22_;
wire [0:0] sb_1__2__0_chanx_right_out_24_;
wire [0:0] sb_1__2__0_chanx_right_out_26_;
wire [0:0] sb_1__2__0_chanx_right_out_28_;
wire [0:0] sb_1__2__0_chanx_right_out_2_;
wire [0:0] sb_1__2__0_chanx_right_out_30_;
wire [0:0] sb_1__2__0_chanx_right_out_32_;
wire [0:0] sb_1__2__0_chanx_right_out_34_;
wire [0:0] sb_1__2__0_chanx_right_out_36_;
wire [0:0] sb_1__2__0_chanx_right_out_38_;
wire [0:0] sb_1__2__0_chanx_right_out_40_;
wire [0:0] sb_1__2__0_chanx_right_out_42_;
wire [0:0] sb_1__2__0_chanx_right_out_44_;
wire [0:0] sb_1__2__0_chanx_right_out_46_;
wire [0:0] sb_1__2__0_chanx_right_out_48_;
wire [0:0] sb_1__2__0_chanx_right_out_4_;
wire [0:0] sb_1__2__0_chanx_right_out_50_;
wire [0:0] sb_1__2__0_chanx_right_out_52_;
wire [0:0] sb_1__2__0_chanx_right_out_54_;
wire [0:0] sb_1__2__0_chanx_right_out_56_;
wire [0:0] sb_1__2__0_chanx_right_out_58_;
wire [0:0] sb_1__2__0_chanx_right_out_60_;
wire [0:0] sb_1__2__0_chanx_right_out_62_;
wire [0:0] sb_1__2__0_chanx_right_out_64_;
wire [0:0] sb_1__2__0_chanx_right_out_66_;
wire [0:0] sb_1__2__0_chanx_right_out_68_;
wire [0:0] sb_1__2__0_chanx_right_out_6_;
wire [0:0] sb_1__2__0_chanx_right_out_70_;
wire [0:0] sb_1__2__0_chanx_right_out_72_;
wire [0:0] sb_1__2__0_chanx_right_out_74_;
wire [0:0] sb_1__2__0_chanx_right_out_76_;
wire [0:0] sb_1__2__0_chanx_right_out_78_;
wire [0:0] sb_1__2__0_chanx_right_out_80_;
wire [0:0] sb_1__2__0_chanx_right_out_82_;
wire [0:0] sb_1__2__0_chanx_right_out_84_;
wire [0:0] sb_1__2__0_chanx_right_out_86_;
wire [0:0] sb_1__2__0_chanx_right_out_88_;
wire [0:0] sb_1__2__0_chanx_right_out_8_;
wire [0:0] sb_1__2__0_chanx_right_out_90_;
wire [0:0] sb_1__2__0_chanx_right_out_92_;
wire [0:0] sb_1__2__0_chanx_right_out_94_;
wire [0:0] sb_1__2__0_chanx_right_out_96_;
wire [0:0] sb_1__2__0_chanx_right_out_98_;
wire [0:0] sb_1__2__0_chany_bottom_out_101_;
wire [0:0] sb_1__2__0_chany_bottom_out_103_;
wire [0:0] sb_1__2__0_chany_bottom_out_105_;
wire [0:0] sb_1__2__0_chany_bottom_out_107_;
wire [0:0] sb_1__2__0_chany_bottom_out_109_;
wire [0:0] sb_1__2__0_chany_bottom_out_111_;
wire [0:0] sb_1__2__0_chany_bottom_out_113_;
wire [0:0] sb_1__2__0_chany_bottom_out_115_;
wire [0:0] sb_1__2__0_chany_bottom_out_117_;
wire [0:0] sb_1__2__0_chany_bottom_out_119_;
wire [0:0] sb_1__2__0_chany_bottom_out_11_;
wire [0:0] sb_1__2__0_chany_bottom_out_121_;
wire [0:0] sb_1__2__0_chany_bottom_out_123_;
wire [0:0] sb_1__2__0_chany_bottom_out_125_;
wire [0:0] sb_1__2__0_chany_bottom_out_127_;
wire [0:0] sb_1__2__0_chany_bottom_out_129_;
wire [0:0] sb_1__2__0_chany_bottom_out_131_;
wire [0:0] sb_1__2__0_chany_bottom_out_133_;
wire [0:0] sb_1__2__0_chany_bottom_out_135_;
wire [0:0] sb_1__2__0_chany_bottom_out_137_;
wire [0:0] sb_1__2__0_chany_bottom_out_139_;
wire [0:0] sb_1__2__0_chany_bottom_out_13_;
wire [0:0] sb_1__2__0_chany_bottom_out_141_;
wire [0:0] sb_1__2__0_chany_bottom_out_143_;
wire [0:0] sb_1__2__0_chany_bottom_out_145_;
wire [0:0] sb_1__2__0_chany_bottom_out_147_;
wire [0:0] sb_1__2__0_chany_bottom_out_149_;
wire [0:0] sb_1__2__0_chany_bottom_out_151_;
wire [0:0] sb_1__2__0_chany_bottom_out_153_;
wire [0:0] sb_1__2__0_chany_bottom_out_155_;
wire [0:0] sb_1__2__0_chany_bottom_out_157_;
wire [0:0] sb_1__2__0_chany_bottom_out_159_;
wire [0:0] sb_1__2__0_chany_bottom_out_15_;
wire [0:0] sb_1__2__0_chany_bottom_out_161_;
wire [0:0] sb_1__2__0_chany_bottom_out_163_;
wire [0:0] sb_1__2__0_chany_bottom_out_165_;
wire [0:0] sb_1__2__0_chany_bottom_out_167_;
wire [0:0] sb_1__2__0_chany_bottom_out_169_;
wire [0:0] sb_1__2__0_chany_bottom_out_171_;
wire [0:0] sb_1__2__0_chany_bottom_out_173_;
wire [0:0] sb_1__2__0_chany_bottom_out_175_;
wire [0:0] sb_1__2__0_chany_bottom_out_177_;
wire [0:0] sb_1__2__0_chany_bottom_out_179_;
wire [0:0] sb_1__2__0_chany_bottom_out_17_;
wire [0:0] sb_1__2__0_chany_bottom_out_181_;
wire [0:0] sb_1__2__0_chany_bottom_out_183_;
wire [0:0] sb_1__2__0_chany_bottom_out_185_;
wire [0:0] sb_1__2__0_chany_bottom_out_187_;
wire [0:0] sb_1__2__0_chany_bottom_out_189_;
wire [0:0] sb_1__2__0_chany_bottom_out_191_;
wire [0:0] sb_1__2__0_chany_bottom_out_193_;
wire [0:0] sb_1__2__0_chany_bottom_out_195_;
wire [0:0] sb_1__2__0_chany_bottom_out_197_;
wire [0:0] sb_1__2__0_chany_bottom_out_199_;
wire [0:0] sb_1__2__0_chany_bottom_out_19_;
wire [0:0] sb_1__2__0_chany_bottom_out_1_;
wire [0:0] sb_1__2__0_chany_bottom_out_21_;
wire [0:0] sb_1__2__0_chany_bottom_out_23_;
wire [0:0] sb_1__2__0_chany_bottom_out_25_;
wire [0:0] sb_1__2__0_chany_bottom_out_27_;
wire [0:0] sb_1__2__0_chany_bottom_out_29_;
wire [0:0] sb_1__2__0_chany_bottom_out_31_;
wire [0:0] sb_1__2__0_chany_bottom_out_33_;
wire [0:0] sb_1__2__0_chany_bottom_out_35_;
wire [0:0] sb_1__2__0_chany_bottom_out_37_;
wire [0:0] sb_1__2__0_chany_bottom_out_39_;
wire [0:0] sb_1__2__0_chany_bottom_out_3_;
wire [0:0] sb_1__2__0_chany_bottom_out_41_;
wire [0:0] sb_1__2__0_chany_bottom_out_43_;
wire [0:0] sb_1__2__0_chany_bottom_out_45_;
wire [0:0] sb_1__2__0_chany_bottom_out_47_;
wire [0:0] sb_1__2__0_chany_bottom_out_49_;
wire [0:0] sb_1__2__0_chany_bottom_out_51_;
wire [0:0] sb_1__2__0_chany_bottom_out_53_;
wire [0:0] sb_1__2__0_chany_bottom_out_55_;
wire [0:0] sb_1__2__0_chany_bottom_out_57_;
wire [0:0] sb_1__2__0_chany_bottom_out_59_;
wire [0:0] sb_1__2__0_chany_bottom_out_5_;
wire [0:0] sb_1__2__0_chany_bottom_out_61_;
wire [0:0] sb_1__2__0_chany_bottom_out_63_;
wire [0:0] sb_1__2__0_chany_bottom_out_65_;
wire [0:0] sb_1__2__0_chany_bottom_out_67_;
wire [0:0] sb_1__2__0_chany_bottom_out_69_;
wire [0:0] sb_1__2__0_chany_bottom_out_71_;
wire [0:0] sb_1__2__0_chany_bottom_out_73_;
wire [0:0] sb_1__2__0_chany_bottom_out_75_;
wire [0:0] sb_1__2__0_chany_bottom_out_77_;
wire [0:0] sb_1__2__0_chany_bottom_out_79_;
wire [0:0] sb_1__2__0_chany_bottom_out_7_;
wire [0:0] sb_1__2__0_chany_bottom_out_81_;
wire [0:0] sb_1__2__0_chany_bottom_out_83_;
wire [0:0] sb_1__2__0_chany_bottom_out_85_;
wire [0:0] sb_1__2__0_chany_bottom_out_87_;
wire [0:0] sb_1__2__0_chany_bottom_out_89_;
wire [0:0] sb_1__2__0_chany_bottom_out_91_;
wire [0:0] sb_1__2__0_chany_bottom_out_93_;
wire [0:0] sb_1__2__0_chany_bottom_out_95_;
wire [0:0] sb_1__2__0_chany_bottom_out_97_;
wire [0:0] sb_1__2__0_chany_bottom_out_99_;
wire [0:0] sb_1__2__0_chany_bottom_out_9_;
wire [0:0] sb_2__0__0_ccff_tail;
wire [0:0] sb_2__0__0_chanx_left_out_101_;
wire [0:0] sb_2__0__0_chanx_left_out_103_;
wire [0:0] sb_2__0__0_chanx_left_out_105_;
wire [0:0] sb_2__0__0_chanx_left_out_107_;
wire [0:0] sb_2__0__0_chanx_left_out_109_;
wire [0:0] sb_2__0__0_chanx_left_out_111_;
wire [0:0] sb_2__0__0_chanx_left_out_113_;
wire [0:0] sb_2__0__0_chanx_left_out_115_;
wire [0:0] sb_2__0__0_chanx_left_out_117_;
wire [0:0] sb_2__0__0_chanx_left_out_119_;
wire [0:0] sb_2__0__0_chanx_left_out_11_;
wire [0:0] sb_2__0__0_chanx_left_out_121_;
wire [0:0] sb_2__0__0_chanx_left_out_123_;
wire [0:0] sb_2__0__0_chanx_left_out_125_;
wire [0:0] sb_2__0__0_chanx_left_out_127_;
wire [0:0] sb_2__0__0_chanx_left_out_129_;
wire [0:0] sb_2__0__0_chanx_left_out_131_;
wire [0:0] sb_2__0__0_chanx_left_out_133_;
wire [0:0] sb_2__0__0_chanx_left_out_135_;
wire [0:0] sb_2__0__0_chanx_left_out_137_;
wire [0:0] sb_2__0__0_chanx_left_out_139_;
wire [0:0] sb_2__0__0_chanx_left_out_13_;
wire [0:0] sb_2__0__0_chanx_left_out_141_;
wire [0:0] sb_2__0__0_chanx_left_out_143_;
wire [0:0] sb_2__0__0_chanx_left_out_145_;
wire [0:0] sb_2__0__0_chanx_left_out_147_;
wire [0:0] sb_2__0__0_chanx_left_out_149_;
wire [0:0] sb_2__0__0_chanx_left_out_151_;
wire [0:0] sb_2__0__0_chanx_left_out_153_;
wire [0:0] sb_2__0__0_chanx_left_out_155_;
wire [0:0] sb_2__0__0_chanx_left_out_157_;
wire [0:0] sb_2__0__0_chanx_left_out_159_;
wire [0:0] sb_2__0__0_chanx_left_out_15_;
wire [0:0] sb_2__0__0_chanx_left_out_161_;
wire [0:0] sb_2__0__0_chanx_left_out_163_;
wire [0:0] sb_2__0__0_chanx_left_out_165_;
wire [0:0] sb_2__0__0_chanx_left_out_167_;
wire [0:0] sb_2__0__0_chanx_left_out_169_;
wire [0:0] sb_2__0__0_chanx_left_out_171_;
wire [0:0] sb_2__0__0_chanx_left_out_173_;
wire [0:0] sb_2__0__0_chanx_left_out_175_;
wire [0:0] sb_2__0__0_chanx_left_out_177_;
wire [0:0] sb_2__0__0_chanx_left_out_179_;
wire [0:0] sb_2__0__0_chanx_left_out_17_;
wire [0:0] sb_2__0__0_chanx_left_out_181_;
wire [0:0] sb_2__0__0_chanx_left_out_183_;
wire [0:0] sb_2__0__0_chanx_left_out_185_;
wire [0:0] sb_2__0__0_chanx_left_out_187_;
wire [0:0] sb_2__0__0_chanx_left_out_189_;
wire [0:0] sb_2__0__0_chanx_left_out_191_;
wire [0:0] sb_2__0__0_chanx_left_out_193_;
wire [0:0] sb_2__0__0_chanx_left_out_195_;
wire [0:0] sb_2__0__0_chanx_left_out_197_;
wire [0:0] sb_2__0__0_chanx_left_out_199_;
wire [0:0] sb_2__0__0_chanx_left_out_19_;
wire [0:0] sb_2__0__0_chanx_left_out_1_;
wire [0:0] sb_2__0__0_chanx_left_out_21_;
wire [0:0] sb_2__0__0_chanx_left_out_23_;
wire [0:0] sb_2__0__0_chanx_left_out_25_;
wire [0:0] sb_2__0__0_chanx_left_out_27_;
wire [0:0] sb_2__0__0_chanx_left_out_29_;
wire [0:0] sb_2__0__0_chanx_left_out_31_;
wire [0:0] sb_2__0__0_chanx_left_out_33_;
wire [0:0] sb_2__0__0_chanx_left_out_35_;
wire [0:0] sb_2__0__0_chanx_left_out_37_;
wire [0:0] sb_2__0__0_chanx_left_out_39_;
wire [0:0] sb_2__0__0_chanx_left_out_3_;
wire [0:0] sb_2__0__0_chanx_left_out_41_;
wire [0:0] sb_2__0__0_chanx_left_out_43_;
wire [0:0] sb_2__0__0_chanx_left_out_45_;
wire [0:0] sb_2__0__0_chanx_left_out_47_;
wire [0:0] sb_2__0__0_chanx_left_out_49_;
wire [0:0] sb_2__0__0_chanx_left_out_51_;
wire [0:0] sb_2__0__0_chanx_left_out_53_;
wire [0:0] sb_2__0__0_chanx_left_out_55_;
wire [0:0] sb_2__0__0_chanx_left_out_57_;
wire [0:0] sb_2__0__0_chanx_left_out_59_;
wire [0:0] sb_2__0__0_chanx_left_out_5_;
wire [0:0] sb_2__0__0_chanx_left_out_61_;
wire [0:0] sb_2__0__0_chanx_left_out_63_;
wire [0:0] sb_2__0__0_chanx_left_out_65_;
wire [0:0] sb_2__0__0_chanx_left_out_67_;
wire [0:0] sb_2__0__0_chanx_left_out_69_;
wire [0:0] sb_2__0__0_chanx_left_out_71_;
wire [0:0] sb_2__0__0_chanx_left_out_73_;
wire [0:0] sb_2__0__0_chanx_left_out_75_;
wire [0:0] sb_2__0__0_chanx_left_out_77_;
wire [0:0] sb_2__0__0_chanx_left_out_79_;
wire [0:0] sb_2__0__0_chanx_left_out_7_;
wire [0:0] sb_2__0__0_chanx_left_out_81_;
wire [0:0] sb_2__0__0_chanx_left_out_83_;
wire [0:0] sb_2__0__0_chanx_left_out_85_;
wire [0:0] sb_2__0__0_chanx_left_out_87_;
wire [0:0] sb_2__0__0_chanx_left_out_89_;
wire [0:0] sb_2__0__0_chanx_left_out_91_;
wire [0:0] sb_2__0__0_chanx_left_out_93_;
wire [0:0] sb_2__0__0_chanx_left_out_95_;
wire [0:0] sb_2__0__0_chanx_left_out_97_;
wire [0:0] sb_2__0__0_chanx_left_out_99_;
wire [0:0] sb_2__0__0_chanx_left_out_9_;
wire [0:0] sb_2__0__0_chany_top_out_0_;
wire [0:0] sb_2__0__0_chany_top_out_100_;
wire [0:0] sb_2__0__0_chany_top_out_102_;
wire [0:0] sb_2__0__0_chany_top_out_104_;
wire [0:0] sb_2__0__0_chany_top_out_106_;
wire [0:0] sb_2__0__0_chany_top_out_108_;
wire [0:0] sb_2__0__0_chany_top_out_10_;
wire [0:0] sb_2__0__0_chany_top_out_110_;
wire [0:0] sb_2__0__0_chany_top_out_112_;
wire [0:0] sb_2__0__0_chany_top_out_114_;
wire [0:0] sb_2__0__0_chany_top_out_116_;
wire [0:0] sb_2__0__0_chany_top_out_118_;
wire [0:0] sb_2__0__0_chany_top_out_120_;
wire [0:0] sb_2__0__0_chany_top_out_122_;
wire [0:0] sb_2__0__0_chany_top_out_124_;
wire [0:0] sb_2__0__0_chany_top_out_126_;
wire [0:0] sb_2__0__0_chany_top_out_128_;
wire [0:0] sb_2__0__0_chany_top_out_12_;
wire [0:0] sb_2__0__0_chany_top_out_130_;
wire [0:0] sb_2__0__0_chany_top_out_132_;
wire [0:0] sb_2__0__0_chany_top_out_134_;
wire [0:0] sb_2__0__0_chany_top_out_136_;
wire [0:0] sb_2__0__0_chany_top_out_138_;
wire [0:0] sb_2__0__0_chany_top_out_140_;
wire [0:0] sb_2__0__0_chany_top_out_142_;
wire [0:0] sb_2__0__0_chany_top_out_144_;
wire [0:0] sb_2__0__0_chany_top_out_146_;
wire [0:0] sb_2__0__0_chany_top_out_148_;
wire [0:0] sb_2__0__0_chany_top_out_14_;
wire [0:0] sb_2__0__0_chany_top_out_150_;
wire [0:0] sb_2__0__0_chany_top_out_152_;
wire [0:0] sb_2__0__0_chany_top_out_154_;
wire [0:0] sb_2__0__0_chany_top_out_156_;
wire [0:0] sb_2__0__0_chany_top_out_158_;
wire [0:0] sb_2__0__0_chany_top_out_160_;
wire [0:0] sb_2__0__0_chany_top_out_162_;
wire [0:0] sb_2__0__0_chany_top_out_164_;
wire [0:0] sb_2__0__0_chany_top_out_166_;
wire [0:0] sb_2__0__0_chany_top_out_168_;
wire [0:0] sb_2__0__0_chany_top_out_16_;
wire [0:0] sb_2__0__0_chany_top_out_170_;
wire [0:0] sb_2__0__0_chany_top_out_172_;
wire [0:0] sb_2__0__0_chany_top_out_174_;
wire [0:0] sb_2__0__0_chany_top_out_176_;
wire [0:0] sb_2__0__0_chany_top_out_178_;
wire [0:0] sb_2__0__0_chany_top_out_180_;
wire [0:0] sb_2__0__0_chany_top_out_182_;
wire [0:0] sb_2__0__0_chany_top_out_184_;
wire [0:0] sb_2__0__0_chany_top_out_186_;
wire [0:0] sb_2__0__0_chany_top_out_188_;
wire [0:0] sb_2__0__0_chany_top_out_18_;
wire [0:0] sb_2__0__0_chany_top_out_190_;
wire [0:0] sb_2__0__0_chany_top_out_192_;
wire [0:0] sb_2__0__0_chany_top_out_194_;
wire [0:0] sb_2__0__0_chany_top_out_196_;
wire [0:0] sb_2__0__0_chany_top_out_198_;
wire [0:0] sb_2__0__0_chany_top_out_20_;
wire [0:0] sb_2__0__0_chany_top_out_22_;
wire [0:0] sb_2__0__0_chany_top_out_24_;
wire [0:0] sb_2__0__0_chany_top_out_26_;
wire [0:0] sb_2__0__0_chany_top_out_28_;
wire [0:0] sb_2__0__0_chany_top_out_2_;
wire [0:0] sb_2__0__0_chany_top_out_30_;
wire [0:0] sb_2__0__0_chany_top_out_32_;
wire [0:0] sb_2__0__0_chany_top_out_34_;
wire [0:0] sb_2__0__0_chany_top_out_36_;
wire [0:0] sb_2__0__0_chany_top_out_38_;
wire [0:0] sb_2__0__0_chany_top_out_40_;
wire [0:0] sb_2__0__0_chany_top_out_42_;
wire [0:0] sb_2__0__0_chany_top_out_44_;
wire [0:0] sb_2__0__0_chany_top_out_46_;
wire [0:0] sb_2__0__0_chany_top_out_48_;
wire [0:0] sb_2__0__0_chany_top_out_4_;
wire [0:0] sb_2__0__0_chany_top_out_50_;
wire [0:0] sb_2__0__0_chany_top_out_52_;
wire [0:0] sb_2__0__0_chany_top_out_54_;
wire [0:0] sb_2__0__0_chany_top_out_56_;
wire [0:0] sb_2__0__0_chany_top_out_58_;
wire [0:0] sb_2__0__0_chany_top_out_60_;
wire [0:0] sb_2__0__0_chany_top_out_62_;
wire [0:0] sb_2__0__0_chany_top_out_64_;
wire [0:0] sb_2__0__0_chany_top_out_66_;
wire [0:0] sb_2__0__0_chany_top_out_68_;
wire [0:0] sb_2__0__0_chany_top_out_6_;
wire [0:0] sb_2__0__0_chany_top_out_70_;
wire [0:0] sb_2__0__0_chany_top_out_72_;
wire [0:0] sb_2__0__0_chany_top_out_74_;
wire [0:0] sb_2__0__0_chany_top_out_76_;
wire [0:0] sb_2__0__0_chany_top_out_78_;
wire [0:0] sb_2__0__0_chany_top_out_80_;
wire [0:0] sb_2__0__0_chany_top_out_82_;
wire [0:0] sb_2__0__0_chany_top_out_84_;
wire [0:0] sb_2__0__0_chany_top_out_86_;
wire [0:0] sb_2__0__0_chany_top_out_88_;
wire [0:0] sb_2__0__0_chany_top_out_8_;
wire [0:0] sb_2__0__0_chany_top_out_90_;
wire [0:0] sb_2__0__0_chany_top_out_92_;
wire [0:0] sb_2__0__0_chany_top_out_94_;
wire [0:0] sb_2__0__0_chany_top_out_96_;
wire [0:0] sb_2__0__0_chany_top_out_98_;
wire [0:0] sb_2__1__0_ccff_tail;
wire [0:0] sb_2__1__0_chanx_left_out_101_;
wire [0:0] sb_2__1__0_chanx_left_out_103_;
wire [0:0] sb_2__1__0_chanx_left_out_105_;
wire [0:0] sb_2__1__0_chanx_left_out_107_;
wire [0:0] sb_2__1__0_chanx_left_out_109_;
wire [0:0] sb_2__1__0_chanx_left_out_111_;
wire [0:0] sb_2__1__0_chanx_left_out_113_;
wire [0:0] sb_2__1__0_chanx_left_out_115_;
wire [0:0] sb_2__1__0_chanx_left_out_117_;
wire [0:0] sb_2__1__0_chanx_left_out_119_;
wire [0:0] sb_2__1__0_chanx_left_out_11_;
wire [0:0] sb_2__1__0_chanx_left_out_121_;
wire [0:0] sb_2__1__0_chanx_left_out_123_;
wire [0:0] sb_2__1__0_chanx_left_out_125_;
wire [0:0] sb_2__1__0_chanx_left_out_127_;
wire [0:0] sb_2__1__0_chanx_left_out_129_;
wire [0:0] sb_2__1__0_chanx_left_out_131_;
wire [0:0] sb_2__1__0_chanx_left_out_133_;
wire [0:0] sb_2__1__0_chanx_left_out_135_;
wire [0:0] sb_2__1__0_chanx_left_out_137_;
wire [0:0] sb_2__1__0_chanx_left_out_139_;
wire [0:0] sb_2__1__0_chanx_left_out_13_;
wire [0:0] sb_2__1__0_chanx_left_out_141_;
wire [0:0] sb_2__1__0_chanx_left_out_143_;
wire [0:0] sb_2__1__0_chanx_left_out_145_;
wire [0:0] sb_2__1__0_chanx_left_out_147_;
wire [0:0] sb_2__1__0_chanx_left_out_149_;
wire [0:0] sb_2__1__0_chanx_left_out_151_;
wire [0:0] sb_2__1__0_chanx_left_out_153_;
wire [0:0] sb_2__1__0_chanx_left_out_155_;
wire [0:0] sb_2__1__0_chanx_left_out_157_;
wire [0:0] sb_2__1__0_chanx_left_out_159_;
wire [0:0] sb_2__1__0_chanx_left_out_15_;
wire [0:0] sb_2__1__0_chanx_left_out_161_;
wire [0:0] sb_2__1__0_chanx_left_out_163_;
wire [0:0] sb_2__1__0_chanx_left_out_165_;
wire [0:0] sb_2__1__0_chanx_left_out_167_;
wire [0:0] sb_2__1__0_chanx_left_out_169_;
wire [0:0] sb_2__1__0_chanx_left_out_171_;
wire [0:0] sb_2__1__0_chanx_left_out_173_;
wire [0:0] sb_2__1__0_chanx_left_out_175_;
wire [0:0] sb_2__1__0_chanx_left_out_177_;
wire [0:0] sb_2__1__0_chanx_left_out_179_;
wire [0:0] sb_2__1__0_chanx_left_out_17_;
wire [0:0] sb_2__1__0_chanx_left_out_181_;
wire [0:0] sb_2__1__0_chanx_left_out_183_;
wire [0:0] sb_2__1__0_chanx_left_out_185_;
wire [0:0] sb_2__1__0_chanx_left_out_187_;
wire [0:0] sb_2__1__0_chanx_left_out_189_;
wire [0:0] sb_2__1__0_chanx_left_out_191_;
wire [0:0] sb_2__1__0_chanx_left_out_193_;
wire [0:0] sb_2__1__0_chanx_left_out_195_;
wire [0:0] sb_2__1__0_chanx_left_out_197_;
wire [0:0] sb_2__1__0_chanx_left_out_199_;
wire [0:0] sb_2__1__0_chanx_left_out_19_;
wire [0:0] sb_2__1__0_chanx_left_out_1_;
wire [0:0] sb_2__1__0_chanx_left_out_21_;
wire [0:0] sb_2__1__0_chanx_left_out_23_;
wire [0:0] sb_2__1__0_chanx_left_out_25_;
wire [0:0] sb_2__1__0_chanx_left_out_27_;
wire [0:0] sb_2__1__0_chanx_left_out_29_;
wire [0:0] sb_2__1__0_chanx_left_out_31_;
wire [0:0] sb_2__1__0_chanx_left_out_33_;
wire [0:0] sb_2__1__0_chanx_left_out_35_;
wire [0:0] sb_2__1__0_chanx_left_out_37_;
wire [0:0] sb_2__1__0_chanx_left_out_39_;
wire [0:0] sb_2__1__0_chanx_left_out_3_;
wire [0:0] sb_2__1__0_chanx_left_out_41_;
wire [0:0] sb_2__1__0_chanx_left_out_43_;
wire [0:0] sb_2__1__0_chanx_left_out_45_;
wire [0:0] sb_2__1__0_chanx_left_out_47_;
wire [0:0] sb_2__1__0_chanx_left_out_49_;
wire [0:0] sb_2__1__0_chanx_left_out_51_;
wire [0:0] sb_2__1__0_chanx_left_out_53_;
wire [0:0] sb_2__1__0_chanx_left_out_55_;
wire [0:0] sb_2__1__0_chanx_left_out_57_;
wire [0:0] sb_2__1__0_chanx_left_out_59_;
wire [0:0] sb_2__1__0_chanx_left_out_5_;
wire [0:0] sb_2__1__0_chanx_left_out_61_;
wire [0:0] sb_2__1__0_chanx_left_out_63_;
wire [0:0] sb_2__1__0_chanx_left_out_65_;
wire [0:0] sb_2__1__0_chanx_left_out_67_;
wire [0:0] sb_2__1__0_chanx_left_out_69_;
wire [0:0] sb_2__1__0_chanx_left_out_71_;
wire [0:0] sb_2__1__0_chanx_left_out_73_;
wire [0:0] sb_2__1__0_chanx_left_out_75_;
wire [0:0] sb_2__1__0_chanx_left_out_77_;
wire [0:0] sb_2__1__0_chanx_left_out_79_;
wire [0:0] sb_2__1__0_chanx_left_out_7_;
wire [0:0] sb_2__1__0_chanx_left_out_81_;
wire [0:0] sb_2__1__0_chanx_left_out_83_;
wire [0:0] sb_2__1__0_chanx_left_out_85_;
wire [0:0] sb_2__1__0_chanx_left_out_87_;
wire [0:0] sb_2__1__0_chanx_left_out_89_;
wire [0:0] sb_2__1__0_chanx_left_out_91_;
wire [0:0] sb_2__1__0_chanx_left_out_93_;
wire [0:0] sb_2__1__0_chanx_left_out_95_;
wire [0:0] sb_2__1__0_chanx_left_out_97_;
wire [0:0] sb_2__1__0_chanx_left_out_99_;
wire [0:0] sb_2__1__0_chanx_left_out_9_;
wire [0:0] sb_2__1__0_chany_bottom_out_101_;
wire [0:0] sb_2__1__0_chany_bottom_out_103_;
wire [0:0] sb_2__1__0_chany_bottom_out_105_;
wire [0:0] sb_2__1__0_chany_bottom_out_107_;
wire [0:0] sb_2__1__0_chany_bottom_out_109_;
wire [0:0] sb_2__1__0_chany_bottom_out_111_;
wire [0:0] sb_2__1__0_chany_bottom_out_113_;
wire [0:0] sb_2__1__0_chany_bottom_out_115_;
wire [0:0] sb_2__1__0_chany_bottom_out_117_;
wire [0:0] sb_2__1__0_chany_bottom_out_119_;
wire [0:0] sb_2__1__0_chany_bottom_out_11_;
wire [0:0] sb_2__1__0_chany_bottom_out_121_;
wire [0:0] sb_2__1__0_chany_bottom_out_123_;
wire [0:0] sb_2__1__0_chany_bottom_out_125_;
wire [0:0] sb_2__1__0_chany_bottom_out_127_;
wire [0:0] sb_2__1__0_chany_bottom_out_129_;
wire [0:0] sb_2__1__0_chany_bottom_out_131_;
wire [0:0] sb_2__1__0_chany_bottom_out_133_;
wire [0:0] sb_2__1__0_chany_bottom_out_135_;
wire [0:0] sb_2__1__0_chany_bottom_out_137_;
wire [0:0] sb_2__1__0_chany_bottom_out_139_;
wire [0:0] sb_2__1__0_chany_bottom_out_13_;
wire [0:0] sb_2__1__0_chany_bottom_out_141_;
wire [0:0] sb_2__1__0_chany_bottom_out_143_;
wire [0:0] sb_2__1__0_chany_bottom_out_145_;
wire [0:0] sb_2__1__0_chany_bottom_out_147_;
wire [0:0] sb_2__1__0_chany_bottom_out_149_;
wire [0:0] sb_2__1__0_chany_bottom_out_151_;
wire [0:0] sb_2__1__0_chany_bottom_out_153_;
wire [0:0] sb_2__1__0_chany_bottom_out_155_;
wire [0:0] sb_2__1__0_chany_bottom_out_157_;
wire [0:0] sb_2__1__0_chany_bottom_out_159_;
wire [0:0] sb_2__1__0_chany_bottom_out_15_;
wire [0:0] sb_2__1__0_chany_bottom_out_161_;
wire [0:0] sb_2__1__0_chany_bottom_out_163_;
wire [0:0] sb_2__1__0_chany_bottom_out_165_;
wire [0:0] sb_2__1__0_chany_bottom_out_167_;
wire [0:0] sb_2__1__0_chany_bottom_out_169_;
wire [0:0] sb_2__1__0_chany_bottom_out_171_;
wire [0:0] sb_2__1__0_chany_bottom_out_173_;
wire [0:0] sb_2__1__0_chany_bottom_out_175_;
wire [0:0] sb_2__1__0_chany_bottom_out_177_;
wire [0:0] sb_2__1__0_chany_bottom_out_179_;
wire [0:0] sb_2__1__0_chany_bottom_out_17_;
wire [0:0] sb_2__1__0_chany_bottom_out_181_;
wire [0:0] sb_2__1__0_chany_bottom_out_183_;
wire [0:0] sb_2__1__0_chany_bottom_out_185_;
wire [0:0] sb_2__1__0_chany_bottom_out_187_;
wire [0:0] sb_2__1__0_chany_bottom_out_189_;
wire [0:0] sb_2__1__0_chany_bottom_out_191_;
wire [0:0] sb_2__1__0_chany_bottom_out_193_;
wire [0:0] sb_2__1__0_chany_bottom_out_195_;
wire [0:0] sb_2__1__0_chany_bottom_out_197_;
wire [0:0] sb_2__1__0_chany_bottom_out_199_;
wire [0:0] sb_2__1__0_chany_bottom_out_19_;
wire [0:0] sb_2__1__0_chany_bottom_out_1_;
wire [0:0] sb_2__1__0_chany_bottom_out_21_;
wire [0:0] sb_2__1__0_chany_bottom_out_23_;
wire [0:0] sb_2__1__0_chany_bottom_out_25_;
wire [0:0] sb_2__1__0_chany_bottom_out_27_;
wire [0:0] sb_2__1__0_chany_bottom_out_29_;
wire [0:0] sb_2__1__0_chany_bottom_out_31_;
wire [0:0] sb_2__1__0_chany_bottom_out_33_;
wire [0:0] sb_2__1__0_chany_bottom_out_35_;
wire [0:0] sb_2__1__0_chany_bottom_out_37_;
wire [0:0] sb_2__1__0_chany_bottom_out_39_;
wire [0:0] sb_2__1__0_chany_bottom_out_3_;
wire [0:0] sb_2__1__0_chany_bottom_out_41_;
wire [0:0] sb_2__1__0_chany_bottom_out_43_;
wire [0:0] sb_2__1__0_chany_bottom_out_45_;
wire [0:0] sb_2__1__0_chany_bottom_out_47_;
wire [0:0] sb_2__1__0_chany_bottom_out_49_;
wire [0:0] sb_2__1__0_chany_bottom_out_51_;
wire [0:0] sb_2__1__0_chany_bottom_out_53_;
wire [0:0] sb_2__1__0_chany_bottom_out_55_;
wire [0:0] sb_2__1__0_chany_bottom_out_57_;
wire [0:0] sb_2__1__0_chany_bottom_out_59_;
wire [0:0] sb_2__1__0_chany_bottom_out_5_;
wire [0:0] sb_2__1__0_chany_bottom_out_61_;
wire [0:0] sb_2__1__0_chany_bottom_out_63_;
wire [0:0] sb_2__1__0_chany_bottom_out_65_;
wire [0:0] sb_2__1__0_chany_bottom_out_67_;
wire [0:0] sb_2__1__0_chany_bottom_out_69_;
wire [0:0] sb_2__1__0_chany_bottom_out_71_;
wire [0:0] sb_2__1__0_chany_bottom_out_73_;
wire [0:0] sb_2__1__0_chany_bottom_out_75_;
wire [0:0] sb_2__1__0_chany_bottom_out_77_;
wire [0:0] sb_2__1__0_chany_bottom_out_79_;
wire [0:0] sb_2__1__0_chany_bottom_out_7_;
wire [0:0] sb_2__1__0_chany_bottom_out_81_;
wire [0:0] sb_2__1__0_chany_bottom_out_83_;
wire [0:0] sb_2__1__0_chany_bottom_out_85_;
wire [0:0] sb_2__1__0_chany_bottom_out_87_;
wire [0:0] sb_2__1__0_chany_bottom_out_89_;
wire [0:0] sb_2__1__0_chany_bottom_out_91_;
wire [0:0] sb_2__1__0_chany_bottom_out_93_;
wire [0:0] sb_2__1__0_chany_bottom_out_95_;
wire [0:0] sb_2__1__0_chany_bottom_out_97_;
wire [0:0] sb_2__1__0_chany_bottom_out_99_;
wire [0:0] sb_2__1__0_chany_bottom_out_9_;
wire [0:0] sb_2__1__0_chany_top_out_0_;
wire [0:0] sb_2__1__0_chany_top_out_100_;
wire [0:0] sb_2__1__0_chany_top_out_102_;
wire [0:0] sb_2__1__0_chany_top_out_104_;
wire [0:0] sb_2__1__0_chany_top_out_106_;
wire [0:0] sb_2__1__0_chany_top_out_108_;
wire [0:0] sb_2__1__0_chany_top_out_10_;
wire [0:0] sb_2__1__0_chany_top_out_110_;
wire [0:0] sb_2__1__0_chany_top_out_112_;
wire [0:0] sb_2__1__0_chany_top_out_114_;
wire [0:0] sb_2__1__0_chany_top_out_116_;
wire [0:0] sb_2__1__0_chany_top_out_118_;
wire [0:0] sb_2__1__0_chany_top_out_120_;
wire [0:0] sb_2__1__0_chany_top_out_122_;
wire [0:0] sb_2__1__0_chany_top_out_124_;
wire [0:0] sb_2__1__0_chany_top_out_126_;
wire [0:0] sb_2__1__0_chany_top_out_128_;
wire [0:0] sb_2__1__0_chany_top_out_12_;
wire [0:0] sb_2__1__0_chany_top_out_130_;
wire [0:0] sb_2__1__0_chany_top_out_132_;
wire [0:0] sb_2__1__0_chany_top_out_134_;
wire [0:0] sb_2__1__0_chany_top_out_136_;
wire [0:0] sb_2__1__0_chany_top_out_138_;
wire [0:0] sb_2__1__0_chany_top_out_140_;
wire [0:0] sb_2__1__0_chany_top_out_142_;
wire [0:0] sb_2__1__0_chany_top_out_144_;
wire [0:0] sb_2__1__0_chany_top_out_146_;
wire [0:0] sb_2__1__0_chany_top_out_148_;
wire [0:0] sb_2__1__0_chany_top_out_14_;
wire [0:0] sb_2__1__0_chany_top_out_150_;
wire [0:0] sb_2__1__0_chany_top_out_152_;
wire [0:0] sb_2__1__0_chany_top_out_154_;
wire [0:0] sb_2__1__0_chany_top_out_156_;
wire [0:0] sb_2__1__0_chany_top_out_158_;
wire [0:0] sb_2__1__0_chany_top_out_160_;
wire [0:0] sb_2__1__0_chany_top_out_162_;
wire [0:0] sb_2__1__0_chany_top_out_164_;
wire [0:0] sb_2__1__0_chany_top_out_166_;
wire [0:0] sb_2__1__0_chany_top_out_168_;
wire [0:0] sb_2__1__0_chany_top_out_16_;
wire [0:0] sb_2__1__0_chany_top_out_170_;
wire [0:0] sb_2__1__0_chany_top_out_172_;
wire [0:0] sb_2__1__0_chany_top_out_174_;
wire [0:0] sb_2__1__0_chany_top_out_176_;
wire [0:0] sb_2__1__0_chany_top_out_178_;
wire [0:0] sb_2__1__0_chany_top_out_180_;
wire [0:0] sb_2__1__0_chany_top_out_182_;
wire [0:0] sb_2__1__0_chany_top_out_184_;
wire [0:0] sb_2__1__0_chany_top_out_186_;
wire [0:0] sb_2__1__0_chany_top_out_188_;
wire [0:0] sb_2__1__0_chany_top_out_18_;
wire [0:0] sb_2__1__0_chany_top_out_190_;
wire [0:0] sb_2__1__0_chany_top_out_192_;
wire [0:0] sb_2__1__0_chany_top_out_194_;
wire [0:0] sb_2__1__0_chany_top_out_196_;
wire [0:0] sb_2__1__0_chany_top_out_198_;
wire [0:0] sb_2__1__0_chany_top_out_20_;
wire [0:0] sb_2__1__0_chany_top_out_22_;
wire [0:0] sb_2__1__0_chany_top_out_24_;
wire [0:0] sb_2__1__0_chany_top_out_26_;
wire [0:0] sb_2__1__0_chany_top_out_28_;
wire [0:0] sb_2__1__0_chany_top_out_2_;
wire [0:0] sb_2__1__0_chany_top_out_30_;
wire [0:0] sb_2__1__0_chany_top_out_32_;
wire [0:0] sb_2__1__0_chany_top_out_34_;
wire [0:0] sb_2__1__0_chany_top_out_36_;
wire [0:0] sb_2__1__0_chany_top_out_38_;
wire [0:0] sb_2__1__0_chany_top_out_40_;
wire [0:0] sb_2__1__0_chany_top_out_42_;
wire [0:0] sb_2__1__0_chany_top_out_44_;
wire [0:0] sb_2__1__0_chany_top_out_46_;
wire [0:0] sb_2__1__0_chany_top_out_48_;
wire [0:0] sb_2__1__0_chany_top_out_4_;
wire [0:0] sb_2__1__0_chany_top_out_50_;
wire [0:0] sb_2__1__0_chany_top_out_52_;
wire [0:0] sb_2__1__0_chany_top_out_54_;
wire [0:0] sb_2__1__0_chany_top_out_56_;
wire [0:0] sb_2__1__0_chany_top_out_58_;
wire [0:0] sb_2__1__0_chany_top_out_60_;
wire [0:0] sb_2__1__0_chany_top_out_62_;
wire [0:0] sb_2__1__0_chany_top_out_64_;
wire [0:0] sb_2__1__0_chany_top_out_66_;
wire [0:0] sb_2__1__0_chany_top_out_68_;
wire [0:0] sb_2__1__0_chany_top_out_6_;
wire [0:0] sb_2__1__0_chany_top_out_70_;
wire [0:0] sb_2__1__0_chany_top_out_72_;
wire [0:0] sb_2__1__0_chany_top_out_74_;
wire [0:0] sb_2__1__0_chany_top_out_76_;
wire [0:0] sb_2__1__0_chany_top_out_78_;
wire [0:0] sb_2__1__0_chany_top_out_80_;
wire [0:0] sb_2__1__0_chany_top_out_82_;
wire [0:0] sb_2__1__0_chany_top_out_84_;
wire [0:0] sb_2__1__0_chany_top_out_86_;
wire [0:0] sb_2__1__0_chany_top_out_88_;
wire [0:0] sb_2__1__0_chany_top_out_8_;
wire [0:0] sb_2__1__0_chany_top_out_90_;
wire [0:0] sb_2__1__0_chany_top_out_92_;
wire [0:0] sb_2__1__0_chany_top_out_94_;
wire [0:0] sb_2__1__0_chany_top_out_96_;
wire [0:0] sb_2__1__0_chany_top_out_98_;
wire [0:0] sb_2__2__0_ccff_tail;
wire [0:0] sb_2__2__0_chanx_left_out_101_;
wire [0:0] sb_2__2__0_chanx_left_out_103_;
wire [0:0] sb_2__2__0_chanx_left_out_105_;
wire [0:0] sb_2__2__0_chanx_left_out_107_;
wire [0:0] sb_2__2__0_chanx_left_out_109_;
wire [0:0] sb_2__2__0_chanx_left_out_111_;
wire [0:0] sb_2__2__0_chanx_left_out_113_;
wire [0:0] sb_2__2__0_chanx_left_out_115_;
wire [0:0] sb_2__2__0_chanx_left_out_117_;
wire [0:0] sb_2__2__0_chanx_left_out_119_;
wire [0:0] sb_2__2__0_chanx_left_out_11_;
wire [0:0] sb_2__2__0_chanx_left_out_121_;
wire [0:0] sb_2__2__0_chanx_left_out_123_;
wire [0:0] sb_2__2__0_chanx_left_out_125_;
wire [0:0] sb_2__2__0_chanx_left_out_127_;
wire [0:0] sb_2__2__0_chanx_left_out_129_;
wire [0:0] sb_2__2__0_chanx_left_out_131_;
wire [0:0] sb_2__2__0_chanx_left_out_133_;
wire [0:0] sb_2__2__0_chanx_left_out_135_;
wire [0:0] sb_2__2__0_chanx_left_out_137_;
wire [0:0] sb_2__2__0_chanx_left_out_139_;
wire [0:0] sb_2__2__0_chanx_left_out_13_;
wire [0:0] sb_2__2__0_chanx_left_out_141_;
wire [0:0] sb_2__2__0_chanx_left_out_143_;
wire [0:0] sb_2__2__0_chanx_left_out_145_;
wire [0:0] sb_2__2__0_chanx_left_out_147_;
wire [0:0] sb_2__2__0_chanx_left_out_149_;
wire [0:0] sb_2__2__0_chanx_left_out_151_;
wire [0:0] sb_2__2__0_chanx_left_out_153_;
wire [0:0] sb_2__2__0_chanx_left_out_155_;
wire [0:0] sb_2__2__0_chanx_left_out_157_;
wire [0:0] sb_2__2__0_chanx_left_out_159_;
wire [0:0] sb_2__2__0_chanx_left_out_15_;
wire [0:0] sb_2__2__0_chanx_left_out_161_;
wire [0:0] sb_2__2__0_chanx_left_out_163_;
wire [0:0] sb_2__2__0_chanx_left_out_165_;
wire [0:0] sb_2__2__0_chanx_left_out_167_;
wire [0:0] sb_2__2__0_chanx_left_out_169_;
wire [0:0] sb_2__2__0_chanx_left_out_171_;
wire [0:0] sb_2__2__0_chanx_left_out_173_;
wire [0:0] sb_2__2__0_chanx_left_out_175_;
wire [0:0] sb_2__2__0_chanx_left_out_177_;
wire [0:0] sb_2__2__0_chanx_left_out_179_;
wire [0:0] sb_2__2__0_chanx_left_out_17_;
wire [0:0] sb_2__2__0_chanx_left_out_181_;
wire [0:0] sb_2__2__0_chanx_left_out_183_;
wire [0:0] sb_2__2__0_chanx_left_out_185_;
wire [0:0] sb_2__2__0_chanx_left_out_187_;
wire [0:0] sb_2__2__0_chanx_left_out_189_;
wire [0:0] sb_2__2__0_chanx_left_out_191_;
wire [0:0] sb_2__2__0_chanx_left_out_193_;
wire [0:0] sb_2__2__0_chanx_left_out_195_;
wire [0:0] sb_2__2__0_chanx_left_out_197_;
wire [0:0] sb_2__2__0_chanx_left_out_199_;
wire [0:0] sb_2__2__0_chanx_left_out_19_;
wire [0:0] sb_2__2__0_chanx_left_out_1_;
wire [0:0] sb_2__2__0_chanx_left_out_21_;
wire [0:0] sb_2__2__0_chanx_left_out_23_;
wire [0:0] sb_2__2__0_chanx_left_out_25_;
wire [0:0] sb_2__2__0_chanx_left_out_27_;
wire [0:0] sb_2__2__0_chanx_left_out_29_;
wire [0:0] sb_2__2__0_chanx_left_out_31_;
wire [0:0] sb_2__2__0_chanx_left_out_33_;
wire [0:0] sb_2__2__0_chanx_left_out_35_;
wire [0:0] sb_2__2__0_chanx_left_out_37_;
wire [0:0] sb_2__2__0_chanx_left_out_39_;
wire [0:0] sb_2__2__0_chanx_left_out_3_;
wire [0:0] sb_2__2__0_chanx_left_out_41_;
wire [0:0] sb_2__2__0_chanx_left_out_43_;
wire [0:0] sb_2__2__0_chanx_left_out_45_;
wire [0:0] sb_2__2__0_chanx_left_out_47_;
wire [0:0] sb_2__2__0_chanx_left_out_49_;
wire [0:0] sb_2__2__0_chanx_left_out_51_;
wire [0:0] sb_2__2__0_chanx_left_out_53_;
wire [0:0] sb_2__2__0_chanx_left_out_55_;
wire [0:0] sb_2__2__0_chanx_left_out_57_;
wire [0:0] sb_2__2__0_chanx_left_out_59_;
wire [0:0] sb_2__2__0_chanx_left_out_5_;
wire [0:0] sb_2__2__0_chanx_left_out_61_;
wire [0:0] sb_2__2__0_chanx_left_out_63_;
wire [0:0] sb_2__2__0_chanx_left_out_65_;
wire [0:0] sb_2__2__0_chanx_left_out_67_;
wire [0:0] sb_2__2__0_chanx_left_out_69_;
wire [0:0] sb_2__2__0_chanx_left_out_71_;
wire [0:0] sb_2__2__0_chanx_left_out_73_;
wire [0:0] sb_2__2__0_chanx_left_out_75_;
wire [0:0] sb_2__2__0_chanx_left_out_77_;
wire [0:0] sb_2__2__0_chanx_left_out_79_;
wire [0:0] sb_2__2__0_chanx_left_out_7_;
wire [0:0] sb_2__2__0_chanx_left_out_81_;
wire [0:0] sb_2__2__0_chanx_left_out_83_;
wire [0:0] sb_2__2__0_chanx_left_out_85_;
wire [0:0] sb_2__2__0_chanx_left_out_87_;
wire [0:0] sb_2__2__0_chanx_left_out_89_;
wire [0:0] sb_2__2__0_chanx_left_out_91_;
wire [0:0] sb_2__2__0_chanx_left_out_93_;
wire [0:0] sb_2__2__0_chanx_left_out_95_;
wire [0:0] sb_2__2__0_chanx_left_out_97_;
wire [0:0] sb_2__2__0_chanx_left_out_99_;
wire [0:0] sb_2__2__0_chanx_left_out_9_;
wire [0:0] sb_2__2__0_chany_bottom_out_101_;
wire [0:0] sb_2__2__0_chany_bottom_out_103_;
wire [0:0] sb_2__2__0_chany_bottom_out_105_;
wire [0:0] sb_2__2__0_chany_bottom_out_107_;
wire [0:0] sb_2__2__0_chany_bottom_out_109_;
wire [0:0] sb_2__2__0_chany_bottom_out_111_;
wire [0:0] sb_2__2__0_chany_bottom_out_113_;
wire [0:0] sb_2__2__0_chany_bottom_out_115_;
wire [0:0] sb_2__2__0_chany_bottom_out_117_;
wire [0:0] sb_2__2__0_chany_bottom_out_119_;
wire [0:0] sb_2__2__0_chany_bottom_out_11_;
wire [0:0] sb_2__2__0_chany_bottom_out_121_;
wire [0:0] sb_2__2__0_chany_bottom_out_123_;
wire [0:0] sb_2__2__0_chany_bottom_out_125_;
wire [0:0] sb_2__2__0_chany_bottom_out_127_;
wire [0:0] sb_2__2__0_chany_bottom_out_129_;
wire [0:0] sb_2__2__0_chany_bottom_out_131_;
wire [0:0] sb_2__2__0_chany_bottom_out_133_;
wire [0:0] sb_2__2__0_chany_bottom_out_135_;
wire [0:0] sb_2__2__0_chany_bottom_out_137_;
wire [0:0] sb_2__2__0_chany_bottom_out_139_;
wire [0:0] sb_2__2__0_chany_bottom_out_13_;
wire [0:0] sb_2__2__0_chany_bottom_out_141_;
wire [0:0] sb_2__2__0_chany_bottom_out_143_;
wire [0:0] sb_2__2__0_chany_bottom_out_145_;
wire [0:0] sb_2__2__0_chany_bottom_out_147_;
wire [0:0] sb_2__2__0_chany_bottom_out_149_;
wire [0:0] sb_2__2__0_chany_bottom_out_151_;
wire [0:0] sb_2__2__0_chany_bottom_out_153_;
wire [0:0] sb_2__2__0_chany_bottom_out_155_;
wire [0:0] sb_2__2__0_chany_bottom_out_157_;
wire [0:0] sb_2__2__0_chany_bottom_out_159_;
wire [0:0] sb_2__2__0_chany_bottom_out_15_;
wire [0:0] sb_2__2__0_chany_bottom_out_161_;
wire [0:0] sb_2__2__0_chany_bottom_out_163_;
wire [0:0] sb_2__2__0_chany_bottom_out_165_;
wire [0:0] sb_2__2__0_chany_bottom_out_167_;
wire [0:0] sb_2__2__0_chany_bottom_out_169_;
wire [0:0] sb_2__2__0_chany_bottom_out_171_;
wire [0:0] sb_2__2__0_chany_bottom_out_173_;
wire [0:0] sb_2__2__0_chany_bottom_out_175_;
wire [0:0] sb_2__2__0_chany_bottom_out_177_;
wire [0:0] sb_2__2__0_chany_bottom_out_179_;
wire [0:0] sb_2__2__0_chany_bottom_out_17_;
wire [0:0] sb_2__2__0_chany_bottom_out_181_;
wire [0:0] sb_2__2__0_chany_bottom_out_183_;
wire [0:0] sb_2__2__0_chany_bottom_out_185_;
wire [0:0] sb_2__2__0_chany_bottom_out_187_;
wire [0:0] sb_2__2__0_chany_bottom_out_189_;
wire [0:0] sb_2__2__0_chany_bottom_out_191_;
wire [0:0] sb_2__2__0_chany_bottom_out_193_;
wire [0:0] sb_2__2__0_chany_bottom_out_195_;
wire [0:0] sb_2__2__0_chany_bottom_out_197_;
wire [0:0] sb_2__2__0_chany_bottom_out_199_;
wire [0:0] sb_2__2__0_chany_bottom_out_19_;
wire [0:0] sb_2__2__0_chany_bottom_out_1_;
wire [0:0] sb_2__2__0_chany_bottom_out_21_;
wire [0:0] sb_2__2__0_chany_bottom_out_23_;
wire [0:0] sb_2__2__0_chany_bottom_out_25_;
wire [0:0] sb_2__2__0_chany_bottom_out_27_;
wire [0:0] sb_2__2__0_chany_bottom_out_29_;
wire [0:0] sb_2__2__0_chany_bottom_out_31_;
wire [0:0] sb_2__2__0_chany_bottom_out_33_;
wire [0:0] sb_2__2__0_chany_bottom_out_35_;
wire [0:0] sb_2__2__0_chany_bottom_out_37_;
wire [0:0] sb_2__2__0_chany_bottom_out_39_;
wire [0:0] sb_2__2__0_chany_bottom_out_3_;
wire [0:0] sb_2__2__0_chany_bottom_out_41_;
wire [0:0] sb_2__2__0_chany_bottom_out_43_;
wire [0:0] sb_2__2__0_chany_bottom_out_45_;
wire [0:0] sb_2__2__0_chany_bottom_out_47_;
wire [0:0] sb_2__2__0_chany_bottom_out_49_;
wire [0:0] sb_2__2__0_chany_bottom_out_51_;
wire [0:0] sb_2__2__0_chany_bottom_out_53_;
wire [0:0] sb_2__2__0_chany_bottom_out_55_;
wire [0:0] sb_2__2__0_chany_bottom_out_57_;
wire [0:0] sb_2__2__0_chany_bottom_out_59_;
wire [0:0] sb_2__2__0_chany_bottom_out_5_;
wire [0:0] sb_2__2__0_chany_bottom_out_61_;
wire [0:0] sb_2__2__0_chany_bottom_out_63_;
wire [0:0] sb_2__2__0_chany_bottom_out_65_;
wire [0:0] sb_2__2__0_chany_bottom_out_67_;
wire [0:0] sb_2__2__0_chany_bottom_out_69_;
wire [0:0] sb_2__2__0_chany_bottom_out_71_;
wire [0:0] sb_2__2__0_chany_bottom_out_73_;
wire [0:0] sb_2__2__0_chany_bottom_out_75_;
wire [0:0] sb_2__2__0_chany_bottom_out_77_;
wire [0:0] sb_2__2__0_chany_bottom_out_79_;
wire [0:0] sb_2__2__0_chany_bottom_out_7_;
wire [0:0] sb_2__2__0_chany_bottom_out_81_;
wire [0:0] sb_2__2__0_chany_bottom_out_83_;
wire [0:0] sb_2__2__0_chany_bottom_out_85_;
wire [0:0] sb_2__2__0_chany_bottom_out_87_;
wire [0:0] sb_2__2__0_chany_bottom_out_89_;
wire [0:0] sb_2__2__0_chany_bottom_out_91_;
wire [0:0] sb_2__2__0_chany_bottom_out_93_;
wire [0:0] sb_2__2__0_chany_bottom_out_95_;
wire [0:0] sb_2__2__0_chany_bottom_out_97_;
wire [0:0] sb_2__2__0_chany_bottom_out_99_;
wire [0:0] sb_2__2__0_chany_bottom_out_9_;

// ----- BEGIN Local short connections -----

assign lut4_out_0 = gfpga_pad_frac_lut6_spypad_lut4_spy[0]; assign lut4_out_1 = gfpga_pad_frac_lut6_spypad_lut4_spy[1]; assign lut4_out_2 = gfpga_pad_frac_lut6_spypad_lut4_spy[2]; assign lut4_out_3 = gfpga_pad_frac_lut6_spypad_lut4_spy[3]; assign lut5_out_0 = gfpga_pad_frac_lut6_spypad_lut5_spy[0]; assign lut5_out_1 = gfpga_pad_frac_lut6_spypad_lut5_spy[1]; assign lut6_out_0 = gfpga_pad_frac_lut6_spypad_lut6_spy[0]; assign grid_clb_1_2_undriven_top_width_0_height_0__pin_40_[0] = sc_head; assign sc_tail = grid_clb_2_1_undriven_bottom_width_0_height_0__pin_64_[0]; assign cc_spypad_0 = grid_io_bottom_0_ccff_tail[0]; assign cc_spypad_1 = grid_io_left_0_ccff_tail[0]; assign cc_spypad_2 = grid_clb_spypad_0_ccff_tail[0]; assign sc_spypad_0 = grid_clb_1_1_undriven_bottom_width_0_height_0__pin_64_[0]; assign shiftreg_spypad_0 = grid_clb_spypad_0_bottom_width_0_height_0__pin_67_lower[0]; assign cout_spypad_0 = grid_clb_1_1_undriven_bottom_width_0_height_0__pin_65_[0]; assign perf_spypad_0 = grid_clb_1_1_undriven_top_width_0_height_0__pin_68_[0]; assign grid_clb_1_1_undriven_top_width_0_height_0__pin_41_[0] = grid_clb_1_2_undriven_bottom_width_0_height_0__pin_65_[0]; assign grid_clb_1_1_undriven_top_width_0_height_0__pin_40_[0] = grid_clb_1_2_undriven_bottom_width_0_height_0__pin_64_[0]; assign grid_clb_2_2_undriven_top_width_0_height_0__pin_40_[0] = grid_clb_1_1_undriven_bottom_width_0_height_0__pin_64_[0];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	grid_clb_spypad grid_clb_1_1 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.Reset(Reset[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.gfpga_pad_frac_lut6_spypad_lut4_spy(gfpga_pad_frac_lut6_spypad_lut4_spy[0:3]),
		.gfpga_pad_frac_lut6_spypad_lut5_spy(gfpga_pad_frac_lut6_spypad_lut5_spy[0:1]),
		.gfpga_pad_frac_lut6_spypad_lut6_spy(gfpga_pad_frac_lut6_spypad_lut6_spy[0]),
		.top_width_0_height_0__pin_40_(grid_clb_1_1_undriven_top_width_0_height_0__pin_40_[0]),
		.top_width_0_height_0__pin_41_(grid_clb_1_1_undriven_top_width_0_height_0__pin_41_[0]),
		.top_width_0_height_0__pin_42_(cbx_1__1__0_bottom_grid_pin_42_[0]),
		.top_width_0_height_0__pin_43_(cbx_1__1__0_bottom_grid_pin_43_[0]),
		.top_width_0_height_0__pin_69_(cbx_1__1__0_bottom_grid_pin_69_[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__0_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__0_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__0_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__0_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__0_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__0_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__0_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__0_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__0_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__0_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__0_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__0_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__0_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__0_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__0_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__0_left_grid_pin_15_[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__0_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__0_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__0_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__0_left_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__0__0_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__0__0_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__0__0_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__0__0_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__0__0_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__0__0_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__0__0_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__0__0_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__0__0_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__0__0_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__0__0_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__0__0_top_grid_pin_31_[0]),
		.bottom_width_0_height_0__pin_32_(cbx_1__0__0_top_grid_pin_32_[0]),
		.bottom_width_0_height_0__pin_33_(cbx_1__0__0_top_grid_pin_33_[0]),
		.bottom_width_0_height_0__pin_34_(cbx_1__0__0_top_grid_pin_34_[0]),
		.bottom_width_0_height_0__pin_35_(cbx_1__0__0_top_grid_pin_35_[0]),
		.bottom_width_0_height_0__pin_36_(cbx_1__0__0_top_grid_pin_36_[0]),
		.bottom_width_0_height_0__pin_37_(cbx_1__0__0_top_grid_pin_37_[0]),
		.bottom_width_0_height_0__pin_38_(cbx_1__0__0_top_grid_pin_38_[0]),
		.bottom_width_0_height_0__pin_39_(cbx_1__0__0_top_grid_pin_39_[0]),
		.ccff_head(cby_1__1__0_ccff_tail[0]),
		.top_width_0_height_0__pin_68_(grid_clb_1_1_undriven_top_width_0_height_0__pin_68_[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_spypad_0_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_spypad_0_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_spypad_0_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_spypad_0_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_spypad_0_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_spypad_0_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_spypad_0_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_spypad_0_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_spypad_0_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_spypad_0_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_spypad_0_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_spypad_0_right_width_0_height_0__pin_49_lower[0]),
		.right_width_0_height_0__pin_50_upper(grid_clb_spypad_0_right_width_0_height_0__pin_50_upper[0]),
		.right_width_0_height_0__pin_50_lower(grid_clb_spypad_0_right_width_0_height_0__pin_50_lower[0]),
		.right_width_0_height_0__pin_51_upper(grid_clb_spypad_0_right_width_0_height_0__pin_51_upper[0]),
		.right_width_0_height_0__pin_51_lower(grid_clb_spypad_0_right_width_0_height_0__pin_51_lower[0]),
		.right_width_0_height_0__pin_52_upper(grid_clb_spypad_0_right_width_0_height_0__pin_52_upper[0]),
		.right_width_0_height_0__pin_52_lower(grid_clb_spypad_0_right_width_0_height_0__pin_52_lower[0]),
		.right_width_0_height_0__pin_53_upper(grid_clb_spypad_0_right_width_0_height_0__pin_53_upper[0]),
		.right_width_0_height_0__pin_53_lower(grid_clb_spypad_0_right_width_0_height_0__pin_53_lower[0]),
		.bottom_width_0_height_0__pin_54_upper(grid_clb_spypad_0_bottom_width_0_height_0__pin_54_upper[0]),
		.bottom_width_0_height_0__pin_54_lower(grid_clb_spypad_0_bottom_width_0_height_0__pin_54_lower[0]),
		.bottom_width_0_height_0__pin_55_upper(grid_clb_spypad_0_bottom_width_0_height_0__pin_55_upper[0]),
		.bottom_width_0_height_0__pin_55_lower(grid_clb_spypad_0_bottom_width_0_height_0__pin_55_lower[0]),
		.bottom_width_0_height_0__pin_56_upper(grid_clb_spypad_0_bottom_width_0_height_0__pin_56_upper[0]),
		.bottom_width_0_height_0__pin_56_lower(grid_clb_spypad_0_bottom_width_0_height_0__pin_56_lower[0]),
		.bottom_width_0_height_0__pin_57_upper(grid_clb_spypad_0_bottom_width_0_height_0__pin_57_upper[0]),
		.bottom_width_0_height_0__pin_57_lower(grid_clb_spypad_0_bottom_width_0_height_0__pin_57_lower[0]),
		.bottom_width_0_height_0__pin_58_upper(grid_clb_spypad_0_bottom_width_0_height_0__pin_58_upper[0]),
		.bottom_width_0_height_0__pin_58_lower(grid_clb_spypad_0_bottom_width_0_height_0__pin_58_lower[0]),
		.bottom_width_0_height_0__pin_59_upper(grid_clb_spypad_0_bottom_width_0_height_0__pin_59_upper[0]),
		.bottom_width_0_height_0__pin_59_lower(grid_clb_spypad_0_bottom_width_0_height_0__pin_59_lower[0]),
		.bottom_width_0_height_0__pin_60_upper(grid_clb_spypad_0_bottom_width_0_height_0__pin_60_upper[0]),
		.bottom_width_0_height_0__pin_60_lower(grid_clb_spypad_0_bottom_width_0_height_0__pin_60_lower[0]),
		.bottom_width_0_height_0__pin_61_upper(grid_clb_spypad_0_bottom_width_0_height_0__pin_61_upper[0]),
		.bottom_width_0_height_0__pin_61_lower(grid_clb_spypad_0_bottom_width_0_height_0__pin_61_lower[0]),
		.bottom_width_0_height_0__pin_62_upper(grid_clb_spypad_0_bottom_width_0_height_0__pin_62_upper[0]),
		.bottom_width_0_height_0__pin_62_lower(grid_clb_spypad_0_bottom_width_0_height_0__pin_62_lower[0]),
		.bottom_width_0_height_0__pin_63_upper(grid_clb_spypad_0_bottom_width_0_height_0__pin_63_upper[0]),
		.bottom_width_0_height_0__pin_63_lower(grid_clb_spypad_0_bottom_width_0_height_0__pin_63_lower[0]),
		.bottom_width_0_height_0__pin_64_(grid_clb_1_1_undriven_bottom_width_0_height_0__pin_64_[0]),
		.bottom_width_0_height_0__pin_65_(grid_clb_1_1_undriven_bottom_width_0_height_0__pin_65_[0]),
		.bottom_width_0_height_0__pin_66_upper(grid_clb_spypad_0_bottom_width_0_height_0__pin_66_upper[0]),
		.bottom_width_0_height_0__pin_66_lower(grid_clb_spypad_0_bottom_width_0_height_0__pin_66_lower[0]),
		.bottom_width_0_height_0__pin_67_upper(grid_clb_spypad_0_bottom_width_0_height_0__pin_67_upper[0]),
		.bottom_width_0_height_0__pin_67_lower(grid_clb_spypad_0_bottom_width_0_height_0__pin_67_lower[0]),
		.ccff_tail(grid_clb_spypad_0_ccff_tail[0]));

	grid_clb grid_clb_1_2 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.Reset(Reset[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_40_(grid_clb_1_2_undriven_top_width_0_height_0__pin_40_[0]),
		.top_width_0_height_0__pin_41_(grid_clb_1_2_undriven_top_width_0_height_0__pin_41_[0]),
		.top_width_0_height_0__pin_42_(cbx_1__2__0_bottom_grid_pin_42_[0]),
		.top_width_0_height_0__pin_43_(cbx_1__2__0_bottom_grid_pin_43_[0]),
		.top_width_0_height_0__pin_68_(cbx_1__2__0_bottom_grid_pin_68_[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__1_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__1_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__1_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__1_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__1_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__1_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__1_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__1_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__1_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__1_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__1_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__1_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__1_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__1_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__1_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__1_left_grid_pin_15_[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__1_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__1_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__1_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__1_left_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__0_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__0_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__0_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__0_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__0_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__0_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__0_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__0_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__0_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__0_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__0_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__0_top_grid_pin_31_[0]),
		.bottom_width_0_height_0__pin_32_(cbx_1__1__0_top_grid_pin_32_[0]),
		.bottom_width_0_height_0__pin_33_(cbx_1__1__0_top_grid_pin_33_[0]),
		.bottom_width_0_height_0__pin_34_(cbx_1__1__0_top_grid_pin_34_[0]),
		.bottom_width_0_height_0__pin_35_(cbx_1__1__0_top_grid_pin_35_[0]),
		.bottom_width_0_height_0__pin_36_(cbx_1__1__0_top_grid_pin_36_[0]),
		.bottom_width_0_height_0__pin_37_(cbx_1__1__0_top_grid_pin_37_[0]),
		.bottom_width_0_height_0__pin_38_(cbx_1__1__0_top_grid_pin_38_[0]),
		.bottom_width_0_height_0__pin_39_(cbx_1__1__0_top_grid_pin_39_[0]),
		.ccff_head(cby_1__1__1_ccff_tail[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_0_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_0_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_0_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_0_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_0_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_0_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_0_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_0_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_0_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_0_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_0_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_0_right_width_0_height_0__pin_49_lower[0]),
		.right_width_0_height_0__pin_50_upper(grid_clb_0_right_width_0_height_0__pin_50_upper[0]),
		.right_width_0_height_0__pin_50_lower(grid_clb_0_right_width_0_height_0__pin_50_lower[0]),
		.right_width_0_height_0__pin_51_upper(grid_clb_0_right_width_0_height_0__pin_51_upper[0]),
		.right_width_0_height_0__pin_51_lower(grid_clb_0_right_width_0_height_0__pin_51_lower[0]),
		.right_width_0_height_0__pin_52_upper(grid_clb_0_right_width_0_height_0__pin_52_upper[0]),
		.right_width_0_height_0__pin_52_lower(grid_clb_0_right_width_0_height_0__pin_52_lower[0]),
		.right_width_0_height_0__pin_53_upper(grid_clb_0_right_width_0_height_0__pin_53_upper[0]),
		.right_width_0_height_0__pin_53_lower(grid_clb_0_right_width_0_height_0__pin_53_lower[0]),
		.bottom_width_0_height_0__pin_54_upper(grid_clb_0_bottom_width_0_height_0__pin_54_upper[0]),
		.bottom_width_0_height_0__pin_54_lower(grid_clb_0_bottom_width_0_height_0__pin_54_lower[0]),
		.bottom_width_0_height_0__pin_55_upper(grid_clb_0_bottom_width_0_height_0__pin_55_upper[0]),
		.bottom_width_0_height_0__pin_55_lower(grid_clb_0_bottom_width_0_height_0__pin_55_lower[0]),
		.bottom_width_0_height_0__pin_56_upper(grid_clb_0_bottom_width_0_height_0__pin_56_upper[0]),
		.bottom_width_0_height_0__pin_56_lower(grid_clb_0_bottom_width_0_height_0__pin_56_lower[0]),
		.bottom_width_0_height_0__pin_57_upper(grid_clb_0_bottom_width_0_height_0__pin_57_upper[0]),
		.bottom_width_0_height_0__pin_57_lower(grid_clb_0_bottom_width_0_height_0__pin_57_lower[0]),
		.bottom_width_0_height_0__pin_58_upper(grid_clb_0_bottom_width_0_height_0__pin_58_upper[0]),
		.bottom_width_0_height_0__pin_58_lower(grid_clb_0_bottom_width_0_height_0__pin_58_lower[0]),
		.bottom_width_0_height_0__pin_59_upper(grid_clb_0_bottom_width_0_height_0__pin_59_upper[0]),
		.bottom_width_0_height_0__pin_59_lower(grid_clb_0_bottom_width_0_height_0__pin_59_lower[0]),
		.bottom_width_0_height_0__pin_60_upper(grid_clb_0_bottom_width_0_height_0__pin_60_upper[0]),
		.bottom_width_0_height_0__pin_60_lower(grid_clb_0_bottom_width_0_height_0__pin_60_lower[0]),
		.bottom_width_0_height_0__pin_61_upper(grid_clb_0_bottom_width_0_height_0__pin_61_upper[0]),
		.bottom_width_0_height_0__pin_61_lower(grid_clb_0_bottom_width_0_height_0__pin_61_lower[0]),
		.bottom_width_0_height_0__pin_62_upper(grid_clb_0_bottom_width_0_height_0__pin_62_upper[0]),
		.bottom_width_0_height_0__pin_62_lower(grid_clb_0_bottom_width_0_height_0__pin_62_lower[0]),
		.bottom_width_0_height_0__pin_63_upper(grid_clb_0_bottom_width_0_height_0__pin_63_upper[0]),
		.bottom_width_0_height_0__pin_63_lower(grid_clb_0_bottom_width_0_height_0__pin_63_lower[0]),
		.bottom_width_0_height_0__pin_64_(grid_clb_1_2_undriven_bottom_width_0_height_0__pin_64_[0]),
		.bottom_width_0_height_0__pin_65_(grid_clb_1_2_undriven_bottom_width_0_height_0__pin_65_[0]),
		.bottom_width_0_height_0__pin_66_upper(grid_clb_0_bottom_width_0_height_0__pin_66_upper[0]),
		.bottom_width_0_height_0__pin_66_lower(grid_clb_0_bottom_width_0_height_0__pin_66_lower[0]),
		.bottom_width_0_height_0__pin_67_upper(grid_clb_0_bottom_width_0_height_0__pin_67_upper[0]),
		.bottom_width_0_height_0__pin_67_lower(grid_clb_0_bottom_width_0_height_0__pin_67_lower[0]),
		.ccff_tail(ccff_tail[0]));

	grid_clb grid_clb_2_1 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.Reset(Reset[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_40_(direct_interc_1_out[0]),
		.top_width_0_height_0__pin_41_(direct_interc_0_out[0]),
		.top_width_0_height_0__pin_42_(cbx_1__1__1_bottom_grid_pin_42_[0]),
		.top_width_0_height_0__pin_43_(cbx_1__1__1_bottom_grid_pin_43_[0]),
		.top_width_0_height_0__pin_68_(cbx_1__1__1_bottom_grid_pin_69_[0]),
		.right_width_0_height_0__pin_0_(cby_2__1__0_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_2__1__0_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_2__1__0_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_2__1__0_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_2__1__0_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_2__1__0_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_2__1__0_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_2__1__0_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_2__1__0_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_2__1__0_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_2__1__0_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_2__1__0_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_2__1__0_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_2__1__0_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_2__1__0_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_2__1__0_left_grid_pin_15_[0]),
		.right_width_0_height_0__pin_16_(cby_2__1__0_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_2__1__0_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_2__1__0_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_2__1__0_left_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__0__1_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__0__1_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__0__1_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__0__1_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__0__1_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__0__1_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__0__1_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__0__1_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__0__1_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__0__1_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__0__1_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__0__1_top_grid_pin_31_[0]),
		.bottom_width_0_height_0__pin_32_(cbx_1__0__1_top_grid_pin_32_[0]),
		.bottom_width_0_height_0__pin_33_(cbx_1__0__1_top_grid_pin_33_[0]),
		.bottom_width_0_height_0__pin_34_(cbx_1__0__1_top_grid_pin_34_[0]),
		.bottom_width_0_height_0__pin_35_(cbx_1__0__1_top_grid_pin_35_[0]),
		.bottom_width_0_height_0__pin_36_(cbx_1__0__1_top_grid_pin_36_[0]),
		.bottom_width_0_height_0__pin_37_(cbx_1__0__1_top_grid_pin_37_[0]),
		.bottom_width_0_height_0__pin_38_(cbx_1__0__1_top_grid_pin_38_[0]),
		.bottom_width_0_height_0__pin_39_(cbx_1__0__1_top_grid_pin_39_[0]),
		.ccff_head(cby_2__1__0_ccff_tail[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_1_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_1_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_1_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_1_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_1_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_1_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_1_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_1_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_1_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_1_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_1_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_1_right_width_0_height_0__pin_49_lower[0]),
		.right_width_0_height_0__pin_50_upper(grid_clb_1_right_width_0_height_0__pin_50_upper[0]),
		.right_width_0_height_0__pin_50_lower(grid_clb_1_right_width_0_height_0__pin_50_lower[0]),
		.right_width_0_height_0__pin_51_upper(grid_clb_1_right_width_0_height_0__pin_51_upper[0]),
		.right_width_0_height_0__pin_51_lower(grid_clb_1_right_width_0_height_0__pin_51_lower[0]),
		.right_width_0_height_0__pin_52_upper(grid_clb_1_right_width_0_height_0__pin_52_upper[0]),
		.right_width_0_height_0__pin_52_lower(grid_clb_1_right_width_0_height_0__pin_52_lower[0]),
		.right_width_0_height_0__pin_53_upper(grid_clb_1_right_width_0_height_0__pin_53_upper[0]),
		.right_width_0_height_0__pin_53_lower(grid_clb_1_right_width_0_height_0__pin_53_lower[0]),
		.bottom_width_0_height_0__pin_54_upper(grid_clb_1_bottom_width_0_height_0__pin_54_upper[0]),
		.bottom_width_0_height_0__pin_54_lower(grid_clb_1_bottom_width_0_height_0__pin_54_lower[0]),
		.bottom_width_0_height_0__pin_55_upper(grid_clb_1_bottom_width_0_height_0__pin_55_upper[0]),
		.bottom_width_0_height_0__pin_55_lower(grid_clb_1_bottom_width_0_height_0__pin_55_lower[0]),
		.bottom_width_0_height_0__pin_56_upper(grid_clb_1_bottom_width_0_height_0__pin_56_upper[0]),
		.bottom_width_0_height_0__pin_56_lower(grid_clb_1_bottom_width_0_height_0__pin_56_lower[0]),
		.bottom_width_0_height_0__pin_57_upper(grid_clb_1_bottom_width_0_height_0__pin_57_upper[0]),
		.bottom_width_0_height_0__pin_57_lower(grid_clb_1_bottom_width_0_height_0__pin_57_lower[0]),
		.bottom_width_0_height_0__pin_58_upper(grid_clb_1_bottom_width_0_height_0__pin_58_upper[0]),
		.bottom_width_0_height_0__pin_58_lower(grid_clb_1_bottom_width_0_height_0__pin_58_lower[0]),
		.bottom_width_0_height_0__pin_59_upper(grid_clb_1_bottom_width_0_height_0__pin_59_upper[0]),
		.bottom_width_0_height_0__pin_59_lower(grid_clb_1_bottom_width_0_height_0__pin_59_lower[0]),
		.bottom_width_0_height_0__pin_60_upper(grid_clb_1_bottom_width_0_height_0__pin_60_upper[0]),
		.bottom_width_0_height_0__pin_60_lower(grid_clb_1_bottom_width_0_height_0__pin_60_lower[0]),
		.bottom_width_0_height_0__pin_61_upper(grid_clb_1_bottom_width_0_height_0__pin_61_upper[0]),
		.bottom_width_0_height_0__pin_61_lower(grid_clb_1_bottom_width_0_height_0__pin_61_lower[0]),
		.bottom_width_0_height_0__pin_62_upper(grid_clb_1_bottom_width_0_height_0__pin_62_upper[0]),
		.bottom_width_0_height_0__pin_62_lower(grid_clb_1_bottom_width_0_height_0__pin_62_lower[0]),
		.bottom_width_0_height_0__pin_63_upper(grid_clb_1_bottom_width_0_height_0__pin_63_upper[0]),
		.bottom_width_0_height_0__pin_63_lower(grid_clb_1_bottom_width_0_height_0__pin_63_lower[0]),
		.bottom_width_0_height_0__pin_64_(grid_clb_2_1_undriven_bottom_width_0_height_0__pin_64_[0]),
		.bottom_width_0_height_0__pin_65_(grid_clb_2_1_undriven_bottom_width_0_height_0__pin_65_[0]),
		.bottom_width_0_height_0__pin_66_upper(grid_clb_1_bottom_width_0_height_0__pin_66_upper[0]),
		.bottom_width_0_height_0__pin_66_lower(grid_clb_1_bottom_width_0_height_0__pin_66_lower[0]),
		.bottom_width_0_height_0__pin_67_upper(grid_clb_1_bottom_width_0_height_0__pin_67_upper[0]),
		.bottom_width_0_height_0__pin_67_lower(grid_clb_1_bottom_width_0_height_0__pin_67_lower[0]),
		.ccff_tail(grid_clb_1_ccff_tail[0]));

	grid_clb grid_clb_2_2 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.Reset(Reset[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_40_(grid_clb_2_2_undriven_top_width_0_height_0__pin_40_[0]),
		.top_width_0_height_0__pin_41_(grid_clb_2_2_undriven_top_width_0_height_0__pin_41_[0]),
		.top_width_0_height_0__pin_42_(cbx_1__2__1_bottom_grid_pin_42_[0]),
		.top_width_0_height_0__pin_43_(cbx_1__2__1_bottom_grid_pin_43_[0]),
		.top_width_0_height_0__pin_68_(cbx_1__2__1_bottom_grid_pin_68_[0]),
		.right_width_0_height_0__pin_0_(cby_2__1__1_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_2__1__1_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_2__1__1_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_2__1__1_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_2__1__1_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_2__1__1_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_2__1__1_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_2__1__1_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_2__1__1_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_2__1__1_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_2__1__1_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_2__1__1_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_2__1__1_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_2__1__1_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_2__1__1_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_2__1__1_left_grid_pin_15_[0]),
		.right_width_0_height_0__pin_16_(cby_2__1__1_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_2__1__1_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_2__1__1_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_2__1__1_left_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__1_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__1_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__1_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__1_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__1_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__1_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__1_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__1_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__1_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__1_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__1_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__1_top_grid_pin_31_[0]),
		.bottom_width_0_height_0__pin_32_(cbx_1__1__1_top_grid_pin_32_[0]),
		.bottom_width_0_height_0__pin_33_(cbx_1__1__1_top_grid_pin_33_[0]),
		.bottom_width_0_height_0__pin_34_(cbx_1__1__1_top_grid_pin_34_[0]),
		.bottom_width_0_height_0__pin_35_(cbx_1__1__1_top_grid_pin_35_[0]),
		.bottom_width_0_height_0__pin_36_(cbx_1__1__1_top_grid_pin_36_[0]),
		.bottom_width_0_height_0__pin_37_(cbx_1__1__1_top_grid_pin_37_[0]),
		.bottom_width_0_height_0__pin_38_(cbx_1__1__1_top_grid_pin_38_[0]),
		.bottom_width_0_height_0__pin_39_(cbx_1__1__1_top_grid_pin_39_[0]),
		.ccff_head(cby_2__1__1_ccff_tail[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_2_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_2_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_2_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_2_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_2_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_2_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_2_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_2_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_2_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_2_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_2_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_2_right_width_0_height_0__pin_49_lower[0]),
		.right_width_0_height_0__pin_50_upper(grid_clb_2_right_width_0_height_0__pin_50_upper[0]),
		.right_width_0_height_0__pin_50_lower(grid_clb_2_right_width_0_height_0__pin_50_lower[0]),
		.right_width_0_height_0__pin_51_upper(grid_clb_2_right_width_0_height_0__pin_51_upper[0]),
		.right_width_0_height_0__pin_51_lower(grid_clb_2_right_width_0_height_0__pin_51_lower[0]),
		.right_width_0_height_0__pin_52_upper(grid_clb_2_right_width_0_height_0__pin_52_upper[0]),
		.right_width_0_height_0__pin_52_lower(grid_clb_2_right_width_0_height_0__pin_52_lower[0]),
		.right_width_0_height_0__pin_53_upper(grid_clb_2_right_width_0_height_0__pin_53_upper[0]),
		.right_width_0_height_0__pin_53_lower(grid_clb_2_right_width_0_height_0__pin_53_lower[0]),
		.bottom_width_0_height_0__pin_54_upper(grid_clb_2_bottom_width_0_height_0__pin_54_upper[0]),
		.bottom_width_0_height_0__pin_54_lower(grid_clb_2_bottom_width_0_height_0__pin_54_lower[0]),
		.bottom_width_0_height_0__pin_55_upper(grid_clb_2_bottom_width_0_height_0__pin_55_upper[0]),
		.bottom_width_0_height_0__pin_55_lower(grid_clb_2_bottom_width_0_height_0__pin_55_lower[0]),
		.bottom_width_0_height_0__pin_56_upper(grid_clb_2_bottom_width_0_height_0__pin_56_upper[0]),
		.bottom_width_0_height_0__pin_56_lower(grid_clb_2_bottom_width_0_height_0__pin_56_lower[0]),
		.bottom_width_0_height_0__pin_57_upper(grid_clb_2_bottom_width_0_height_0__pin_57_upper[0]),
		.bottom_width_0_height_0__pin_57_lower(grid_clb_2_bottom_width_0_height_0__pin_57_lower[0]),
		.bottom_width_0_height_0__pin_58_upper(grid_clb_2_bottom_width_0_height_0__pin_58_upper[0]),
		.bottom_width_0_height_0__pin_58_lower(grid_clb_2_bottom_width_0_height_0__pin_58_lower[0]),
		.bottom_width_0_height_0__pin_59_upper(grid_clb_2_bottom_width_0_height_0__pin_59_upper[0]),
		.bottom_width_0_height_0__pin_59_lower(grid_clb_2_bottom_width_0_height_0__pin_59_lower[0]),
		.bottom_width_0_height_0__pin_60_upper(grid_clb_2_bottom_width_0_height_0__pin_60_upper[0]),
		.bottom_width_0_height_0__pin_60_lower(grid_clb_2_bottom_width_0_height_0__pin_60_lower[0]),
		.bottom_width_0_height_0__pin_61_upper(grid_clb_2_bottom_width_0_height_0__pin_61_upper[0]),
		.bottom_width_0_height_0__pin_61_lower(grid_clb_2_bottom_width_0_height_0__pin_61_lower[0]),
		.bottom_width_0_height_0__pin_62_upper(grid_clb_2_bottom_width_0_height_0__pin_62_upper[0]),
		.bottom_width_0_height_0__pin_62_lower(grid_clb_2_bottom_width_0_height_0__pin_62_lower[0]),
		.bottom_width_0_height_0__pin_63_upper(grid_clb_2_bottom_width_0_height_0__pin_63_upper[0]),
		.bottom_width_0_height_0__pin_63_lower(grid_clb_2_bottom_width_0_height_0__pin_63_lower[0]),
		.bottom_width_0_height_0__pin_64_(grid_clb_2_bottom_width_0_height_0__pin_64_[0]),
		.bottom_width_0_height_0__pin_65_(grid_clb_2_bottom_width_0_height_0__pin_65_[0]),
		.bottom_width_0_height_0__pin_66_upper(grid_clb_2_bottom_width_0_height_0__pin_66_upper[0]),
		.bottom_width_0_height_0__pin_66_lower(grid_clb_2_bottom_width_0_height_0__pin_66_lower[0]),
		.bottom_width_0_height_0__pin_67_upper(grid_clb_2_bottom_width_0_height_0__pin_67_upper[0]),
		.bottom_width_0_height_0__pin_67_lower(grid_clb_2_bottom_width_0_height_0__pin_67_lower[0]),
		.ccff_tail(grid_clb_2_ccff_tail[0]));

	grid_io_top grid_io_top_1_3 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[0]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[0]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[0]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[0]),
		.bottom_width_0_height_0__pin_0_(cbx_1__2__0_top_grid_pin_0_[0]),
		.ccff_head(cbx_1__2__0_ccff_tail[0]),
		.bottom_width_0_height_0__pin_1_upper(grid_io_top_0_bottom_width_0_height_0__pin_1_upper[0]),
		.bottom_width_0_height_0__pin_1_lower(grid_io_top_0_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_top_0_ccff_tail[0]));

	grid_io_top grid_io_top_2_3 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[1]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[1]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[1]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[1]),
		.bottom_width_0_height_0__pin_0_(cbx_1__2__1_top_grid_pin_0_[0]),
		.ccff_head(cbx_1__2__1_ccff_tail[0]),
		.bottom_width_0_height_0__pin_1_upper(grid_io_top_1_bottom_width_0_height_0__pin_1_upper[0]),
		.bottom_width_0_height_0__pin_1_lower(grid_io_top_1_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_top_1_ccff_tail[0]));

	grid_io_right grid_io_right_3_1 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[2]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[2]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[2]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[2]),
		.left_width_0_height_0__pin_0_(cby_2__1__0_right_grid_pin_0_[0]),
		.ccff_head(grid_io_bottom_1_ccff_tail[0]),
		.left_width_0_height_0__pin_1_upper(grid_io_right_0_left_width_0_height_0__pin_1_upper[0]),
		.left_width_0_height_0__pin_1_lower(grid_io_right_0_left_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_right_0_ccff_tail[0]));

	grid_io_right grid_io_right_3_2 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[3]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[3]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[3]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[3]),
		.left_width_0_height_0__pin_0_(cby_2__1__1_right_grid_pin_0_[0]),
		.ccff_head(grid_io_right_0_ccff_tail[0]),
		.left_width_0_height_0__pin_1_upper(grid_io_right_1_left_width_0_height_0__pin_1_upper[0]),
		.left_width_0_height_0__pin_1_lower(grid_io_right_1_left_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_right_1_ccff_tail[0]));

	grid_io_bottom grid_io_bottom_1_0 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[4]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[4]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[4]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[4]),
		.top_width_0_height_0__pin_0_(cbx_1__0__0_bottom_grid_pin_0_[0]),
		.ccff_head(ccff_head[0]),
		.top_width_0_height_0__pin_1_upper(grid_io_bottom_0_top_width_0_height_0__pin_1_upper[0]),
		.top_width_0_height_0__pin_1_lower(grid_io_bottom_0_top_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_bottom_0_ccff_tail[0]));

	grid_io_bottom grid_io_bottom_2_0 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[5]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[5]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[5]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[5]),
		.top_width_0_height_0__pin_0_(cbx_1__0__1_bottom_grid_pin_0_[0]),
		.ccff_head(grid_io_bottom_0_ccff_tail[0]),
		.top_width_0_height_0__pin_1_upper(grid_io_bottom_1_top_width_0_height_0__pin_1_upper[0]),
		.top_width_0_height_0__pin_1_lower(grid_io_bottom_1_top_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_bottom_1_ccff_tail[0]));

	grid_io_left grid_io_left_0_1 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[6]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[6]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[6]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[6]),
		.right_width_0_height_0__pin_0_(cby_0__1__0_left_grid_pin_0_[0]),
		.ccff_head(cby_0__1__0_ccff_tail[0]),
		.right_width_0_height_0__pin_1_upper(grid_io_left_0_right_width_0_height_0__pin_1_upper[0]),
		.right_width_0_height_0__pin_1_lower(grid_io_left_0_right_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_left_0_ccff_tail[0]));

	grid_io_left grid_io_left_0_2 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[7]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[7]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[7]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[7]),
		.right_width_0_height_0__pin_0_(cby_0__1__1_left_grid_pin_0_[0]),
		.ccff_head(cby_0__1__1_ccff_tail[0]),
		.right_width_0_height_0__pin_1_upper(grid_io_left_1_right_width_0_height_0__pin_1_upper[0]),
		.right_width_0_height_0__pin_1_lower(grid_io_left_1_right_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_left_1_ccff_tail[0]));

	sb_0__0_ sb_0__0_ (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.chany_top_in_1_(cby_0__1__0_chany_out_1_[0]),
		.chany_top_in_3_(cby_0__1__0_chany_out_3_[0]),
		.chany_top_in_5_(cby_0__1__0_chany_out_5_[0]),
		.chany_top_in_7_(cby_0__1__0_chany_out_7_[0]),
		.chany_top_in_9_(cby_0__1__0_chany_out_9_[0]),
		.chany_top_in_11_(cby_0__1__0_chany_out_11_[0]),
		.chany_top_in_13_(cby_0__1__0_chany_out_13_[0]),
		.chany_top_in_15_(cby_0__1__0_chany_out_15_[0]),
		.chany_top_in_17_(cby_0__1__0_chany_out_17_[0]),
		.chany_top_in_19_(cby_0__1__0_chany_out_19_[0]),
		.chany_top_in_21_(cby_0__1__0_chany_out_21_[0]),
		.chany_top_in_23_(cby_0__1__0_chany_out_23_[0]),
		.chany_top_in_25_(cby_0__1__0_chany_out_25_[0]),
		.chany_top_in_27_(cby_0__1__0_chany_out_27_[0]),
		.chany_top_in_29_(cby_0__1__0_chany_out_29_[0]),
		.chany_top_in_31_(cby_0__1__0_chany_out_31_[0]),
		.chany_top_in_33_(cby_0__1__0_chany_out_33_[0]),
		.chany_top_in_35_(cby_0__1__0_chany_out_35_[0]),
		.chany_top_in_37_(cby_0__1__0_chany_out_37_[0]),
		.chany_top_in_39_(cby_0__1__0_chany_out_39_[0]),
		.chany_top_in_41_(cby_0__1__0_chany_out_41_[0]),
		.chany_top_in_43_(cby_0__1__0_chany_out_43_[0]),
		.chany_top_in_45_(cby_0__1__0_chany_out_45_[0]),
		.chany_top_in_47_(cby_0__1__0_chany_out_47_[0]),
		.chany_top_in_49_(cby_0__1__0_chany_out_49_[0]),
		.chany_top_in_51_(cby_0__1__0_chany_out_51_[0]),
		.chany_top_in_53_(cby_0__1__0_chany_out_53_[0]),
		.chany_top_in_55_(cby_0__1__0_chany_out_55_[0]),
		.chany_top_in_57_(cby_0__1__0_chany_out_57_[0]),
		.chany_top_in_59_(cby_0__1__0_chany_out_59_[0]),
		.chany_top_in_61_(cby_0__1__0_chany_out_61_[0]),
		.chany_top_in_63_(cby_0__1__0_chany_out_63_[0]),
		.chany_top_in_65_(cby_0__1__0_chany_out_65_[0]),
		.chany_top_in_67_(cby_0__1__0_chany_out_67_[0]),
		.chany_top_in_69_(cby_0__1__0_chany_out_69_[0]),
		.chany_top_in_71_(cby_0__1__0_chany_out_71_[0]),
		.chany_top_in_73_(cby_0__1__0_chany_out_73_[0]),
		.chany_top_in_75_(cby_0__1__0_chany_out_75_[0]),
		.chany_top_in_77_(cby_0__1__0_chany_out_77_[0]),
		.chany_top_in_79_(cby_0__1__0_chany_out_79_[0]),
		.chany_top_in_81_(cby_0__1__0_chany_out_81_[0]),
		.chany_top_in_83_(cby_0__1__0_chany_out_83_[0]),
		.chany_top_in_85_(cby_0__1__0_chany_out_85_[0]),
		.chany_top_in_87_(cby_0__1__0_chany_out_87_[0]),
		.chany_top_in_89_(cby_0__1__0_chany_out_89_[0]),
		.chany_top_in_91_(cby_0__1__0_chany_out_91_[0]),
		.chany_top_in_93_(cby_0__1__0_chany_out_93_[0]),
		.chany_top_in_95_(cby_0__1__0_chany_out_95_[0]),
		.chany_top_in_97_(cby_0__1__0_chany_out_97_[0]),
		.chany_top_in_99_(cby_0__1__0_chany_out_99_[0]),
		.chany_top_in_101_(cby_0__1__0_chany_out_101_[0]),
		.chany_top_in_103_(cby_0__1__0_chany_out_103_[0]),
		.chany_top_in_105_(cby_0__1__0_chany_out_105_[0]),
		.chany_top_in_107_(cby_0__1__0_chany_out_107_[0]),
		.chany_top_in_109_(cby_0__1__0_chany_out_109_[0]),
		.chany_top_in_111_(cby_0__1__0_chany_out_111_[0]),
		.chany_top_in_113_(cby_0__1__0_chany_out_113_[0]),
		.chany_top_in_115_(cby_0__1__0_chany_out_115_[0]),
		.chany_top_in_117_(cby_0__1__0_chany_out_117_[0]),
		.chany_top_in_119_(cby_0__1__0_chany_out_119_[0]),
		.chany_top_in_121_(cby_0__1__0_chany_out_121_[0]),
		.chany_top_in_123_(cby_0__1__0_chany_out_123_[0]),
		.chany_top_in_125_(cby_0__1__0_chany_out_125_[0]),
		.chany_top_in_127_(cby_0__1__0_chany_out_127_[0]),
		.chany_top_in_129_(cby_0__1__0_chany_out_129_[0]),
		.chany_top_in_131_(cby_0__1__0_chany_out_131_[0]),
		.chany_top_in_133_(cby_0__1__0_chany_out_133_[0]),
		.chany_top_in_135_(cby_0__1__0_chany_out_135_[0]),
		.chany_top_in_137_(cby_0__1__0_chany_out_137_[0]),
		.chany_top_in_139_(cby_0__1__0_chany_out_139_[0]),
		.chany_top_in_141_(cby_0__1__0_chany_out_141_[0]),
		.chany_top_in_143_(cby_0__1__0_chany_out_143_[0]),
		.chany_top_in_145_(cby_0__1__0_chany_out_145_[0]),
		.chany_top_in_147_(cby_0__1__0_chany_out_147_[0]),
		.chany_top_in_149_(cby_0__1__0_chany_out_149_[0]),
		.chany_top_in_151_(cby_0__1__0_chany_out_151_[0]),
		.chany_top_in_153_(cby_0__1__0_chany_out_153_[0]),
		.chany_top_in_155_(cby_0__1__0_chany_out_155_[0]),
		.chany_top_in_157_(cby_0__1__0_chany_out_157_[0]),
		.chany_top_in_159_(cby_0__1__0_chany_out_159_[0]),
		.chany_top_in_161_(cby_0__1__0_chany_out_161_[0]),
		.chany_top_in_163_(cby_0__1__0_chany_out_163_[0]),
		.chany_top_in_165_(cby_0__1__0_chany_out_165_[0]),
		.chany_top_in_167_(cby_0__1__0_chany_out_167_[0]),
		.chany_top_in_169_(cby_0__1__0_chany_out_169_[0]),
		.chany_top_in_171_(cby_0__1__0_chany_out_171_[0]),
		.chany_top_in_173_(cby_0__1__0_chany_out_173_[0]),
		.chany_top_in_175_(cby_0__1__0_chany_out_175_[0]),
		.chany_top_in_177_(cby_0__1__0_chany_out_177_[0]),
		.chany_top_in_179_(cby_0__1__0_chany_out_179_[0]),
		.chany_top_in_181_(cby_0__1__0_chany_out_181_[0]),
		.chany_top_in_183_(cby_0__1__0_chany_out_183_[0]),
		.chany_top_in_185_(cby_0__1__0_chany_out_185_[0]),
		.chany_top_in_187_(cby_0__1__0_chany_out_187_[0]),
		.chany_top_in_189_(cby_0__1__0_chany_out_189_[0]),
		.chany_top_in_191_(cby_0__1__0_chany_out_191_[0]),
		.chany_top_in_193_(cby_0__1__0_chany_out_193_[0]),
		.chany_top_in_195_(cby_0__1__0_chany_out_195_[0]),
		.chany_top_in_197_(cby_0__1__0_chany_out_197_[0]),
		.chany_top_in_199_(cby_0__1__0_chany_out_199_[0]),
		.top_left_grid_pin_1_(grid_io_left_0_right_width_0_height_0__pin_1_lower[0]),
		.chanx_right_in_1_(cbx_1__0__0_chanx_out_1_[0]),
		.chanx_right_in_3_(cbx_1__0__0_chanx_out_3_[0]),
		.chanx_right_in_5_(cbx_1__0__0_chanx_out_5_[0]),
		.chanx_right_in_7_(cbx_1__0__0_chanx_out_7_[0]),
		.chanx_right_in_9_(cbx_1__0__0_chanx_out_9_[0]),
		.chanx_right_in_11_(cbx_1__0__0_chanx_out_11_[0]),
		.chanx_right_in_13_(cbx_1__0__0_chanx_out_13_[0]),
		.chanx_right_in_15_(cbx_1__0__0_chanx_out_15_[0]),
		.chanx_right_in_17_(cbx_1__0__0_chanx_out_17_[0]),
		.chanx_right_in_19_(cbx_1__0__0_chanx_out_19_[0]),
		.chanx_right_in_21_(cbx_1__0__0_chanx_out_21_[0]),
		.chanx_right_in_23_(cbx_1__0__0_chanx_out_23_[0]),
		.chanx_right_in_25_(cbx_1__0__0_chanx_out_25_[0]),
		.chanx_right_in_27_(cbx_1__0__0_chanx_out_27_[0]),
		.chanx_right_in_29_(cbx_1__0__0_chanx_out_29_[0]),
		.chanx_right_in_31_(cbx_1__0__0_chanx_out_31_[0]),
		.chanx_right_in_33_(cbx_1__0__0_chanx_out_33_[0]),
		.chanx_right_in_35_(cbx_1__0__0_chanx_out_35_[0]),
		.chanx_right_in_37_(cbx_1__0__0_chanx_out_37_[0]),
		.chanx_right_in_39_(cbx_1__0__0_chanx_out_39_[0]),
		.chanx_right_in_41_(cbx_1__0__0_chanx_out_41_[0]),
		.chanx_right_in_43_(cbx_1__0__0_chanx_out_43_[0]),
		.chanx_right_in_45_(cbx_1__0__0_chanx_out_45_[0]),
		.chanx_right_in_47_(cbx_1__0__0_chanx_out_47_[0]),
		.chanx_right_in_49_(cbx_1__0__0_chanx_out_49_[0]),
		.chanx_right_in_51_(cbx_1__0__0_chanx_out_51_[0]),
		.chanx_right_in_53_(cbx_1__0__0_chanx_out_53_[0]),
		.chanx_right_in_55_(cbx_1__0__0_chanx_out_55_[0]),
		.chanx_right_in_57_(cbx_1__0__0_chanx_out_57_[0]),
		.chanx_right_in_59_(cbx_1__0__0_chanx_out_59_[0]),
		.chanx_right_in_61_(cbx_1__0__0_chanx_out_61_[0]),
		.chanx_right_in_63_(cbx_1__0__0_chanx_out_63_[0]),
		.chanx_right_in_65_(cbx_1__0__0_chanx_out_65_[0]),
		.chanx_right_in_67_(cbx_1__0__0_chanx_out_67_[0]),
		.chanx_right_in_69_(cbx_1__0__0_chanx_out_69_[0]),
		.chanx_right_in_71_(cbx_1__0__0_chanx_out_71_[0]),
		.chanx_right_in_73_(cbx_1__0__0_chanx_out_73_[0]),
		.chanx_right_in_75_(cbx_1__0__0_chanx_out_75_[0]),
		.chanx_right_in_77_(cbx_1__0__0_chanx_out_77_[0]),
		.chanx_right_in_79_(cbx_1__0__0_chanx_out_79_[0]),
		.chanx_right_in_81_(cbx_1__0__0_chanx_out_81_[0]),
		.chanx_right_in_83_(cbx_1__0__0_chanx_out_83_[0]),
		.chanx_right_in_85_(cbx_1__0__0_chanx_out_85_[0]),
		.chanx_right_in_87_(cbx_1__0__0_chanx_out_87_[0]),
		.chanx_right_in_89_(cbx_1__0__0_chanx_out_89_[0]),
		.chanx_right_in_91_(cbx_1__0__0_chanx_out_91_[0]),
		.chanx_right_in_93_(cbx_1__0__0_chanx_out_93_[0]),
		.chanx_right_in_95_(cbx_1__0__0_chanx_out_95_[0]),
		.chanx_right_in_97_(cbx_1__0__0_chanx_out_97_[0]),
		.chanx_right_in_99_(cbx_1__0__0_chanx_out_99_[0]),
		.chanx_right_in_101_(cbx_1__0__0_chanx_out_101_[0]),
		.chanx_right_in_103_(cbx_1__0__0_chanx_out_103_[0]),
		.chanx_right_in_105_(cbx_1__0__0_chanx_out_105_[0]),
		.chanx_right_in_107_(cbx_1__0__0_chanx_out_107_[0]),
		.chanx_right_in_109_(cbx_1__0__0_chanx_out_109_[0]),
		.chanx_right_in_111_(cbx_1__0__0_chanx_out_111_[0]),
		.chanx_right_in_113_(cbx_1__0__0_chanx_out_113_[0]),
		.chanx_right_in_115_(cbx_1__0__0_chanx_out_115_[0]),
		.chanx_right_in_117_(cbx_1__0__0_chanx_out_117_[0]),
		.chanx_right_in_119_(cbx_1__0__0_chanx_out_119_[0]),
		.chanx_right_in_121_(cbx_1__0__0_chanx_out_121_[0]),
		.chanx_right_in_123_(cbx_1__0__0_chanx_out_123_[0]),
		.chanx_right_in_125_(cbx_1__0__0_chanx_out_125_[0]),
		.chanx_right_in_127_(cbx_1__0__0_chanx_out_127_[0]),
		.chanx_right_in_129_(cbx_1__0__0_chanx_out_129_[0]),
		.chanx_right_in_131_(cbx_1__0__0_chanx_out_131_[0]),
		.chanx_right_in_133_(cbx_1__0__0_chanx_out_133_[0]),
		.chanx_right_in_135_(cbx_1__0__0_chanx_out_135_[0]),
		.chanx_right_in_137_(cbx_1__0__0_chanx_out_137_[0]),
		.chanx_right_in_139_(cbx_1__0__0_chanx_out_139_[0]),
		.chanx_right_in_141_(cbx_1__0__0_chanx_out_141_[0]),
		.chanx_right_in_143_(cbx_1__0__0_chanx_out_143_[0]),
		.chanx_right_in_145_(cbx_1__0__0_chanx_out_145_[0]),
		.chanx_right_in_147_(cbx_1__0__0_chanx_out_147_[0]),
		.chanx_right_in_149_(cbx_1__0__0_chanx_out_149_[0]),
		.chanx_right_in_151_(cbx_1__0__0_chanx_out_151_[0]),
		.chanx_right_in_153_(cbx_1__0__0_chanx_out_153_[0]),
		.chanx_right_in_155_(cbx_1__0__0_chanx_out_155_[0]),
		.chanx_right_in_157_(cbx_1__0__0_chanx_out_157_[0]),
		.chanx_right_in_159_(cbx_1__0__0_chanx_out_159_[0]),
		.chanx_right_in_161_(cbx_1__0__0_chanx_out_161_[0]),
		.chanx_right_in_163_(cbx_1__0__0_chanx_out_163_[0]),
		.chanx_right_in_165_(cbx_1__0__0_chanx_out_165_[0]),
		.chanx_right_in_167_(cbx_1__0__0_chanx_out_167_[0]),
		.chanx_right_in_169_(cbx_1__0__0_chanx_out_169_[0]),
		.chanx_right_in_171_(cbx_1__0__0_chanx_out_171_[0]),
		.chanx_right_in_173_(cbx_1__0__0_chanx_out_173_[0]),
		.chanx_right_in_175_(cbx_1__0__0_chanx_out_175_[0]),
		.chanx_right_in_177_(cbx_1__0__0_chanx_out_177_[0]),
		.chanx_right_in_179_(cbx_1__0__0_chanx_out_179_[0]),
		.chanx_right_in_181_(cbx_1__0__0_chanx_out_181_[0]),
		.chanx_right_in_183_(cbx_1__0__0_chanx_out_183_[0]),
		.chanx_right_in_185_(cbx_1__0__0_chanx_out_185_[0]),
		.chanx_right_in_187_(cbx_1__0__0_chanx_out_187_[0]),
		.chanx_right_in_189_(cbx_1__0__0_chanx_out_189_[0]),
		.chanx_right_in_191_(cbx_1__0__0_chanx_out_191_[0]),
		.chanx_right_in_193_(cbx_1__0__0_chanx_out_193_[0]),
		.chanx_right_in_195_(cbx_1__0__0_chanx_out_195_[0]),
		.chanx_right_in_197_(cbx_1__0__0_chanx_out_197_[0]),
		.chanx_right_in_199_(cbx_1__0__0_chanx_out_199_[0]),
		.right_top_grid_pin_54_(grid_clb_spypad_0_bottom_width_0_height_0__pin_54_upper[0]),
		.right_top_grid_pin_55_(grid_clb_spypad_0_bottom_width_0_height_0__pin_55_upper[0]),
		.right_top_grid_pin_56_(grid_clb_spypad_0_bottom_width_0_height_0__pin_56_upper[0]),
		.right_top_grid_pin_57_(grid_clb_spypad_0_bottom_width_0_height_0__pin_57_upper[0]),
		.right_top_grid_pin_58_(grid_clb_spypad_0_bottom_width_0_height_0__pin_58_upper[0]),
		.right_top_grid_pin_59_(grid_clb_spypad_0_bottom_width_0_height_0__pin_59_upper[0]),
		.right_top_grid_pin_60_(grid_clb_spypad_0_bottom_width_0_height_0__pin_60_upper[0]),
		.right_top_grid_pin_61_(grid_clb_spypad_0_bottom_width_0_height_0__pin_61_upper[0]),
		.right_top_grid_pin_62_(grid_clb_spypad_0_bottom_width_0_height_0__pin_62_upper[0]),
		.right_top_grid_pin_63_(grid_clb_spypad_0_bottom_width_0_height_0__pin_63_upper[0]),
		.right_top_grid_pin_66_(grid_clb_spypad_0_bottom_width_0_height_0__pin_66_upper[0]),
		.right_top_grid_pin_67_(grid_clb_spypad_0_bottom_width_0_height_0__pin_67_upper[0]),
		.right_bottom_grid_pin_1_(grid_io_bottom_0_top_width_0_height_0__pin_1_upper[0]),
		.ccff_head(grid_io_left_1_ccff_tail[0]),
		.chany_top_out_0_(sb_0__0__0_chany_top_out_0_[0]),
		.chany_top_out_2_(sb_0__0__0_chany_top_out_2_[0]),
		.chany_top_out_4_(sb_0__0__0_chany_top_out_4_[0]),
		.chany_top_out_6_(sb_0__0__0_chany_top_out_6_[0]),
		.chany_top_out_8_(sb_0__0__0_chany_top_out_8_[0]),
		.chany_top_out_10_(sb_0__0__0_chany_top_out_10_[0]),
		.chany_top_out_12_(sb_0__0__0_chany_top_out_12_[0]),
		.chany_top_out_14_(sb_0__0__0_chany_top_out_14_[0]),
		.chany_top_out_16_(sb_0__0__0_chany_top_out_16_[0]),
		.chany_top_out_18_(sb_0__0__0_chany_top_out_18_[0]),
		.chany_top_out_20_(sb_0__0__0_chany_top_out_20_[0]),
		.chany_top_out_22_(sb_0__0__0_chany_top_out_22_[0]),
		.chany_top_out_24_(sb_0__0__0_chany_top_out_24_[0]),
		.chany_top_out_26_(sb_0__0__0_chany_top_out_26_[0]),
		.chany_top_out_28_(sb_0__0__0_chany_top_out_28_[0]),
		.chany_top_out_30_(sb_0__0__0_chany_top_out_30_[0]),
		.chany_top_out_32_(sb_0__0__0_chany_top_out_32_[0]),
		.chany_top_out_34_(sb_0__0__0_chany_top_out_34_[0]),
		.chany_top_out_36_(sb_0__0__0_chany_top_out_36_[0]),
		.chany_top_out_38_(sb_0__0__0_chany_top_out_38_[0]),
		.chany_top_out_40_(sb_0__0__0_chany_top_out_40_[0]),
		.chany_top_out_42_(sb_0__0__0_chany_top_out_42_[0]),
		.chany_top_out_44_(sb_0__0__0_chany_top_out_44_[0]),
		.chany_top_out_46_(sb_0__0__0_chany_top_out_46_[0]),
		.chany_top_out_48_(sb_0__0__0_chany_top_out_48_[0]),
		.chany_top_out_50_(sb_0__0__0_chany_top_out_50_[0]),
		.chany_top_out_52_(sb_0__0__0_chany_top_out_52_[0]),
		.chany_top_out_54_(sb_0__0__0_chany_top_out_54_[0]),
		.chany_top_out_56_(sb_0__0__0_chany_top_out_56_[0]),
		.chany_top_out_58_(sb_0__0__0_chany_top_out_58_[0]),
		.chany_top_out_60_(sb_0__0__0_chany_top_out_60_[0]),
		.chany_top_out_62_(sb_0__0__0_chany_top_out_62_[0]),
		.chany_top_out_64_(sb_0__0__0_chany_top_out_64_[0]),
		.chany_top_out_66_(sb_0__0__0_chany_top_out_66_[0]),
		.chany_top_out_68_(sb_0__0__0_chany_top_out_68_[0]),
		.chany_top_out_70_(sb_0__0__0_chany_top_out_70_[0]),
		.chany_top_out_72_(sb_0__0__0_chany_top_out_72_[0]),
		.chany_top_out_74_(sb_0__0__0_chany_top_out_74_[0]),
		.chany_top_out_76_(sb_0__0__0_chany_top_out_76_[0]),
		.chany_top_out_78_(sb_0__0__0_chany_top_out_78_[0]),
		.chany_top_out_80_(sb_0__0__0_chany_top_out_80_[0]),
		.chany_top_out_82_(sb_0__0__0_chany_top_out_82_[0]),
		.chany_top_out_84_(sb_0__0__0_chany_top_out_84_[0]),
		.chany_top_out_86_(sb_0__0__0_chany_top_out_86_[0]),
		.chany_top_out_88_(sb_0__0__0_chany_top_out_88_[0]),
		.chany_top_out_90_(sb_0__0__0_chany_top_out_90_[0]),
		.chany_top_out_92_(sb_0__0__0_chany_top_out_92_[0]),
		.chany_top_out_94_(sb_0__0__0_chany_top_out_94_[0]),
		.chany_top_out_96_(sb_0__0__0_chany_top_out_96_[0]),
		.chany_top_out_98_(sb_0__0__0_chany_top_out_98_[0]),
		.chany_top_out_100_(sb_0__0__0_chany_top_out_100_[0]),
		.chany_top_out_102_(sb_0__0__0_chany_top_out_102_[0]),
		.chany_top_out_104_(sb_0__0__0_chany_top_out_104_[0]),
		.chany_top_out_106_(sb_0__0__0_chany_top_out_106_[0]),
		.chany_top_out_108_(sb_0__0__0_chany_top_out_108_[0]),
		.chany_top_out_110_(sb_0__0__0_chany_top_out_110_[0]),
		.chany_top_out_112_(sb_0__0__0_chany_top_out_112_[0]),
		.chany_top_out_114_(sb_0__0__0_chany_top_out_114_[0]),
		.chany_top_out_116_(sb_0__0__0_chany_top_out_116_[0]),
		.chany_top_out_118_(sb_0__0__0_chany_top_out_118_[0]),
		.chany_top_out_120_(sb_0__0__0_chany_top_out_120_[0]),
		.chany_top_out_122_(sb_0__0__0_chany_top_out_122_[0]),
		.chany_top_out_124_(sb_0__0__0_chany_top_out_124_[0]),
		.chany_top_out_126_(sb_0__0__0_chany_top_out_126_[0]),
		.chany_top_out_128_(sb_0__0__0_chany_top_out_128_[0]),
		.chany_top_out_130_(sb_0__0__0_chany_top_out_130_[0]),
		.chany_top_out_132_(sb_0__0__0_chany_top_out_132_[0]),
		.chany_top_out_134_(sb_0__0__0_chany_top_out_134_[0]),
		.chany_top_out_136_(sb_0__0__0_chany_top_out_136_[0]),
		.chany_top_out_138_(sb_0__0__0_chany_top_out_138_[0]),
		.chany_top_out_140_(sb_0__0__0_chany_top_out_140_[0]),
		.chany_top_out_142_(sb_0__0__0_chany_top_out_142_[0]),
		.chany_top_out_144_(sb_0__0__0_chany_top_out_144_[0]),
		.chany_top_out_146_(sb_0__0__0_chany_top_out_146_[0]),
		.chany_top_out_148_(sb_0__0__0_chany_top_out_148_[0]),
		.chany_top_out_150_(sb_0__0__0_chany_top_out_150_[0]),
		.chany_top_out_152_(sb_0__0__0_chany_top_out_152_[0]),
		.chany_top_out_154_(sb_0__0__0_chany_top_out_154_[0]),
		.chany_top_out_156_(sb_0__0__0_chany_top_out_156_[0]),
		.chany_top_out_158_(sb_0__0__0_chany_top_out_158_[0]),
		.chany_top_out_160_(sb_0__0__0_chany_top_out_160_[0]),
		.chany_top_out_162_(sb_0__0__0_chany_top_out_162_[0]),
		.chany_top_out_164_(sb_0__0__0_chany_top_out_164_[0]),
		.chany_top_out_166_(sb_0__0__0_chany_top_out_166_[0]),
		.chany_top_out_168_(sb_0__0__0_chany_top_out_168_[0]),
		.chany_top_out_170_(sb_0__0__0_chany_top_out_170_[0]),
		.chany_top_out_172_(sb_0__0__0_chany_top_out_172_[0]),
		.chany_top_out_174_(sb_0__0__0_chany_top_out_174_[0]),
		.chany_top_out_176_(sb_0__0__0_chany_top_out_176_[0]),
		.chany_top_out_178_(sb_0__0__0_chany_top_out_178_[0]),
		.chany_top_out_180_(sb_0__0__0_chany_top_out_180_[0]),
		.chany_top_out_182_(sb_0__0__0_chany_top_out_182_[0]),
		.chany_top_out_184_(sb_0__0__0_chany_top_out_184_[0]),
		.chany_top_out_186_(sb_0__0__0_chany_top_out_186_[0]),
		.chany_top_out_188_(sb_0__0__0_chany_top_out_188_[0]),
		.chany_top_out_190_(sb_0__0__0_chany_top_out_190_[0]),
		.chany_top_out_192_(sb_0__0__0_chany_top_out_192_[0]),
		.chany_top_out_194_(sb_0__0__0_chany_top_out_194_[0]),
		.chany_top_out_196_(sb_0__0__0_chany_top_out_196_[0]),
		.chany_top_out_198_(sb_0__0__0_chany_top_out_198_[0]),
		.chanx_right_out_0_(sb_0__0__0_chanx_right_out_0_[0]),
		.chanx_right_out_2_(sb_0__0__0_chanx_right_out_2_[0]),
		.chanx_right_out_4_(sb_0__0__0_chanx_right_out_4_[0]),
		.chanx_right_out_6_(sb_0__0__0_chanx_right_out_6_[0]),
		.chanx_right_out_8_(sb_0__0__0_chanx_right_out_8_[0]),
		.chanx_right_out_10_(sb_0__0__0_chanx_right_out_10_[0]),
		.chanx_right_out_12_(sb_0__0__0_chanx_right_out_12_[0]),
		.chanx_right_out_14_(sb_0__0__0_chanx_right_out_14_[0]),
		.chanx_right_out_16_(sb_0__0__0_chanx_right_out_16_[0]),
		.chanx_right_out_18_(sb_0__0__0_chanx_right_out_18_[0]),
		.chanx_right_out_20_(sb_0__0__0_chanx_right_out_20_[0]),
		.chanx_right_out_22_(sb_0__0__0_chanx_right_out_22_[0]),
		.chanx_right_out_24_(sb_0__0__0_chanx_right_out_24_[0]),
		.chanx_right_out_26_(sb_0__0__0_chanx_right_out_26_[0]),
		.chanx_right_out_28_(sb_0__0__0_chanx_right_out_28_[0]),
		.chanx_right_out_30_(sb_0__0__0_chanx_right_out_30_[0]),
		.chanx_right_out_32_(sb_0__0__0_chanx_right_out_32_[0]),
		.chanx_right_out_34_(sb_0__0__0_chanx_right_out_34_[0]),
		.chanx_right_out_36_(sb_0__0__0_chanx_right_out_36_[0]),
		.chanx_right_out_38_(sb_0__0__0_chanx_right_out_38_[0]),
		.chanx_right_out_40_(sb_0__0__0_chanx_right_out_40_[0]),
		.chanx_right_out_42_(sb_0__0__0_chanx_right_out_42_[0]),
		.chanx_right_out_44_(sb_0__0__0_chanx_right_out_44_[0]),
		.chanx_right_out_46_(sb_0__0__0_chanx_right_out_46_[0]),
		.chanx_right_out_48_(sb_0__0__0_chanx_right_out_48_[0]),
		.chanx_right_out_50_(sb_0__0__0_chanx_right_out_50_[0]),
		.chanx_right_out_52_(sb_0__0__0_chanx_right_out_52_[0]),
		.chanx_right_out_54_(sb_0__0__0_chanx_right_out_54_[0]),
		.chanx_right_out_56_(sb_0__0__0_chanx_right_out_56_[0]),
		.chanx_right_out_58_(sb_0__0__0_chanx_right_out_58_[0]),
		.chanx_right_out_60_(sb_0__0__0_chanx_right_out_60_[0]),
		.chanx_right_out_62_(sb_0__0__0_chanx_right_out_62_[0]),
		.chanx_right_out_64_(sb_0__0__0_chanx_right_out_64_[0]),
		.chanx_right_out_66_(sb_0__0__0_chanx_right_out_66_[0]),
		.chanx_right_out_68_(sb_0__0__0_chanx_right_out_68_[0]),
		.chanx_right_out_70_(sb_0__0__0_chanx_right_out_70_[0]),
		.chanx_right_out_72_(sb_0__0__0_chanx_right_out_72_[0]),
		.chanx_right_out_74_(sb_0__0__0_chanx_right_out_74_[0]),
		.chanx_right_out_76_(sb_0__0__0_chanx_right_out_76_[0]),
		.chanx_right_out_78_(sb_0__0__0_chanx_right_out_78_[0]),
		.chanx_right_out_80_(sb_0__0__0_chanx_right_out_80_[0]),
		.chanx_right_out_82_(sb_0__0__0_chanx_right_out_82_[0]),
		.chanx_right_out_84_(sb_0__0__0_chanx_right_out_84_[0]),
		.chanx_right_out_86_(sb_0__0__0_chanx_right_out_86_[0]),
		.chanx_right_out_88_(sb_0__0__0_chanx_right_out_88_[0]),
		.chanx_right_out_90_(sb_0__0__0_chanx_right_out_90_[0]),
		.chanx_right_out_92_(sb_0__0__0_chanx_right_out_92_[0]),
		.chanx_right_out_94_(sb_0__0__0_chanx_right_out_94_[0]),
		.chanx_right_out_96_(sb_0__0__0_chanx_right_out_96_[0]),
		.chanx_right_out_98_(sb_0__0__0_chanx_right_out_98_[0]),
		.chanx_right_out_100_(sb_0__0__0_chanx_right_out_100_[0]),
		.chanx_right_out_102_(sb_0__0__0_chanx_right_out_102_[0]),
		.chanx_right_out_104_(sb_0__0__0_chanx_right_out_104_[0]),
		.chanx_right_out_106_(sb_0__0__0_chanx_right_out_106_[0]),
		.chanx_right_out_108_(sb_0__0__0_chanx_right_out_108_[0]),
		.chanx_right_out_110_(sb_0__0__0_chanx_right_out_110_[0]),
		.chanx_right_out_112_(sb_0__0__0_chanx_right_out_112_[0]),
		.chanx_right_out_114_(sb_0__0__0_chanx_right_out_114_[0]),
		.chanx_right_out_116_(sb_0__0__0_chanx_right_out_116_[0]),
		.chanx_right_out_118_(sb_0__0__0_chanx_right_out_118_[0]),
		.chanx_right_out_120_(sb_0__0__0_chanx_right_out_120_[0]),
		.chanx_right_out_122_(sb_0__0__0_chanx_right_out_122_[0]),
		.chanx_right_out_124_(sb_0__0__0_chanx_right_out_124_[0]),
		.chanx_right_out_126_(sb_0__0__0_chanx_right_out_126_[0]),
		.chanx_right_out_128_(sb_0__0__0_chanx_right_out_128_[0]),
		.chanx_right_out_130_(sb_0__0__0_chanx_right_out_130_[0]),
		.chanx_right_out_132_(sb_0__0__0_chanx_right_out_132_[0]),
		.chanx_right_out_134_(sb_0__0__0_chanx_right_out_134_[0]),
		.chanx_right_out_136_(sb_0__0__0_chanx_right_out_136_[0]),
		.chanx_right_out_138_(sb_0__0__0_chanx_right_out_138_[0]),
		.chanx_right_out_140_(sb_0__0__0_chanx_right_out_140_[0]),
		.chanx_right_out_142_(sb_0__0__0_chanx_right_out_142_[0]),
		.chanx_right_out_144_(sb_0__0__0_chanx_right_out_144_[0]),
		.chanx_right_out_146_(sb_0__0__0_chanx_right_out_146_[0]),
		.chanx_right_out_148_(sb_0__0__0_chanx_right_out_148_[0]),
		.chanx_right_out_150_(sb_0__0__0_chanx_right_out_150_[0]),
		.chanx_right_out_152_(sb_0__0__0_chanx_right_out_152_[0]),
		.chanx_right_out_154_(sb_0__0__0_chanx_right_out_154_[0]),
		.chanx_right_out_156_(sb_0__0__0_chanx_right_out_156_[0]),
		.chanx_right_out_158_(sb_0__0__0_chanx_right_out_158_[0]),
		.chanx_right_out_160_(sb_0__0__0_chanx_right_out_160_[0]),
		.chanx_right_out_162_(sb_0__0__0_chanx_right_out_162_[0]),
		.chanx_right_out_164_(sb_0__0__0_chanx_right_out_164_[0]),
		.chanx_right_out_166_(sb_0__0__0_chanx_right_out_166_[0]),
		.chanx_right_out_168_(sb_0__0__0_chanx_right_out_168_[0]),
		.chanx_right_out_170_(sb_0__0__0_chanx_right_out_170_[0]),
		.chanx_right_out_172_(sb_0__0__0_chanx_right_out_172_[0]),
		.chanx_right_out_174_(sb_0__0__0_chanx_right_out_174_[0]),
		.chanx_right_out_176_(sb_0__0__0_chanx_right_out_176_[0]),
		.chanx_right_out_178_(sb_0__0__0_chanx_right_out_178_[0]),
		.chanx_right_out_180_(sb_0__0__0_chanx_right_out_180_[0]),
		.chanx_right_out_182_(sb_0__0__0_chanx_right_out_182_[0]),
		.chanx_right_out_184_(sb_0__0__0_chanx_right_out_184_[0]),
		.chanx_right_out_186_(sb_0__0__0_chanx_right_out_186_[0]),
		.chanx_right_out_188_(sb_0__0__0_chanx_right_out_188_[0]),
		.chanx_right_out_190_(sb_0__0__0_chanx_right_out_190_[0]),
		.chanx_right_out_192_(sb_0__0__0_chanx_right_out_192_[0]),
		.chanx_right_out_194_(sb_0__0__0_chanx_right_out_194_[0]),
		.chanx_right_out_196_(sb_0__0__0_chanx_right_out_196_[0]),
		.chanx_right_out_198_(sb_0__0__0_chanx_right_out_198_[0]),
		.ccff_tail(sb_0__0__0_ccff_tail[0]));

	sb_0__1_ sb_0__1_ (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.chany_top_in_1_(cby_0__1__1_chany_out_1_[0]),
		.chany_top_in_3_(cby_0__1__1_chany_out_3_[0]),
		.chany_top_in_5_(cby_0__1__1_chany_out_5_[0]),
		.chany_top_in_7_(cby_0__1__1_chany_out_7_[0]),
		.chany_top_in_9_(cby_0__1__1_chany_out_9_[0]),
		.chany_top_in_11_(cby_0__1__1_chany_out_11_[0]),
		.chany_top_in_13_(cby_0__1__1_chany_out_13_[0]),
		.chany_top_in_15_(cby_0__1__1_chany_out_15_[0]),
		.chany_top_in_17_(cby_0__1__1_chany_out_17_[0]),
		.chany_top_in_19_(cby_0__1__1_chany_out_19_[0]),
		.chany_top_in_21_(cby_0__1__1_chany_out_21_[0]),
		.chany_top_in_23_(cby_0__1__1_chany_out_23_[0]),
		.chany_top_in_25_(cby_0__1__1_chany_out_25_[0]),
		.chany_top_in_27_(cby_0__1__1_chany_out_27_[0]),
		.chany_top_in_29_(cby_0__1__1_chany_out_29_[0]),
		.chany_top_in_31_(cby_0__1__1_chany_out_31_[0]),
		.chany_top_in_33_(cby_0__1__1_chany_out_33_[0]),
		.chany_top_in_35_(cby_0__1__1_chany_out_35_[0]),
		.chany_top_in_37_(cby_0__1__1_chany_out_37_[0]),
		.chany_top_in_39_(cby_0__1__1_chany_out_39_[0]),
		.chany_top_in_41_(cby_0__1__1_chany_out_41_[0]),
		.chany_top_in_43_(cby_0__1__1_chany_out_43_[0]),
		.chany_top_in_45_(cby_0__1__1_chany_out_45_[0]),
		.chany_top_in_47_(cby_0__1__1_chany_out_47_[0]),
		.chany_top_in_49_(cby_0__1__1_chany_out_49_[0]),
		.chany_top_in_51_(cby_0__1__1_chany_out_51_[0]),
		.chany_top_in_53_(cby_0__1__1_chany_out_53_[0]),
		.chany_top_in_55_(cby_0__1__1_chany_out_55_[0]),
		.chany_top_in_57_(cby_0__1__1_chany_out_57_[0]),
		.chany_top_in_59_(cby_0__1__1_chany_out_59_[0]),
		.chany_top_in_61_(cby_0__1__1_chany_out_61_[0]),
		.chany_top_in_63_(cby_0__1__1_chany_out_63_[0]),
		.chany_top_in_65_(cby_0__1__1_chany_out_65_[0]),
		.chany_top_in_67_(cby_0__1__1_chany_out_67_[0]),
		.chany_top_in_69_(cby_0__1__1_chany_out_69_[0]),
		.chany_top_in_71_(cby_0__1__1_chany_out_71_[0]),
		.chany_top_in_73_(cby_0__1__1_chany_out_73_[0]),
		.chany_top_in_75_(cby_0__1__1_chany_out_75_[0]),
		.chany_top_in_77_(cby_0__1__1_chany_out_77_[0]),
		.chany_top_in_79_(cby_0__1__1_chany_out_79_[0]),
		.chany_top_in_81_(cby_0__1__1_chany_out_81_[0]),
		.chany_top_in_83_(cby_0__1__1_chany_out_83_[0]),
		.chany_top_in_85_(cby_0__1__1_chany_out_85_[0]),
		.chany_top_in_87_(cby_0__1__1_chany_out_87_[0]),
		.chany_top_in_89_(cby_0__1__1_chany_out_89_[0]),
		.chany_top_in_91_(cby_0__1__1_chany_out_91_[0]),
		.chany_top_in_93_(cby_0__1__1_chany_out_93_[0]),
		.chany_top_in_95_(cby_0__1__1_chany_out_95_[0]),
		.chany_top_in_97_(cby_0__1__1_chany_out_97_[0]),
		.chany_top_in_99_(cby_0__1__1_chany_out_99_[0]),
		.chany_top_in_101_(cby_0__1__1_chany_out_101_[0]),
		.chany_top_in_103_(cby_0__1__1_chany_out_103_[0]),
		.chany_top_in_105_(cby_0__1__1_chany_out_105_[0]),
		.chany_top_in_107_(cby_0__1__1_chany_out_107_[0]),
		.chany_top_in_109_(cby_0__1__1_chany_out_109_[0]),
		.chany_top_in_111_(cby_0__1__1_chany_out_111_[0]),
		.chany_top_in_113_(cby_0__1__1_chany_out_113_[0]),
		.chany_top_in_115_(cby_0__1__1_chany_out_115_[0]),
		.chany_top_in_117_(cby_0__1__1_chany_out_117_[0]),
		.chany_top_in_119_(cby_0__1__1_chany_out_119_[0]),
		.chany_top_in_121_(cby_0__1__1_chany_out_121_[0]),
		.chany_top_in_123_(cby_0__1__1_chany_out_123_[0]),
		.chany_top_in_125_(cby_0__1__1_chany_out_125_[0]),
		.chany_top_in_127_(cby_0__1__1_chany_out_127_[0]),
		.chany_top_in_129_(cby_0__1__1_chany_out_129_[0]),
		.chany_top_in_131_(cby_0__1__1_chany_out_131_[0]),
		.chany_top_in_133_(cby_0__1__1_chany_out_133_[0]),
		.chany_top_in_135_(cby_0__1__1_chany_out_135_[0]),
		.chany_top_in_137_(cby_0__1__1_chany_out_137_[0]),
		.chany_top_in_139_(cby_0__1__1_chany_out_139_[0]),
		.chany_top_in_141_(cby_0__1__1_chany_out_141_[0]),
		.chany_top_in_143_(cby_0__1__1_chany_out_143_[0]),
		.chany_top_in_145_(cby_0__1__1_chany_out_145_[0]),
		.chany_top_in_147_(cby_0__1__1_chany_out_147_[0]),
		.chany_top_in_149_(cby_0__1__1_chany_out_149_[0]),
		.chany_top_in_151_(cby_0__1__1_chany_out_151_[0]),
		.chany_top_in_153_(cby_0__1__1_chany_out_153_[0]),
		.chany_top_in_155_(cby_0__1__1_chany_out_155_[0]),
		.chany_top_in_157_(cby_0__1__1_chany_out_157_[0]),
		.chany_top_in_159_(cby_0__1__1_chany_out_159_[0]),
		.chany_top_in_161_(cby_0__1__1_chany_out_161_[0]),
		.chany_top_in_163_(cby_0__1__1_chany_out_163_[0]),
		.chany_top_in_165_(cby_0__1__1_chany_out_165_[0]),
		.chany_top_in_167_(cby_0__1__1_chany_out_167_[0]),
		.chany_top_in_169_(cby_0__1__1_chany_out_169_[0]),
		.chany_top_in_171_(cby_0__1__1_chany_out_171_[0]),
		.chany_top_in_173_(cby_0__1__1_chany_out_173_[0]),
		.chany_top_in_175_(cby_0__1__1_chany_out_175_[0]),
		.chany_top_in_177_(cby_0__1__1_chany_out_177_[0]),
		.chany_top_in_179_(cby_0__1__1_chany_out_179_[0]),
		.chany_top_in_181_(cby_0__1__1_chany_out_181_[0]),
		.chany_top_in_183_(cby_0__1__1_chany_out_183_[0]),
		.chany_top_in_185_(cby_0__1__1_chany_out_185_[0]),
		.chany_top_in_187_(cby_0__1__1_chany_out_187_[0]),
		.chany_top_in_189_(cby_0__1__1_chany_out_189_[0]),
		.chany_top_in_191_(cby_0__1__1_chany_out_191_[0]),
		.chany_top_in_193_(cby_0__1__1_chany_out_193_[0]),
		.chany_top_in_195_(cby_0__1__1_chany_out_195_[0]),
		.chany_top_in_197_(cby_0__1__1_chany_out_197_[0]),
		.chany_top_in_199_(cby_0__1__1_chany_out_199_[0]),
		.top_left_grid_pin_1_(grid_io_left_1_right_width_0_height_0__pin_1_lower[0]),
		.chanx_right_in_1_(cbx_1__1__0_chanx_out_1_[0]),
		.chanx_right_in_3_(cbx_1__1__0_chanx_out_3_[0]),
		.chanx_right_in_5_(cbx_1__1__0_chanx_out_5_[0]),
		.chanx_right_in_7_(cbx_1__1__0_chanx_out_7_[0]),
		.chanx_right_in_9_(cbx_1__1__0_chanx_out_9_[0]),
		.chanx_right_in_11_(cbx_1__1__0_chanx_out_11_[0]),
		.chanx_right_in_13_(cbx_1__1__0_chanx_out_13_[0]),
		.chanx_right_in_15_(cbx_1__1__0_chanx_out_15_[0]),
		.chanx_right_in_17_(cbx_1__1__0_chanx_out_17_[0]),
		.chanx_right_in_19_(cbx_1__1__0_chanx_out_19_[0]),
		.chanx_right_in_21_(cbx_1__1__0_chanx_out_21_[0]),
		.chanx_right_in_23_(cbx_1__1__0_chanx_out_23_[0]),
		.chanx_right_in_25_(cbx_1__1__0_chanx_out_25_[0]),
		.chanx_right_in_27_(cbx_1__1__0_chanx_out_27_[0]),
		.chanx_right_in_29_(cbx_1__1__0_chanx_out_29_[0]),
		.chanx_right_in_31_(cbx_1__1__0_chanx_out_31_[0]),
		.chanx_right_in_33_(cbx_1__1__0_chanx_out_33_[0]),
		.chanx_right_in_35_(cbx_1__1__0_chanx_out_35_[0]),
		.chanx_right_in_37_(cbx_1__1__0_chanx_out_37_[0]),
		.chanx_right_in_39_(cbx_1__1__0_chanx_out_39_[0]),
		.chanx_right_in_41_(cbx_1__1__0_chanx_out_41_[0]),
		.chanx_right_in_43_(cbx_1__1__0_chanx_out_43_[0]),
		.chanx_right_in_45_(cbx_1__1__0_chanx_out_45_[0]),
		.chanx_right_in_47_(cbx_1__1__0_chanx_out_47_[0]),
		.chanx_right_in_49_(cbx_1__1__0_chanx_out_49_[0]),
		.chanx_right_in_51_(cbx_1__1__0_chanx_out_51_[0]),
		.chanx_right_in_53_(cbx_1__1__0_chanx_out_53_[0]),
		.chanx_right_in_55_(cbx_1__1__0_chanx_out_55_[0]),
		.chanx_right_in_57_(cbx_1__1__0_chanx_out_57_[0]),
		.chanx_right_in_59_(cbx_1__1__0_chanx_out_59_[0]),
		.chanx_right_in_61_(cbx_1__1__0_chanx_out_61_[0]),
		.chanx_right_in_63_(cbx_1__1__0_chanx_out_63_[0]),
		.chanx_right_in_65_(cbx_1__1__0_chanx_out_65_[0]),
		.chanx_right_in_67_(cbx_1__1__0_chanx_out_67_[0]),
		.chanx_right_in_69_(cbx_1__1__0_chanx_out_69_[0]),
		.chanx_right_in_71_(cbx_1__1__0_chanx_out_71_[0]),
		.chanx_right_in_73_(cbx_1__1__0_chanx_out_73_[0]),
		.chanx_right_in_75_(cbx_1__1__0_chanx_out_75_[0]),
		.chanx_right_in_77_(cbx_1__1__0_chanx_out_77_[0]),
		.chanx_right_in_79_(cbx_1__1__0_chanx_out_79_[0]),
		.chanx_right_in_81_(cbx_1__1__0_chanx_out_81_[0]),
		.chanx_right_in_83_(cbx_1__1__0_chanx_out_83_[0]),
		.chanx_right_in_85_(cbx_1__1__0_chanx_out_85_[0]),
		.chanx_right_in_87_(cbx_1__1__0_chanx_out_87_[0]),
		.chanx_right_in_89_(cbx_1__1__0_chanx_out_89_[0]),
		.chanx_right_in_91_(cbx_1__1__0_chanx_out_91_[0]),
		.chanx_right_in_93_(cbx_1__1__0_chanx_out_93_[0]),
		.chanx_right_in_95_(cbx_1__1__0_chanx_out_95_[0]),
		.chanx_right_in_97_(cbx_1__1__0_chanx_out_97_[0]),
		.chanx_right_in_99_(cbx_1__1__0_chanx_out_99_[0]),
		.chanx_right_in_101_(cbx_1__1__0_chanx_out_101_[0]),
		.chanx_right_in_103_(cbx_1__1__0_chanx_out_103_[0]),
		.chanx_right_in_105_(cbx_1__1__0_chanx_out_105_[0]),
		.chanx_right_in_107_(cbx_1__1__0_chanx_out_107_[0]),
		.chanx_right_in_109_(cbx_1__1__0_chanx_out_109_[0]),
		.chanx_right_in_111_(cbx_1__1__0_chanx_out_111_[0]),
		.chanx_right_in_113_(cbx_1__1__0_chanx_out_113_[0]),
		.chanx_right_in_115_(cbx_1__1__0_chanx_out_115_[0]),
		.chanx_right_in_117_(cbx_1__1__0_chanx_out_117_[0]),
		.chanx_right_in_119_(cbx_1__1__0_chanx_out_119_[0]),
		.chanx_right_in_121_(cbx_1__1__0_chanx_out_121_[0]),
		.chanx_right_in_123_(cbx_1__1__0_chanx_out_123_[0]),
		.chanx_right_in_125_(cbx_1__1__0_chanx_out_125_[0]),
		.chanx_right_in_127_(cbx_1__1__0_chanx_out_127_[0]),
		.chanx_right_in_129_(cbx_1__1__0_chanx_out_129_[0]),
		.chanx_right_in_131_(cbx_1__1__0_chanx_out_131_[0]),
		.chanx_right_in_133_(cbx_1__1__0_chanx_out_133_[0]),
		.chanx_right_in_135_(cbx_1__1__0_chanx_out_135_[0]),
		.chanx_right_in_137_(cbx_1__1__0_chanx_out_137_[0]),
		.chanx_right_in_139_(cbx_1__1__0_chanx_out_139_[0]),
		.chanx_right_in_141_(cbx_1__1__0_chanx_out_141_[0]),
		.chanx_right_in_143_(cbx_1__1__0_chanx_out_143_[0]),
		.chanx_right_in_145_(cbx_1__1__0_chanx_out_145_[0]),
		.chanx_right_in_147_(cbx_1__1__0_chanx_out_147_[0]),
		.chanx_right_in_149_(cbx_1__1__0_chanx_out_149_[0]),
		.chanx_right_in_151_(cbx_1__1__0_chanx_out_151_[0]),
		.chanx_right_in_153_(cbx_1__1__0_chanx_out_153_[0]),
		.chanx_right_in_155_(cbx_1__1__0_chanx_out_155_[0]),
		.chanx_right_in_157_(cbx_1__1__0_chanx_out_157_[0]),
		.chanx_right_in_159_(cbx_1__1__0_chanx_out_159_[0]),
		.chanx_right_in_161_(cbx_1__1__0_chanx_out_161_[0]),
		.chanx_right_in_163_(cbx_1__1__0_chanx_out_163_[0]),
		.chanx_right_in_165_(cbx_1__1__0_chanx_out_165_[0]),
		.chanx_right_in_167_(cbx_1__1__0_chanx_out_167_[0]),
		.chanx_right_in_169_(cbx_1__1__0_chanx_out_169_[0]),
		.chanx_right_in_171_(cbx_1__1__0_chanx_out_171_[0]),
		.chanx_right_in_173_(cbx_1__1__0_chanx_out_173_[0]),
		.chanx_right_in_175_(cbx_1__1__0_chanx_out_175_[0]),
		.chanx_right_in_177_(cbx_1__1__0_chanx_out_177_[0]),
		.chanx_right_in_179_(cbx_1__1__0_chanx_out_179_[0]),
		.chanx_right_in_181_(cbx_1__1__0_chanx_out_181_[0]),
		.chanx_right_in_183_(cbx_1__1__0_chanx_out_183_[0]),
		.chanx_right_in_185_(cbx_1__1__0_chanx_out_185_[0]),
		.chanx_right_in_187_(cbx_1__1__0_chanx_out_187_[0]),
		.chanx_right_in_189_(cbx_1__1__0_chanx_out_189_[0]),
		.chanx_right_in_191_(cbx_1__1__0_chanx_out_191_[0]),
		.chanx_right_in_193_(cbx_1__1__0_chanx_out_193_[0]),
		.chanx_right_in_195_(cbx_1__1__0_chanx_out_195_[0]),
		.chanx_right_in_197_(cbx_1__1__0_chanx_out_197_[0]),
		.chanx_right_in_199_(cbx_1__1__0_chanx_out_199_[0]),
		.right_top_grid_pin_54_(grid_clb_0_bottom_width_0_height_0__pin_54_upper[0]),
		.right_top_grid_pin_55_(grid_clb_0_bottom_width_0_height_0__pin_55_upper[0]),
		.right_top_grid_pin_56_(grid_clb_0_bottom_width_0_height_0__pin_56_upper[0]),
		.right_top_grid_pin_57_(grid_clb_0_bottom_width_0_height_0__pin_57_upper[0]),
		.right_top_grid_pin_58_(grid_clb_0_bottom_width_0_height_0__pin_58_upper[0]),
		.right_top_grid_pin_59_(grid_clb_0_bottom_width_0_height_0__pin_59_upper[0]),
		.right_top_grid_pin_60_(grid_clb_0_bottom_width_0_height_0__pin_60_upper[0]),
		.right_top_grid_pin_61_(grid_clb_0_bottom_width_0_height_0__pin_61_upper[0]),
		.right_top_grid_pin_62_(grid_clb_0_bottom_width_0_height_0__pin_62_upper[0]),
		.right_top_grid_pin_63_(grid_clb_0_bottom_width_0_height_0__pin_63_upper[0]),
		.right_top_grid_pin_66_(grid_clb_0_bottom_width_0_height_0__pin_66_upper[0]),
		.right_top_grid_pin_67_(grid_clb_0_bottom_width_0_height_0__pin_67_upper[0]),
		.chany_bottom_in_0_(cby_0__1__0_chany_out_0_[0]),
		.chany_bottom_in_2_(cby_0__1__0_chany_out_2_[0]),
		.chany_bottom_in_4_(cby_0__1__0_chany_out_4_[0]),
		.chany_bottom_in_6_(cby_0__1__0_chany_out_6_[0]),
		.chany_bottom_in_8_(cby_0__1__0_chany_out_8_[0]),
		.chany_bottom_in_10_(cby_0__1__0_chany_out_10_[0]),
		.chany_bottom_in_12_(cby_0__1__0_chany_out_12_[0]),
		.chany_bottom_in_14_(cby_0__1__0_chany_out_14_[0]),
		.chany_bottom_in_16_(cby_0__1__0_chany_out_16_[0]),
		.chany_bottom_in_18_(cby_0__1__0_chany_out_18_[0]),
		.chany_bottom_in_20_(cby_0__1__0_chany_out_20_[0]),
		.chany_bottom_in_22_(cby_0__1__0_chany_out_22_[0]),
		.chany_bottom_in_24_(cby_0__1__0_chany_out_24_[0]),
		.chany_bottom_in_26_(cby_0__1__0_chany_out_26_[0]),
		.chany_bottom_in_28_(cby_0__1__0_chany_out_28_[0]),
		.chany_bottom_in_30_(cby_0__1__0_chany_out_30_[0]),
		.chany_bottom_in_32_(cby_0__1__0_chany_out_32_[0]),
		.chany_bottom_in_34_(cby_0__1__0_chany_out_34_[0]),
		.chany_bottom_in_36_(cby_0__1__0_chany_out_36_[0]),
		.chany_bottom_in_38_(cby_0__1__0_chany_out_38_[0]),
		.chany_bottom_in_40_(cby_0__1__0_chany_out_40_[0]),
		.chany_bottom_in_42_(cby_0__1__0_chany_out_42_[0]),
		.chany_bottom_in_44_(cby_0__1__0_chany_out_44_[0]),
		.chany_bottom_in_46_(cby_0__1__0_chany_out_46_[0]),
		.chany_bottom_in_48_(cby_0__1__0_chany_out_48_[0]),
		.chany_bottom_in_50_(cby_0__1__0_chany_out_50_[0]),
		.chany_bottom_in_52_(cby_0__1__0_chany_out_52_[0]),
		.chany_bottom_in_54_(cby_0__1__0_chany_out_54_[0]),
		.chany_bottom_in_56_(cby_0__1__0_chany_out_56_[0]),
		.chany_bottom_in_58_(cby_0__1__0_chany_out_58_[0]),
		.chany_bottom_in_60_(cby_0__1__0_chany_out_60_[0]),
		.chany_bottom_in_62_(cby_0__1__0_chany_out_62_[0]),
		.chany_bottom_in_64_(cby_0__1__0_chany_out_64_[0]),
		.chany_bottom_in_66_(cby_0__1__0_chany_out_66_[0]),
		.chany_bottom_in_68_(cby_0__1__0_chany_out_68_[0]),
		.chany_bottom_in_70_(cby_0__1__0_chany_out_70_[0]),
		.chany_bottom_in_72_(cby_0__1__0_chany_out_72_[0]),
		.chany_bottom_in_74_(cby_0__1__0_chany_out_74_[0]),
		.chany_bottom_in_76_(cby_0__1__0_chany_out_76_[0]),
		.chany_bottom_in_78_(cby_0__1__0_chany_out_78_[0]),
		.chany_bottom_in_80_(cby_0__1__0_chany_out_80_[0]),
		.chany_bottom_in_82_(cby_0__1__0_chany_out_82_[0]),
		.chany_bottom_in_84_(cby_0__1__0_chany_out_84_[0]),
		.chany_bottom_in_86_(cby_0__1__0_chany_out_86_[0]),
		.chany_bottom_in_88_(cby_0__1__0_chany_out_88_[0]),
		.chany_bottom_in_90_(cby_0__1__0_chany_out_90_[0]),
		.chany_bottom_in_92_(cby_0__1__0_chany_out_92_[0]),
		.chany_bottom_in_94_(cby_0__1__0_chany_out_94_[0]),
		.chany_bottom_in_96_(cby_0__1__0_chany_out_96_[0]),
		.chany_bottom_in_98_(cby_0__1__0_chany_out_98_[0]),
		.chany_bottom_in_100_(cby_0__1__0_chany_out_100_[0]),
		.chany_bottom_in_102_(cby_0__1__0_chany_out_102_[0]),
		.chany_bottom_in_104_(cby_0__1__0_chany_out_104_[0]),
		.chany_bottom_in_106_(cby_0__1__0_chany_out_106_[0]),
		.chany_bottom_in_108_(cby_0__1__0_chany_out_108_[0]),
		.chany_bottom_in_110_(cby_0__1__0_chany_out_110_[0]),
		.chany_bottom_in_112_(cby_0__1__0_chany_out_112_[0]),
		.chany_bottom_in_114_(cby_0__1__0_chany_out_114_[0]),
		.chany_bottom_in_116_(cby_0__1__0_chany_out_116_[0]),
		.chany_bottom_in_118_(cby_0__1__0_chany_out_118_[0]),
		.chany_bottom_in_120_(cby_0__1__0_chany_out_120_[0]),
		.chany_bottom_in_122_(cby_0__1__0_chany_out_122_[0]),
		.chany_bottom_in_124_(cby_0__1__0_chany_out_124_[0]),
		.chany_bottom_in_126_(cby_0__1__0_chany_out_126_[0]),
		.chany_bottom_in_128_(cby_0__1__0_chany_out_128_[0]),
		.chany_bottom_in_130_(cby_0__1__0_chany_out_130_[0]),
		.chany_bottom_in_132_(cby_0__1__0_chany_out_132_[0]),
		.chany_bottom_in_134_(cby_0__1__0_chany_out_134_[0]),
		.chany_bottom_in_136_(cby_0__1__0_chany_out_136_[0]),
		.chany_bottom_in_138_(cby_0__1__0_chany_out_138_[0]),
		.chany_bottom_in_140_(cby_0__1__0_chany_out_140_[0]),
		.chany_bottom_in_142_(cby_0__1__0_chany_out_142_[0]),
		.chany_bottom_in_144_(cby_0__1__0_chany_out_144_[0]),
		.chany_bottom_in_146_(cby_0__1__0_chany_out_146_[0]),
		.chany_bottom_in_148_(cby_0__1__0_chany_out_148_[0]),
		.chany_bottom_in_150_(cby_0__1__0_chany_out_150_[0]),
		.chany_bottom_in_152_(cby_0__1__0_chany_out_152_[0]),
		.chany_bottom_in_154_(cby_0__1__0_chany_out_154_[0]),
		.chany_bottom_in_156_(cby_0__1__0_chany_out_156_[0]),
		.chany_bottom_in_158_(cby_0__1__0_chany_out_158_[0]),
		.chany_bottom_in_160_(cby_0__1__0_chany_out_160_[0]),
		.chany_bottom_in_162_(cby_0__1__0_chany_out_162_[0]),
		.chany_bottom_in_164_(cby_0__1__0_chany_out_164_[0]),
		.chany_bottom_in_166_(cby_0__1__0_chany_out_166_[0]),
		.chany_bottom_in_168_(cby_0__1__0_chany_out_168_[0]),
		.chany_bottom_in_170_(cby_0__1__0_chany_out_170_[0]),
		.chany_bottom_in_172_(cby_0__1__0_chany_out_172_[0]),
		.chany_bottom_in_174_(cby_0__1__0_chany_out_174_[0]),
		.chany_bottom_in_176_(cby_0__1__0_chany_out_176_[0]),
		.chany_bottom_in_178_(cby_0__1__0_chany_out_178_[0]),
		.chany_bottom_in_180_(cby_0__1__0_chany_out_180_[0]),
		.chany_bottom_in_182_(cby_0__1__0_chany_out_182_[0]),
		.chany_bottom_in_184_(cby_0__1__0_chany_out_184_[0]),
		.chany_bottom_in_186_(cby_0__1__0_chany_out_186_[0]),
		.chany_bottom_in_188_(cby_0__1__0_chany_out_188_[0]),
		.chany_bottom_in_190_(cby_0__1__0_chany_out_190_[0]),
		.chany_bottom_in_192_(cby_0__1__0_chany_out_192_[0]),
		.chany_bottom_in_194_(cby_0__1__0_chany_out_194_[0]),
		.chany_bottom_in_196_(cby_0__1__0_chany_out_196_[0]),
		.chany_bottom_in_198_(cby_0__1__0_chany_out_198_[0]),
		.bottom_left_grid_pin_1_(grid_io_left_0_right_width_0_height_0__pin_1_upper[0]),
		.ccff_head(sb_0__2__0_ccff_tail[0]),
		.chany_top_out_0_(sb_0__1__0_chany_top_out_0_[0]),
		.chany_top_out_2_(sb_0__1__0_chany_top_out_2_[0]),
		.chany_top_out_4_(sb_0__1__0_chany_top_out_4_[0]),
		.chany_top_out_6_(sb_0__1__0_chany_top_out_6_[0]),
		.chany_top_out_8_(sb_0__1__0_chany_top_out_8_[0]),
		.chany_top_out_10_(sb_0__1__0_chany_top_out_10_[0]),
		.chany_top_out_12_(sb_0__1__0_chany_top_out_12_[0]),
		.chany_top_out_14_(sb_0__1__0_chany_top_out_14_[0]),
		.chany_top_out_16_(sb_0__1__0_chany_top_out_16_[0]),
		.chany_top_out_18_(sb_0__1__0_chany_top_out_18_[0]),
		.chany_top_out_20_(sb_0__1__0_chany_top_out_20_[0]),
		.chany_top_out_22_(sb_0__1__0_chany_top_out_22_[0]),
		.chany_top_out_24_(sb_0__1__0_chany_top_out_24_[0]),
		.chany_top_out_26_(sb_0__1__0_chany_top_out_26_[0]),
		.chany_top_out_28_(sb_0__1__0_chany_top_out_28_[0]),
		.chany_top_out_30_(sb_0__1__0_chany_top_out_30_[0]),
		.chany_top_out_32_(sb_0__1__0_chany_top_out_32_[0]),
		.chany_top_out_34_(sb_0__1__0_chany_top_out_34_[0]),
		.chany_top_out_36_(sb_0__1__0_chany_top_out_36_[0]),
		.chany_top_out_38_(sb_0__1__0_chany_top_out_38_[0]),
		.chany_top_out_40_(sb_0__1__0_chany_top_out_40_[0]),
		.chany_top_out_42_(sb_0__1__0_chany_top_out_42_[0]),
		.chany_top_out_44_(sb_0__1__0_chany_top_out_44_[0]),
		.chany_top_out_46_(sb_0__1__0_chany_top_out_46_[0]),
		.chany_top_out_48_(sb_0__1__0_chany_top_out_48_[0]),
		.chany_top_out_50_(sb_0__1__0_chany_top_out_50_[0]),
		.chany_top_out_52_(sb_0__1__0_chany_top_out_52_[0]),
		.chany_top_out_54_(sb_0__1__0_chany_top_out_54_[0]),
		.chany_top_out_56_(sb_0__1__0_chany_top_out_56_[0]),
		.chany_top_out_58_(sb_0__1__0_chany_top_out_58_[0]),
		.chany_top_out_60_(sb_0__1__0_chany_top_out_60_[0]),
		.chany_top_out_62_(sb_0__1__0_chany_top_out_62_[0]),
		.chany_top_out_64_(sb_0__1__0_chany_top_out_64_[0]),
		.chany_top_out_66_(sb_0__1__0_chany_top_out_66_[0]),
		.chany_top_out_68_(sb_0__1__0_chany_top_out_68_[0]),
		.chany_top_out_70_(sb_0__1__0_chany_top_out_70_[0]),
		.chany_top_out_72_(sb_0__1__0_chany_top_out_72_[0]),
		.chany_top_out_74_(sb_0__1__0_chany_top_out_74_[0]),
		.chany_top_out_76_(sb_0__1__0_chany_top_out_76_[0]),
		.chany_top_out_78_(sb_0__1__0_chany_top_out_78_[0]),
		.chany_top_out_80_(sb_0__1__0_chany_top_out_80_[0]),
		.chany_top_out_82_(sb_0__1__0_chany_top_out_82_[0]),
		.chany_top_out_84_(sb_0__1__0_chany_top_out_84_[0]),
		.chany_top_out_86_(sb_0__1__0_chany_top_out_86_[0]),
		.chany_top_out_88_(sb_0__1__0_chany_top_out_88_[0]),
		.chany_top_out_90_(sb_0__1__0_chany_top_out_90_[0]),
		.chany_top_out_92_(sb_0__1__0_chany_top_out_92_[0]),
		.chany_top_out_94_(sb_0__1__0_chany_top_out_94_[0]),
		.chany_top_out_96_(sb_0__1__0_chany_top_out_96_[0]),
		.chany_top_out_98_(sb_0__1__0_chany_top_out_98_[0]),
		.chany_top_out_100_(sb_0__1__0_chany_top_out_100_[0]),
		.chany_top_out_102_(sb_0__1__0_chany_top_out_102_[0]),
		.chany_top_out_104_(sb_0__1__0_chany_top_out_104_[0]),
		.chany_top_out_106_(sb_0__1__0_chany_top_out_106_[0]),
		.chany_top_out_108_(sb_0__1__0_chany_top_out_108_[0]),
		.chany_top_out_110_(sb_0__1__0_chany_top_out_110_[0]),
		.chany_top_out_112_(sb_0__1__0_chany_top_out_112_[0]),
		.chany_top_out_114_(sb_0__1__0_chany_top_out_114_[0]),
		.chany_top_out_116_(sb_0__1__0_chany_top_out_116_[0]),
		.chany_top_out_118_(sb_0__1__0_chany_top_out_118_[0]),
		.chany_top_out_120_(sb_0__1__0_chany_top_out_120_[0]),
		.chany_top_out_122_(sb_0__1__0_chany_top_out_122_[0]),
		.chany_top_out_124_(sb_0__1__0_chany_top_out_124_[0]),
		.chany_top_out_126_(sb_0__1__0_chany_top_out_126_[0]),
		.chany_top_out_128_(sb_0__1__0_chany_top_out_128_[0]),
		.chany_top_out_130_(sb_0__1__0_chany_top_out_130_[0]),
		.chany_top_out_132_(sb_0__1__0_chany_top_out_132_[0]),
		.chany_top_out_134_(sb_0__1__0_chany_top_out_134_[0]),
		.chany_top_out_136_(sb_0__1__0_chany_top_out_136_[0]),
		.chany_top_out_138_(sb_0__1__0_chany_top_out_138_[0]),
		.chany_top_out_140_(sb_0__1__0_chany_top_out_140_[0]),
		.chany_top_out_142_(sb_0__1__0_chany_top_out_142_[0]),
		.chany_top_out_144_(sb_0__1__0_chany_top_out_144_[0]),
		.chany_top_out_146_(sb_0__1__0_chany_top_out_146_[0]),
		.chany_top_out_148_(sb_0__1__0_chany_top_out_148_[0]),
		.chany_top_out_150_(sb_0__1__0_chany_top_out_150_[0]),
		.chany_top_out_152_(sb_0__1__0_chany_top_out_152_[0]),
		.chany_top_out_154_(sb_0__1__0_chany_top_out_154_[0]),
		.chany_top_out_156_(sb_0__1__0_chany_top_out_156_[0]),
		.chany_top_out_158_(sb_0__1__0_chany_top_out_158_[0]),
		.chany_top_out_160_(sb_0__1__0_chany_top_out_160_[0]),
		.chany_top_out_162_(sb_0__1__0_chany_top_out_162_[0]),
		.chany_top_out_164_(sb_0__1__0_chany_top_out_164_[0]),
		.chany_top_out_166_(sb_0__1__0_chany_top_out_166_[0]),
		.chany_top_out_168_(sb_0__1__0_chany_top_out_168_[0]),
		.chany_top_out_170_(sb_0__1__0_chany_top_out_170_[0]),
		.chany_top_out_172_(sb_0__1__0_chany_top_out_172_[0]),
		.chany_top_out_174_(sb_0__1__0_chany_top_out_174_[0]),
		.chany_top_out_176_(sb_0__1__0_chany_top_out_176_[0]),
		.chany_top_out_178_(sb_0__1__0_chany_top_out_178_[0]),
		.chany_top_out_180_(sb_0__1__0_chany_top_out_180_[0]),
		.chany_top_out_182_(sb_0__1__0_chany_top_out_182_[0]),
		.chany_top_out_184_(sb_0__1__0_chany_top_out_184_[0]),
		.chany_top_out_186_(sb_0__1__0_chany_top_out_186_[0]),
		.chany_top_out_188_(sb_0__1__0_chany_top_out_188_[0]),
		.chany_top_out_190_(sb_0__1__0_chany_top_out_190_[0]),
		.chany_top_out_192_(sb_0__1__0_chany_top_out_192_[0]),
		.chany_top_out_194_(sb_0__1__0_chany_top_out_194_[0]),
		.chany_top_out_196_(sb_0__1__0_chany_top_out_196_[0]),
		.chany_top_out_198_(sb_0__1__0_chany_top_out_198_[0]),
		.chanx_right_out_0_(sb_0__1__0_chanx_right_out_0_[0]),
		.chanx_right_out_2_(sb_0__1__0_chanx_right_out_2_[0]),
		.chanx_right_out_4_(sb_0__1__0_chanx_right_out_4_[0]),
		.chanx_right_out_6_(sb_0__1__0_chanx_right_out_6_[0]),
		.chanx_right_out_8_(sb_0__1__0_chanx_right_out_8_[0]),
		.chanx_right_out_10_(sb_0__1__0_chanx_right_out_10_[0]),
		.chanx_right_out_12_(sb_0__1__0_chanx_right_out_12_[0]),
		.chanx_right_out_14_(sb_0__1__0_chanx_right_out_14_[0]),
		.chanx_right_out_16_(sb_0__1__0_chanx_right_out_16_[0]),
		.chanx_right_out_18_(sb_0__1__0_chanx_right_out_18_[0]),
		.chanx_right_out_20_(sb_0__1__0_chanx_right_out_20_[0]),
		.chanx_right_out_22_(sb_0__1__0_chanx_right_out_22_[0]),
		.chanx_right_out_24_(sb_0__1__0_chanx_right_out_24_[0]),
		.chanx_right_out_26_(sb_0__1__0_chanx_right_out_26_[0]),
		.chanx_right_out_28_(sb_0__1__0_chanx_right_out_28_[0]),
		.chanx_right_out_30_(sb_0__1__0_chanx_right_out_30_[0]),
		.chanx_right_out_32_(sb_0__1__0_chanx_right_out_32_[0]),
		.chanx_right_out_34_(sb_0__1__0_chanx_right_out_34_[0]),
		.chanx_right_out_36_(sb_0__1__0_chanx_right_out_36_[0]),
		.chanx_right_out_38_(sb_0__1__0_chanx_right_out_38_[0]),
		.chanx_right_out_40_(sb_0__1__0_chanx_right_out_40_[0]),
		.chanx_right_out_42_(sb_0__1__0_chanx_right_out_42_[0]),
		.chanx_right_out_44_(sb_0__1__0_chanx_right_out_44_[0]),
		.chanx_right_out_46_(sb_0__1__0_chanx_right_out_46_[0]),
		.chanx_right_out_48_(sb_0__1__0_chanx_right_out_48_[0]),
		.chanx_right_out_50_(sb_0__1__0_chanx_right_out_50_[0]),
		.chanx_right_out_52_(sb_0__1__0_chanx_right_out_52_[0]),
		.chanx_right_out_54_(sb_0__1__0_chanx_right_out_54_[0]),
		.chanx_right_out_56_(sb_0__1__0_chanx_right_out_56_[0]),
		.chanx_right_out_58_(sb_0__1__0_chanx_right_out_58_[0]),
		.chanx_right_out_60_(sb_0__1__0_chanx_right_out_60_[0]),
		.chanx_right_out_62_(sb_0__1__0_chanx_right_out_62_[0]),
		.chanx_right_out_64_(sb_0__1__0_chanx_right_out_64_[0]),
		.chanx_right_out_66_(sb_0__1__0_chanx_right_out_66_[0]),
		.chanx_right_out_68_(sb_0__1__0_chanx_right_out_68_[0]),
		.chanx_right_out_70_(sb_0__1__0_chanx_right_out_70_[0]),
		.chanx_right_out_72_(sb_0__1__0_chanx_right_out_72_[0]),
		.chanx_right_out_74_(sb_0__1__0_chanx_right_out_74_[0]),
		.chanx_right_out_76_(sb_0__1__0_chanx_right_out_76_[0]),
		.chanx_right_out_78_(sb_0__1__0_chanx_right_out_78_[0]),
		.chanx_right_out_80_(sb_0__1__0_chanx_right_out_80_[0]),
		.chanx_right_out_82_(sb_0__1__0_chanx_right_out_82_[0]),
		.chanx_right_out_84_(sb_0__1__0_chanx_right_out_84_[0]),
		.chanx_right_out_86_(sb_0__1__0_chanx_right_out_86_[0]),
		.chanx_right_out_88_(sb_0__1__0_chanx_right_out_88_[0]),
		.chanx_right_out_90_(sb_0__1__0_chanx_right_out_90_[0]),
		.chanx_right_out_92_(sb_0__1__0_chanx_right_out_92_[0]),
		.chanx_right_out_94_(sb_0__1__0_chanx_right_out_94_[0]),
		.chanx_right_out_96_(sb_0__1__0_chanx_right_out_96_[0]),
		.chanx_right_out_98_(sb_0__1__0_chanx_right_out_98_[0]),
		.chanx_right_out_100_(sb_0__1__0_chanx_right_out_100_[0]),
		.chanx_right_out_102_(sb_0__1__0_chanx_right_out_102_[0]),
		.chanx_right_out_104_(sb_0__1__0_chanx_right_out_104_[0]),
		.chanx_right_out_106_(sb_0__1__0_chanx_right_out_106_[0]),
		.chanx_right_out_108_(sb_0__1__0_chanx_right_out_108_[0]),
		.chanx_right_out_110_(sb_0__1__0_chanx_right_out_110_[0]),
		.chanx_right_out_112_(sb_0__1__0_chanx_right_out_112_[0]),
		.chanx_right_out_114_(sb_0__1__0_chanx_right_out_114_[0]),
		.chanx_right_out_116_(sb_0__1__0_chanx_right_out_116_[0]),
		.chanx_right_out_118_(sb_0__1__0_chanx_right_out_118_[0]),
		.chanx_right_out_120_(sb_0__1__0_chanx_right_out_120_[0]),
		.chanx_right_out_122_(sb_0__1__0_chanx_right_out_122_[0]),
		.chanx_right_out_124_(sb_0__1__0_chanx_right_out_124_[0]),
		.chanx_right_out_126_(sb_0__1__0_chanx_right_out_126_[0]),
		.chanx_right_out_128_(sb_0__1__0_chanx_right_out_128_[0]),
		.chanx_right_out_130_(sb_0__1__0_chanx_right_out_130_[0]),
		.chanx_right_out_132_(sb_0__1__0_chanx_right_out_132_[0]),
		.chanx_right_out_134_(sb_0__1__0_chanx_right_out_134_[0]),
		.chanx_right_out_136_(sb_0__1__0_chanx_right_out_136_[0]),
		.chanx_right_out_138_(sb_0__1__0_chanx_right_out_138_[0]),
		.chanx_right_out_140_(sb_0__1__0_chanx_right_out_140_[0]),
		.chanx_right_out_142_(sb_0__1__0_chanx_right_out_142_[0]),
		.chanx_right_out_144_(sb_0__1__0_chanx_right_out_144_[0]),
		.chanx_right_out_146_(sb_0__1__0_chanx_right_out_146_[0]),
		.chanx_right_out_148_(sb_0__1__0_chanx_right_out_148_[0]),
		.chanx_right_out_150_(sb_0__1__0_chanx_right_out_150_[0]),
		.chanx_right_out_152_(sb_0__1__0_chanx_right_out_152_[0]),
		.chanx_right_out_154_(sb_0__1__0_chanx_right_out_154_[0]),
		.chanx_right_out_156_(sb_0__1__0_chanx_right_out_156_[0]),
		.chanx_right_out_158_(sb_0__1__0_chanx_right_out_158_[0]),
		.chanx_right_out_160_(sb_0__1__0_chanx_right_out_160_[0]),
		.chanx_right_out_162_(sb_0__1__0_chanx_right_out_162_[0]),
		.chanx_right_out_164_(sb_0__1__0_chanx_right_out_164_[0]),
		.chanx_right_out_166_(sb_0__1__0_chanx_right_out_166_[0]),
		.chanx_right_out_168_(sb_0__1__0_chanx_right_out_168_[0]),
		.chanx_right_out_170_(sb_0__1__0_chanx_right_out_170_[0]),
		.chanx_right_out_172_(sb_0__1__0_chanx_right_out_172_[0]),
		.chanx_right_out_174_(sb_0__1__0_chanx_right_out_174_[0]),
		.chanx_right_out_176_(sb_0__1__0_chanx_right_out_176_[0]),
		.chanx_right_out_178_(sb_0__1__0_chanx_right_out_178_[0]),
		.chanx_right_out_180_(sb_0__1__0_chanx_right_out_180_[0]),
		.chanx_right_out_182_(sb_0__1__0_chanx_right_out_182_[0]),
		.chanx_right_out_184_(sb_0__1__0_chanx_right_out_184_[0]),
		.chanx_right_out_186_(sb_0__1__0_chanx_right_out_186_[0]),
		.chanx_right_out_188_(sb_0__1__0_chanx_right_out_188_[0]),
		.chanx_right_out_190_(sb_0__1__0_chanx_right_out_190_[0]),
		.chanx_right_out_192_(sb_0__1__0_chanx_right_out_192_[0]),
		.chanx_right_out_194_(sb_0__1__0_chanx_right_out_194_[0]),
		.chanx_right_out_196_(sb_0__1__0_chanx_right_out_196_[0]),
		.chanx_right_out_198_(sb_0__1__0_chanx_right_out_198_[0]),
		.chany_bottom_out_1_(sb_0__1__0_chany_bottom_out_1_[0]),
		.chany_bottom_out_3_(sb_0__1__0_chany_bottom_out_3_[0]),
		.chany_bottom_out_5_(sb_0__1__0_chany_bottom_out_5_[0]),
		.chany_bottom_out_7_(sb_0__1__0_chany_bottom_out_7_[0]),
		.chany_bottom_out_9_(sb_0__1__0_chany_bottom_out_9_[0]),
		.chany_bottom_out_11_(sb_0__1__0_chany_bottom_out_11_[0]),
		.chany_bottom_out_13_(sb_0__1__0_chany_bottom_out_13_[0]),
		.chany_bottom_out_15_(sb_0__1__0_chany_bottom_out_15_[0]),
		.chany_bottom_out_17_(sb_0__1__0_chany_bottom_out_17_[0]),
		.chany_bottom_out_19_(sb_0__1__0_chany_bottom_out_19_[0]),
		.chany_bottom_out_21_(sb_0__1__0_chany_bottom_out_21_[0]),
		.chany_bottom_out_23_(sb_0__1__0_chany_bottom_out_23_[0]),
		.chany_bottom_out_25_(sb_0__1__0_chany_bottom_out_25_[0]),
		.chany_bottom_out_27_(sb_0__1__0_chany_bottom_out_27_[0]),
		.chany_bottom_out_29_(sb_0__1__0_chany_bottom_out_29_[0]),
		.chany_bottom_out_31_(sb_0__1__0_chany_bottom_out_31_[0]),
		.chany_bottom_out_33_(sb_0__1__0_chany_bottom_out_33_[0]),
		.chany_bottom_out_35_(sb_0__1__0_chany_bottom_out_35_[0]),
		.chany_bottom_out_37_(sb_0__1__0_chany_bottom_out_37_[0]),
		.chany_bottom_out_39_(sb_0__1__0_chany_bottom_out_39_[0]),
		.chany_bottom_out_41_(sb_0__1__0_chany_bottom_out_41_[0]),
		.chany_bottom_out_43_(sb_0__1__0_chany_bottom_out_43_[0]),
		.chany_bottom_out_45_(sb_0__1__0_chany_bottom_out_45_[0]),
		.chany_bottom_out_47_(sb_0__1__0_chany_bottom_out_47_[0]),
		.chany_bottom_out_49_(sb_0__1__0_chany_bottom_out_49_[0]),
		.chany_bottom_out_51_(sb_0__1__0_chany_bottom_out_51_[0]),
		.chany_bottom_out_53_(sb_0__1__0_chany_bottom_out_53_[0]),
		.chany_bottom_out_55_(sb_0__1__0_chany_bottom_out_55_[0]),
		.chany_bottom_out_57_(sb_0__1__0_chany_bottom_out_57_[0]),
		.chany_bottom_out_59_(sb_0__1__0_chany_bottom_out_59_[0]),
		.chany_bottom_out_61_(sb_0__1__0_chany_bottom_out_61_[0]),
		.chany_bottom_out_63_(sb_0__1__0_chany_bottom_out_63_[0]),
		.chany_bottom_out_65_(sb_0__1__0_chany_bottom_out_65_[0]),
		.chany_bottom_out_67_(sb_0__1__0_chany_bottom_out_67_[0]),
		.chany_bottom_out_69_(sb_0__1__0_chany_bottom_out_69_[0]),
		.chany_bottom_out_71_(sb_0__1__0_chany_bottom_out_71_[0]),
		.chany_bottom_out_73_(sb_0__1__0_chany_bottom_out_73_[0]),
		.chany_bottom_out_75_(sb_0__1__0_chany_bottom_out_75_[0]),
		.chany_bottom_out_77_(sb_0__1__0_chany_bottom_out_77_[0]),
		.chany_bottom_out_79_(sb_0__1__0_chany_bottom_out_79_[0]),
		.chany_bottom_out_81_(sb_0__1__0_chany_bottom_out_81_[0]),
		.chany_bottom_out_83_(sb_0__1__0_chany_bottom_out_83_[0]),
		.chany_bottom_out_85_(sb_0__1__0_chany_bottom_out_85_[0]),
		.chany_bottom_out_87_(sb_0__1__0_chany_bottom_out_87_[0]),
		.chany_bottom_out_89_(sb_0__1__0_chany_bottom_out_89_[0]),
		.chany_bottom_out_91_(sb_0__1__0_chany_bottom_out_91_[0]),
		.chany_bottom_out_93_(sb_0__1__0_chany_bottom_out_93_[0]),
		.chany_bottom_out_95_(sb_0__1__0_chany_bottom_out_95_[0]),
		.chany_bottom_out_97_(sb_0__1__0_chany_bottom_out_97_[0]),
		.chany_bottom_out_99_(sb_0__1__0_chany_bottom_out_99_[0]),
		.chany_bottom_out_101_(sb_0__1__0_chany_bottom_out_101_[0]),
		.chany_bottom_out_103_(sb_0__1__0_chany_bottom_out_103_[0]),
		.chany_bottom_out_105_(sb_0__1__0_chany_bottom_out_105_[0]),
		.chany_bottom_out_107_(sb_0__1__0_chany_bottom_out_107_[0]),
		.chany_bottom_out_109_(sb_0__1__0_chany_bottom_out_109_[0]),
		.chany_bottom_out_111_(sb_0__1__0_chany_bottom_out_111_[0]),
		.chany_bottom_out_113_(sb_0__1__0_chany_bottom_out_113_[0]),
		.chany_bottom_out_115_(sb_0__1__0_chany_bottom_out_115_[0]),
		.chany_bottom_out_117_(sb_0__1__0_chany_bottom_out_117_[0]),
		.chany_bottom_out_119_(sb_0__1__0_chany_bottom_out_119_[0]),
		.chany_bottom_out_121_(sb_0__1__0_chany_bottom_out_121_[0]),
		.chany_bottom_out_123_(sb_0__1__0_chany_bottom_out_123_[0]),
		.chany_bottom_out_125_(sb_0__1__0_chany_bottom_out_125_[0]),
		.chany_bottom_out_127_(sb_0__1__0_chany_bottom_out_127_[0]),
		.chany_bottom_out_129_(sb_0__1__0_chany_bottom_out_129_[0]),
		.chany_bottom_out_131_(sb_0__1__0_chany_bottom_out_131_[0]),
		.chany_bottom_out_133_(sb_0__1__0_chany_bottom_out_133_[0]),
		.chany_bottom_out_135_(sb_0__1__0_chany_bottom_out_135_[0]),
		.chany_bottom_out_137_(sb_0__1__0_chany_bottom_out_137_[0]),
		.chany_bottom_out_139_(sb_0__1__0_chany_bottom_out_139_[0]),
		.chany_bottom_out_141_(sb_0__1__0_chany_bottom_out_141_[0]),
		.chany_bottom_out_143_(sb_0__1__0_chany_bottom_out_143_[0]),
		.chany_bottom_out_145_(sb_0__1__0_chany_bottom_out_145_[0]),
		.chany_bottom_out_147_(sb_0__1__0_chany_bottom_out_147_[0]),
		.chany_bottom_out_149_(sb_0__1__0_chany_bottom_out_149_[0]),
		.chany_bottom_out_151_(sb_0__1__0_chany_bottom_out_151_[0]),
		.chany_bottom_out_153_(sb_0__1__0_chany_bottom_out_153_[0]),
		.chany_bottom_out_155_(sb_0__1__0_chany_bottom_out_155_[0]),
		.chany_bottom_out_157_(sb_0__1__0_chany_bottom_out_157_[0]),
		.chany_bottom_out_159_(sb_0__1__0_chany_bottom_out_159_[0]),
		.chany_bottom_out_161_(sb_0__1__0_chany_bottom_out_161_[0]),
		.chany_bottom_out_163_(sb_0__1__0_chany_bottom_out_163_[0]),
		.chany_bottom_out_165_(sb_0__1__0_chany_bottom_out_165_[0]),
		.chany_bottom_out_167_(sb_0__1__0_chany_bottom_out_167_[0]),
		.chany_bottom_out_169_(sb_0__1__0_chany_bottom_out_169_[0]),
		.chany_bottom_out_171_(sb_0__1__0_chany_bottom_out_171_[0]),
		.chany_bottom_out_173_(sb_0__1__0_chany_bottom_out_173_[0]),
		.chany_bottom_out_175_(sb_0__1__0_chany_bottom_out_175_[0]),
		.chany_bottom_out_177_(sb_0__1__0_chany_bottom_out_177_[0]),
		.chany_bottom_out_179_(sb_0__1__0_chany_bottom_out_179_[0]),
		.chany_bottom_out_181_(sb_0__1__0_chany_bottom_out_181_[0]),
		.chany_bottom_out_183_(sb_0__1__0_chany_bottom_out_183_[0]),
		.chany_bottom_out_185_(sb_0__1__0_chany_bottom_out_185_[0]),
		.chany_bottom_out_187_(sb_0__1__0_chany_bottom_out_187_[0]),
		.chany_bottom_out_189_(sb_0__1__0_chany_bottom_out_189_[0]),
		.chany_bottom_out_191_(sb_0__1__0_chany_bottom_out_191_[0]),
		.chany_bottom_out_193_(sb_0__1__0_chany_bottom_out_193_[0]),
		.chany_bottom_out_195_(sb_0__1__0_chany_bottom_out_195_[0]),
		.chany_bottom_out_197_(sb_0__1__0_chany_bottom_out_197_[0]),
		.chany_bottom_out_199_(sb_0__1__0_chany_bottom_out_199_[0]),
		.ccff_tail(sb_0__1__0_ccff_tail[0]));

	sb_0__2_ sb_0__2_ (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.chanx_right_in_1_(cbx_1__2__0_chanx_out_1_[0]),
		.chanx_right_in_3_(cbx_1__2__0_chanx_out_3_[0]),
		.chanx_right_in_5_(cbx_1__2__0_chanx_out_5_[0]),
		.chanx_right_in_7_(cbx_1__2__0_chanx_out_7_[0]),
		.chanx_right_in_9_(cbx_1__2__0_chanx_out_9_[0]),
		.chanx_right_in_11_(cbx_1__2__0_chanx_out_11_[0]),
		.chanx_right_in_13_(cbx_1__2__0_chanx_out_13_[0]),
		.chanx_right_in_15_(cbx_1__2__0_chanx_out_15_[0]),
		.chanx_right_in_17_(cbx_1__2__0_chanx_out_17_[0]),
		.chanx_right_in_19_(cbx_1__2__0_chanx_out_19_[0]),
		.chanx_right_in_21_(cbx_1__2__0_chanx_out_21_[0]),
		.chanx_right_in_23_(cbx_1__2__0_chanx_out_23_[0]),
		.chanx_right_in_25_(cbx_1__2__0_chanx_out_25_[0]),
		.chanx_right_in_27_(cbx_1__2__0_chanx_out_27_[0]),
		.chanx_right_in_29_(cbx_1__2__0_chanx_out_29_[0]),
		.chanx_right_in_31_(cbx_1__2__0_chanx_out_31_[0]),
		.chanx_right_in_33_(cbx_1__2__0_chanx_out_33_[0]),
		.chanx_right_in_35_(cbx_1__2__0_chanx_out_35_[0]),
		.chanx_right_in_37_(cbx_1__2__0_chanx_out_37_[0]),
		.chanx_right_in_39_(cbx_1__2__0_chanx_out_39_[0]),
		.chanx_right_in_41_(cbx_1__2__0_chanx_out_41_[0]),
		.chanx_right_in_43_(cbx_1__2__0_chanx_out_43_[0]),
		.chanx_right_in_45_(cbx_1__2__0_chanx_out_45_[0]),
		.chanx_right_in_47_(cbx_1__2__0_chanx_out_47_[0]),
		.chanx_right_in_49_(cbx_1__2__0_chanx_out_49_[0]),
		.chanx_right_in_51_(cbx_1__2__0_chanx_out_51_[0]),
		.chanx_right_in_53_(cbx_1__2__0_chanx_out_53_[0]),
		.chanx_right_in_55_(cbx_1__2__0_chanx_out_55_[0]),
		.chanx_right_in_57_(cbx_1__2__0_chanx_out_57_[0]),
		.chanx_right_in_59_(cbx_1__2__0_chanx_out_59_[0]),
		.chanx_right_in_61_(cbx_1__2__0_chanx_out_61_[0]),
		.chanx_right_in_63_(cbx_1__2__0_chanx_out_63_[0]),
		.chanx_right_in_65_(cbx_1__2__0_chanx_out_65_[0]),
		.chanx_right_in_67_(cbx_1__2__0_chanx_out_67_[0]),
		.chanx_right_in_69_(cbx_1__2__0_chanx_out_69_[0]),
		.chanx_right_in_71_(cbx_1__2__0_chanx_out_71_[0]),
		.chanx_right_in_73_(cbx_1__2__0_chanx_out_73_[0]),
		.chanx_right_in_75_(cbx_1__2__0_chanx_out_75_[0]),
		.chanx_right_in_77_(cbx_1__2__0_chanx_out_77_[0]),
		.chanx_right_in_79_(cbx_1__2__0_chanx_out_79_[0]),
		.chanx_right_in_81_(cbx_1__2__0_chanx_out_81_[0]),
		.chanx_right_in_83_(cbx_1__2__0_chanx_out_83_[0]),
		.chanx_right_in_85_(cbx_1__2__0_chanx_out_85_[0]),
		.chanx_right_in_87_(cbx_1__2__0_chanx_out_87_[0]),
		.chanx_right_in_89_(cbx_1__2__0_chanx_out_89_[0]),
		.chanx_right_in_91_(cbx_1__2__0_chanx_out_91_[0]),
		.chanx_right_in_93_(cbx_1__2__0_chanx_out_93_[0]),
		.chanx_right_in_95_(cbx_1__2__0_chanx_out_95_[0]),
		.chanx_right_in_97_(cbx_1__2__0_chanx_out_97_[0]),
		.chanx_right_in_99_(cbx_1__2__0_chanx_out_99_[0]),
		.chanx_right_in_101_(cbx_1__2__0_chanx_out_101_[0]),
		.chanx_right_in_103_(cbx_1__2__0_chanx_out_103_[0]),
		.chanx_right_in_105_(cbx_1__2__0_chanx_out_105_[0]),
		.chanx_right_in_107_(cbx_1__2__0_chanx_out_107_[0]),
		.chanx_right_in_109_(cbx_1__2__0_chanx_out_109_[0]),
		.chanx_right_in_111_(cbx_1__2__0_chanx_out_111_[0]),
		.chanx_right_in_113_(cbx_1__2__0_chanx_out_113_[0]),
		.chanx_right_in_115_(cbx_1__2__0_chanx_out_115_[0]),
		.chanx_right_in_117_(cbx_1__2__0_chanx_out_117_[0]),
		.chanx_right_in_119_(cbx_1__2__0_chanx_out_119_[0]),
		.chanx_right_in_121_(cbx_1__2__0_chanx_out_121_[0]),
		.chanx_right_in_123_(cbx_1__2__0_chanx_out_123_[0]),
		.chanx_right_in_125_(cbx_1__2__0_chanx_out_125_[0]),
		.chanx_right_in_127_(cbx_1__2__0_chanx_out_127_[0]),
		.chanx_right_in_129_(cbx_1__2__0_chanx_out_129_[0]),
		.chanx_right_in_131_(cbx_1__2__0_chanx_out_131_[0]),
		.chanx_right_in_133_(cbx_1__2__0_chanx_out_133_[0]),
		.chanx_right_in_135_(cbx_1__2__0_chanx_out_135_[0]),
		.chanx_right_in_137_(cbx_1__2__0_chanx_out_137_[0]),
		.chanx_right_in_139_(cbx_1__2__0_chanx_out_139_[0]),
		.chanx_right_in_141_(cbx_1__2__0_chanx_out_141_[0]),
		.chanx_right_in_143_(cbx_1__2__0_chanx_out_143_[0]),
		.chanx_right_in_145_(cbx_1__2__0_chanx_out_145_[0]),
		.chanx_right_in_147_(cbx_1__2__0_chanx_out_147_[0]),
		.chanx_right_in_149_(cbx_1__2__0_chanx_out_149_[0]),
		.chanx_right_in_151_(cbx_1__2__0_chanx_out_151_[0]),
		.chanx_right_in_153_(cbx_1__2__0_chanx_out_153_[0]),
		.chanx_right_in_155_(cbx_1__2__0_chanx_out_155_[0]),
		.chanx_right_in_157_(cbx_1__2__0_chanx_out_157_[0]),
		.chanx_right_in_159_(cbx_1__2__0_chanx_out_159_[0]),
		.chanx_right_in_161_(cbx_1__2__0_chanx_out_161_[0]),
		.chanx_right_in_163_(cbx_1__2__0_chanx_out_163_[0]),
		.chanx_right_in_165_(cbx_1__2__0_chanx_out_165_[0]),
		.chanx_right_in_167_(cbx_1__2__0_chanx_out_167_[0]),
		.chanx_right_in_169_(cbx_1__2__0_chanx_out_169_[0]),
		.chanx_right_in_171_(cbx_1__2__0_chanx_out_171_[0]),
		.chanx_right_in_173_(cbx_1__2__0_chanx_out_173_[0]),
		.chanx_right_in_175_(cbx_1__2__0_chanx_out_175_[0]),
		.chanx_right_in_177_(cbx_1__2__0_chanx_out_177_[0]),
		.chanx_right_in_179_(cbx_1__2__0_chanx_out_179_[0]),
		.chanx_right_in_181_(cbx_1__2__0_chanx_out_181_[0]),
		.chanx_right_in_183_(cbx_1__2__0_chanx_out_183_[0]),
		.chanx_right_in_185_(cbx_1__2__0_chanx_out_185_[0]),
		.chanx_right_in_187_(cbx_1__2__0_chanx_out_187_[0]),
		.chanx_right_in_189_(cbx_1__2__0_chanx_out_189_[0]),
		.chanx_right_in_191_(cbx_1__2__0_chanx_out_191_[0]),
		.chanx_right_in_193_(cbx_1__2__0_chanx_out_193_[0]),
		.chanx_right_in_195_(cbx_1__2__0_chanx_out_195_[0]),
		.chanx_right_in_197_(cbx_1__2__0_chanx_out_197_[0]),
		.chanx_right_in_199_(cbx_1__2__0_chanx_out_199_[0]),
		.right_top_grid_pin_1_(grid_io_top_0_bottom_width_0_height_0__pin_1_upper[0]),
		.chany_bottom_in_0_(cby_0__1__1_chany_out_0_[0]),
		.chany_bottom_in_2_(cby_0__1__1_chany_out_2_[0]),
		.chany_bottom_in_4_(cby_0__1__1_chany_out_4_[0]),
		.chany_bottom_in_6_(cby_0__1__1_chany_out_6_[0]),
		.chany_bottom_in_8_(cby_0__1__1_chany_out_8_[0]),
		.chany_bottom_in_10_(cby_0__1__1_chany_out_10_[0]),
		.chany_bottom_in_12_(cby_0__1__1_chany_out_12_[0]),
		.chany_bottom_in_14_(cby_0__1__1_chany_out_14_[0]),
		.chany_bottom_in_16_(cby_0__1__1_chany_out_16_[0]),
		.chany_bottom_in_18_(cby_0__1__1_chany_out_18_[0]),
		.chany_bottom_in_20_(cby_0__1__1_chany_out_20_[0]),
		.chany_bottom_in_22_(cby_0__1__1_chany_out_22_[0]),
		.chany_bottom_in_24_(cby_0__1__1_chany_out_24_[0]),
		.chany_bottom_in_26_(cby_0__1__1_chany_out_26_[0]),
		.chany_bottom_in_28_(cby_0__1__1_chany_out_28_[0]),
		.chany_bottom_in_30_(cby_0__1__1_chany_out_30_[0]),
		.chany_bottom_in_32_(cby_0__1__1_chany_out_32_[0]),
		.chany_bottom_in_34_(cby_0__1__1_chany_out_34_[0]),
		.chany_bottom_in_36_(cby_0__1__1_chany_out_36_[0]),
		.chany_bottom_in_38_(cby_0__1__1_chany_out_38_[0]),
		.chany_bottom_in_40_(cby_0__1__1_chany_out_40_[0]),
		.chany_bottom_in_42_(cby_0__1__1_chany_out_42_[0]),
		.chany_bottom_in_44_(cby_0__1__1_chany_out_44_[0]),
		.chany_bottom_in_46_(cby_0__1__1_chany_out_46_[0]),
		.chany_bottom_in_48_(cby_0__1__1_chany_out_48_[0]),
		.chany_bottom_in_50_(cby_0__1__1_chany_out_50_[0]),
		.chany_bottom_in_52_(cby_0__1__1_chany_out_52_[0]),
		.chany_bottom_in_54_(cby_0__1__1_chany_out_54_[0]),
		.chany_bottom_in_56_(cby_0__1__1_chany_out_56_[0]),
		.chany_bottom_in_58_(cby_0__1__1_chany_out_58_[0]),
		.chany_bottom_in_60_(cby_0__1__1_chany_out_60_[0]),
		.chany_bottom_in_62_(cby_0__1__1_chany_out_62_[0]),
		.chany_bottom_in_64_(cby_0__1__1_chany_out_64_[0]),
		.chany_bottom_in_66_(cby_0__1__1_chany_out_66_[0]),
		.chany_bottom_in_68_(cby_0__1__1_chany_out_68_[0]),
		.chany_bottom_in_70_(cby_0__1__1_chany_out_70_[0]),
		.chany_bottom_in_72_(cby_0__1__1_chany_out_72_[0]),
		.chany_bottom_in_74_(cby_0__1__1_chany_out_74_[0]),
		.chany_bottom_in_76_(cby_0__1__1_chany_out_76_[0]),
		.chany_bottom_in_78_(cby_0__1__1_chany_out_78_[0]),
		.chany_bottom_in_80_(cby_0__1__1_chany_out_80_[0]),
		.chany_bottom_in_82_(cby_0__1__1_chany_out_82_[0]),
		.chany_bottom_in_84_(cby_0__1__1_chany_out_84_[0]),
		.chany_bottom_in_86_(cby_0__1__1_chany_out_86_[0]),
		.chany_bottom_in_88_(cby_0__1__1_chany_out_88_[0]),
		.chany_bottom_in_90_(cby_0__1__1_chany_out_90_[0]),
		.chany_bottom_in_92_(cby_0__1__1_chany_out_92_[0]),
		.chany_bottom_in_94_(cby_0__1__1_chany_out_94_[0]),
		.chany_bottom_in_96_(cby_0__1__1_chany_out_96_[0]),
		.chany_bottom_in_98_(cby_0__1__1_chany_out_98_[0]),
		.chany_bottom_in_100_(cby_0__1__1_chany_out_100_[0]),
		.chany_bottom_in_102_(cby_0__1__1_chany_out_102_[0]),
		.chany_bottom_in_104_(cby_0__1__1_chany_out_104_[0]),
		.chany_bottom_in_106_(cby_0__1__1_chany_out_106_[0]),
		.chany_bottom_in_108_(cby_0__1__1_chany_out_108_[0]),
		.chany_bottom_in_110_(cby_0__1__1_chany_out_110_[0]),
		.chany_bottom_in_112_(cby_0__1__1_chany_out_112_[0]),
		.chany_bottom_in_114_(cby_0__1__1_chany_out_114_[0]),
		.chany_bottom_in_116_(cby_0__1__1_chany_out_116_[0]),
		.chany_bottom_in_118_(cby_0__1__1_chany_out_118_[0]),
		.chany_bottom_in_120_(cby_0__1__1_chany_out_120_[0]),
		.chany_bottom_in_122_(cby_0__1__1_chany_out_122_[0]),
		.chany_bottom_in_124_(cby_0__1__1_chany_out_124_[0]),
		.chany_bottom_in_126_(cby_0__1__1_chany_out_126_[0]),
		.chany_bottom_in_128_(cby_0__1__1_chany_out_128_[0]),
		.chany_bottom_in_130_(cby_0__1__1_chany_out_130_[0]),
		.chany_bottom_in_132_(cby_0__1__1_chany_out_132_[0]),
		.chany_bottom_in_134_(cby_0__1__1_chany_out_134_[0]),
		.chany_bottom_in_136_(cby_0__1__1_chany_out_136_[0]),
		.chany_bottom_in_138_(cby_0__1__1_chany_out_138_[0]),
		.chany_bottom_in_140_(cby_0__1__1_chany_out_140_[0]),
		.chany_bottom_in_142_(cby_0__1__1_chany_out_142_[0]),
		.chany_bottom_in_144_(cby_0__1__1_chany_out_144_[0]),
		.chany_bottom_in_146_(cby_0__1__1_chany_out_146_[0]),
		.chany_bottom_in_148_(cby_0__1__1_chany_out_148_[0]),
		.chany_bottom_in_150_(cby_0__1__1_chany_out_150_[0]),
		.chany_bottom_in_152_(cby_0__1__1_chany_out_152_[0]),
		.chany_bottom_in_154_(cby_0__1__1_chany_out_154_[0]),
		.chany_bottom_in_156_(cby_0__1__1_chany_out_156_[0]),
		.chany_bottom_in_158_(cby_0__1__1_chany_out_158_[0]),
		.chany_bottom_in_160_(cby_0__1__1_chany_out_160_[0]),
		.chany_bottom_in_162_(cby_0__1__1_chany_out_162_[0]),
		.chany_bottom_in_164_(cby_0__1__1_chany_out_164_[0]),
		.chany_bottom_in_166_(cby_0__1__1_chany_out_166_[0]),
		.chany_bottom_in_168_(cby_0__1__1_chany_out_168_[0]),
		.chany_bottom_in_170_(cby_0__1__1_chany_out_170_[0]),
		.chany_bottom_in_172_(cby_0__1__1_chany_out_172_[0]),
		.chany_bottom_in_174_(cby_0__1__1_chany_out_174_[0]),
		.chany_bottom_in_176_(cby_0__1__1_chany_out_176_[0]),
		.chany_bottom_in_178_(cby_0__1__1_chany_out_178_[0]),
		.chany_bottom_in_180_(cby_0__1__1_chany_out_180_[0]),
		.chany_bottom_in_182_(cby_0__1__1_chany_out_182_[0]),
		.chany_bottom_in_184_(cby_0__1__1_chany_out_184_[0]),
		.chany_bottom_in_186_(cby_0__1__1_chany_out_186_[0]),
		.chany_bottom_in_188_(cby_0__1__1_chany_out_188_[0]),
		.chany_bottom_in_190_(cby_0__1__1_chany_out_190_[0]),
		.chany_bottom_in_192_(cby_0__1__1_chany_out_192_[0]),
		.chany_bottom_in_194_(cby_0__1__1_chany_out_194_[0]),
		.chany_bottom_in_196_(cby_0__1__1_chany_out_196_[0]),
		.chany_bottom_in_198_(cby_0__1__1_chany_out_198_[0]),
		.bottom_left_grid_pin_1_(grid_io_left_1_right_width_0_height_0__pin_1_upper[0]),
		.ccff_head(grid_io_top_0_ccff_tail[0]),
		.chanx_right_out_0_(sb_0__2__0_chanx_right_out_0_[0]),
		.chanx_right_out_2_(sb_0__2__0_chanx_right_out_2_[0]),
		.chanx_right_out_4_(sb_0__2__0_chanx_right_out_4_[0]),
		.chanx_right_out_6_(sb_0__2__0_chanx_right_out_6_[0]),
		.chanx_right_out_8_(sb_0__2__0_chanx_right_out_8_[0]),
		.chanx_right_out_10_(sb_0__2__0_chanx_right_out_10_[0]),
		.chanx_right_out_12_(sb_0__2__0_chanx_right_out_12_[0]),
		.chanx_right_out_14_(sb_0__2__0_chanx_right_out_14_[0]),
		.chanx_right_out_16_(sb_0__2__0_chanx_right_out_16_[0]),
		.chanx_right_out_18_(sb_0__2__0_chanx_right_out_18_[0]),
		.chanx_right_out_20_(sb_0__2__0_chanx_right_out_20_[0]),
		.chanx_right_out_22_(sb_0__2__0_chanx_right_out_22_[0]),
		.chanx_right_out_24_(sb_0__2__0_chanx_right_out_24_[0]),
		.chanx_right_out_26_(sb_0__2__0_chanx_right_out_26_[0]),
		.chanx_right_out_28_(sb_0__2__0_chanx_right_out_28_[0]),
		.chanx_right_out_30_(sb_0__2__0_chanx_right_out_30_[0]),
		.chanx_right_out_32_(sb_0__2__0_chanx_right_out_32_[0]),
		.chanx_right_out_34_(sb_0__2__0_chanx_right_out_34_[0]),
		.chanx_right_out_36_(sb_0__2__0_chanx_right_out_36_[0]),
		.chanx_right_out_38_(sb_0__2__0_chanx_right_out_38_[0]),
		.chanx_right_out_40_(sb_0__2__0_chanx_right_out_40_[0]),
		.chanx_right_out_42_(sb_0__2__0_chanx_right_out_42_[0]),
		.chanx_right_out_44_(sb_0__2__0_chanx_right_out_44_[0]),
		.chanx_right_out_46_(sb_0__2__0_chanx_right_out_46_[0]),
		.chanx_right_out_48_(sb_0__2__0_chanx_right_out_48_[0]),
		.chanx_right_out_50_(sb_0__2__0_chanx_right_out_50_[0]),
		.chanx_right_out_52_(sb_0__2__0_chanx_right_out_52_[0]),
		.chanx_right_out_54_(sb_0__2__0_chanx_right_out_54_[0]),
		.chanx_right_out_56_(sb_0__2__0_chanx_right_out_56_[0]),
		.chanx_right_out_58_(sb_0__2__0_chanx_right_out_58_[0]),
		.chanx_right_out_60_(sb_0__2__0_chanx_right_out_60_[0]),
		.chanx_right_out_62_(sb_0__2__0_chanx_right_out_62_[0]),
		.chanx_right_out_64_(sb_0__2__0_chanx_right_out_64_[0]),
		.chanx_right_out_66_(sb_0__2__0_chanx_right_out_66_[0]),
		.chanx_right_out_68_(sb_0__2__0_chanx_right_out_68_[0]),
		.chanx_right_out_70_(sb_0__2__0_chanx_right_out_70_[0]),
		.chanx_right_out_72_(sb_0__2__0_chanx_right_out_72_[0]),
		.chanx_right_out_74_(sb_0__2__0_chanx_right_out_74_[0]),
		.chanx_right_out_76_(sb_0__2__0_chanx_right_out_76_[0]),
		.chanx_right_out_78_(sb_0__2__0_chanx_right_out_78_[0]),
		.chanx_right_out_80_(sb_0__2__0_chanx_right_out_80_[0]),
		.chanx_right_out_82_(sb_0__2__0_chanx_right_out_82_[0]),
		.chanx_right_out_84_(sb_0__2__0_chanx_right_out_84_[0]),
		.chanx_right_out_86_(sb_0__2__0_chanx_right_out_86_[0]),
		.chanx_right_out_88_(sb_0__2__0_chanx_right_out_88_[0]),
		.chanx_right_out_90_(sb_0__2__0_chanx_right_out_90_[0]),
		.chanx_right_out_92_(sb_0__2__0_chanx_right_out_92_[0]),
		.chanx_right_out_94_(sb_0__2__0_chanx_right_out_94_[0]),
		.chanx_right_out_96_(sb_0__2__0_chanx_right_out_96_[0]),
		.chanx_right_out_98_(sb_0__2__0_chanx_right_out_98_[0]),
		.chanx_right_out_100_(sb_0__2__0_chanx_right_out_100_[0]),
		.chanx_right_out_102_(sb_0__2__0_chanx_right_out_102_[0]),
		.chanx_right_out_104_(sb_0__2__0_chanx_right_out_104_[0]),
		.chanx_right_out_106_(sb_0__2__0_chanx_right_out_106_[0]),
		.chanx_right_out_108_(sb_0__2__0_chanx_right_out_108_[0]),
		.chanx_right_out_110_(sb_0__2__0_chanx_right_out_110_[0]),
		.chanx_right_out_112_(sb_0__2__0_chanx_right_out_112_[0]),
		.chanx_right_out_114_(sb_0__2__0_chanx_right_out_114_[0]),
		.chanx_right_out_116_(sb_0__2__0_chanx_right_out_116_[0]),
		.chanx_right_out_118_(sb_0__2__0_chanx_right_out_118_[0]),
		.chanx_right_out_120_(sb_0__2__0_chanx_right_out_120_[0]),
		.chanx_right_out_122_(sb_0__2__0_chanx_right_out_122_[0]),
		.chanx_right_out_124_(sb_0__2__0_chanx_right_out_124_[0]),
		.chanx_right_out_126_(sb_0__2__0_chanx_right_out_126_[0]),
		.chanx_right_out_128_(sb_0__2__0_chanx_right_out_128_[0]),
		.chanx_right_out_130_(sb_0__2__0_chanx_right_out_130_[0]),
		.chanx_right_out_132_(sb_0__2__0_chanx_right_out_132_[0]),
		.chanx_right_out_134_(sb_0__2__0_chanx_right_out_134_[0]),
		.chanx_right_out_136_(sb_0__2__0_chanx_right_out_136_[0]),
		.chanx_right_out_138_(sb_0__2__0_chanx_right_out_138_[0]),
		.chanx_right_out_140_(sb_0__2__0_chanx_right_out_140_[0]),
		.chanx_right_out_142_(sb_0__2__0_chanx_right_out_142_[0]),
		.chanx_right_out_144_(sb_0__2__0_chanx_right_out_144_[0]),
		.chanx_right_out_146_(sb_0__2__0_chanx_right_out_146_[0]),
		.chanx_right_out_148_(sb_0__2__0_chanx_right_out_148_[0]),
		.chanx_right_out_150_(sb_0__2__0_chanx_right_out_150_[0]),
		.chanx_right_out_152_(sb_0__2__0_chanx_right_out_152_[0]),
		.chanx_right_out_154_(sb_0__2__0_chanx_right_out_154_[0]),
		.chanx_right_out_156_(sb_0__2__0_chanx_right_out_156_[0]),
		.chanx_right_out_158_(sb_0__2__0_chanx_right_out_158_[0]),
		.chanx_right_out_160_(sb_0__2__0_chanx_right_out_160_[0]),
		.chanx_right_out_162_(sb_0__2__0_chanx_right_out_162_[0]),
		.chanx_right_out_164_(sb_0__2__0_chanx_right_out_164_[0]),
		.chanx_right_out_166_(sb_0__2__0_chanx_right_out_166_[0]),
		.chanx_right_out_168_(sb_0__2__0_chanx_right_out_168_[0]),
		.chanx_right_out_170_(sb_0__2__0_chanx_right_out_170_[0]),
		.chanx_right_out_172_(sb_0__2__0_chanx_right_out_172_[0]),
		.chanx_right_out_174_(sb_0__2__0_chanx_right_out_174_[0]),
		.chanx_right_out_176_(sb_0__2__0_chanx_right_out_176_[0]),
		.chanx_right_out_178_(sb_0__2__0_chanx_right_out_178_[0]),
		.chanx_right_out_180_(sb_0__2__0_chanx_right_out_180_[0]),
		.chanx_right_out_182_(sb_0__2__0_chanx_right_out_182_[0]),
		.chanx_right_out_184_(sb_0__2__0_chanx_right_out_184_[0]),
		.chanx_right_out_186_(sb_0__2__0_chanx_right_out_186_[0]),
		.chanx_right_out_188_(sb_0__2__0_chanx_right_out_188_[0]),
		.chanx_right_out_190_(sb_0__2__0_chanx_right_out_190_[0]),
		.chanx_right_out_192_(sb_0__2__0_chanx_right_out_192_[0]),
		.chanx_right_out_194_(sb_0__2__0_chanx_right_out_194_[0]),
		.chanx_right_out_196_(sb_0__2__0_chanx_right_out_196_[0]),
		.chanx_right_out_198_(sb_0__2__0_chanx_right_out_198_[0]),
		.chany_bottom_out_1_(sb_0__2__0_chany_bottom_out_1_[0]),
		.chany_bottom_out_3_(sb_0__2__0_chany_bottom_out_3_[0]),
		.chany_bottom_out_5_(sb_0__2__0_chany_bottom_out_5_[0]),
		.chany_bottom_out_7_(sb_0__2__0_chany_bottom_out_7_[0]),
		.chany_bottom_out_9_(sb_0__2__0_chany_bottom_out_9_[0]),
		.chany_bottom_out_11_(sb_0__2__0_chany_bottom_out_11_[0]),
		.chany_bottom_out_13_(sb_0__2__0_chany_bottom_out_13_[0]),
		.chany_bottom_out_15_(sb_0__2__0_chany_bottom_out_15_[0]),
		.chany_bottom_out_17_(sb_0__2__0_chany_bottom_out_17_[0]),
		.chany_bottom_out_19_(sb_0__2__0_chany_bottom_out_19_[0]),
		.chany_bottom_out_21_(sb_0__2__0_chany_bottom_out_21_[0]),
		.chany_bottom_out_23_(sb_0__2__0_chany_bottom_out_23_[0]),
		.chany_bottom_out_25_(sb_0__2__0_chany_bottom_out_25_[0]),
		.chany_bottom_out_27_(sb_0__2__0_chany_bottom_out_27_[0]),
		.chany_bottom_out_29_(sb_0__2__0_chany_bottom_out_29_[0]),
		.chany_bottom_out_31_(sb_0__2__0_chany_bottom_out_31_[0]),
		.chany_bottom_out_33_(sb_0__2__0_chany_bottom_out_33_[0]),
		.chany_bottom_out_35_(sb_0__2__0_chany_bottom_out_35_[0]),
		.chany_bottom_out_37_(sb_0__2__0_chany_bottom_out_37_[0]),
		.chany_bottom_out_39_(sb_0__2__0_chany_bottom_out_39_[0]),
		.chany_bottom_out_41_(sb_0__2__0_chany_bottom_out_41_[0]),
		.chany_bottom_out_43_(sb_0__2__0_chany_bottom_out_43_[0]),
		.chany_bottom_out_45_(sb_0__2__0_chany_bottom_out_45_[0]),
		.chany_bottom_out_47_(sb_0__2__0_chany_bottom_out_47_[0]),
		.chany_bottom_out_49_(sb_0__2__0_chany_bottom_out_49_[0]),
		.chany_bottom_out_51_(sb_0__2__0_chany_bottom_out_51_[0]),
		.chany_bottom_out_53_(sb_0__2__0_chany_bottom_out_53_[0]),
		.chany_bottom_out_55_(sb_0__2__0_chany_bottom_out_55_[0]),
		.chany_bottom_out_57_(sb_0__2__0_chany_bottom_out_57_[0]),
		.chany_bottom_out_59_(sb_0__2__0_chany_bottom_out_59_[0]),
		.chany_bottom_out_61_(sb_0__2__0_chany_bottom_out_61_[0]),
		.chany_bottom_out_63_(sb_0__2__0_chany_bottom_out_63_[0]),
		.chany_bottom_out_65_(sb_0__2__0_chany_bottom_out_65_[0]),
		.chany_bottom_out_67_(sb_0__2__0_chany_bottom_out_67_[0]),
		.chany_bottom_out_69_(sb_0__2__0_chany_bottom_out_69_[0]),
		.chany_bottom_out_71_(sb_0__2__0_chany_bottom_out_71_[0]),
		.chany_bottom_out_73_(sb_0__2__0_chany_bottom_out_73_[0]),
		.chany_bottom_out_75_(sb_0__2__0_chany_bottom_out_75_[0]),
		.chany_bottom_out_77_(sb_0__2__0_chany_bottom_out_77_[0]),
		.chany_bottom_out_79_(sb_0__2__0_chany_bottom_out_79_[0]),
		.chany_bottom_out_81_(sb_0__2__0_chany_bottom_out_81_[0]),
		.chany_bottom_out_83_(sb_0__2__0_chany_bottom_out_83_[0]),
		.chany_bottom_out_85_(sb_0__2__0_chany_bottom_out_85_[0]),
		.chany_bottom_out_87_(sb_0__2__0_chany_bottom_out_87_[0]),
		.chany_bottom_out_89_(sb_0__2__0_chany_bottom_out_89_[0]),
		.chany_bottom_out_91_(sb_0__2__0_chany_bottom_out_91_[0]),
		.chany_bottom_out_93_(sb_0__2__0_chany_bottom_out_93_[0]),
		.chany_bottom_out_95_(sb_0__2__0_chany_bottom_out_95_[0]),
		.chany_bottom_out_97_(sb_0__2__0_chany_bottom_out_97_[0]),
		.chany_bottom_out_99_(sb_0__2__0_chany_bottom_out_99_[0]),
		.chany_bottom_out_101_(sb_0__2__0_chany_bottom_out_101_[0]),
		.chany_bottom_out_103_(sb_0__2__0_chany_bottom_out_103_[0]),
		.chany_bottom_out_105_(sb_0__2__0_chany_bottom_out_105_[0]),
		.chany_bottom_out_107_(sb_0__2__0_chany_bottom_out_107_[0]),
		.chany_bottom_out_109_(sb_0__2__0_chany_bottom_out_109_[0]),
		.chany_bottom_out_111_(sb_0__2__0_chany_bottom_out_111_[0]),
		.chany_bottom_out_113_(sb_0__2__0_chany_bottom_out_113_[0]),
		.chany_bottom_out_115_(sb_0__2__0_chany_bottom_out_115_[0]),
		.chany_bottom_out_117_(sb_0__2__0_chany_bottom_out_117_[0]),
		.chany_bottom_out_119_(sb_0__2__0_chany_bottom_out_119_[0]),
		.chany_bottom_out_121_(sb_0__2__0_chany_bottom_out_121_[0]),
		.chany_bottom_out_123_(sb_0__2__0_chany_bottom_out_123_[0]),
		.chany_bottom_out_125_(sb_0__2__0_chany_bottom_out_125_[0]),
		.chany_bottom_out_127_(sb_0__2__0_chany_bottom_out_127_[0]),
		.chany_bottom_out_129_(sb_0__2__0_chany_bottom_out_129_[0]),
		.chany_bottom_out_131_(sb_0__2__0_chany_bottom_out_131_[0]),
		.chany_bottom_out_133_(sb_0__2__0_chany_bottom_out_133_[0]),
		.chany_bottom_out_135_(sb_0__2__0_chany_bottom_out_135_[0]),
		.chany_bottom_out_137_(sb_0__2__0_chany_bottom_out_137_[0]),
		.chany_bottom_out_139_(sb_0__2__0_chany_bottom_out_139_[0]),
		.chany_bottom_out_141_(sb_0__2__0_chany_bottom_out_141_[0]),
		.chany_bottom_out_143_(sb_0__2__0_chany_bottom_out_143_[0]),
		.chany_bottom_out_145_(sb_0__2__0_chany_bottom_out_145_[0]),
		.chany_bottom_out_147_(sb_0__2__0_chany_bottom_out_147_[0]),
		.chany_bottom_out_149_(sb_0__2__0_chany_bottom_out_149_[0]),
		.chany_bottom_out_151_(sb_0__2__0_chany_bottom_out_151_[0]),
		.chany_bottom_out_153_(sb_0__2__0_chany_bottom_out_153_[0]),
		.chany_bottom_out_155_(sb_0__2__0_chany_bottom_out_155_[0]),
		.chany_bottom_out_157_(sb_0__2__0_chany_bottom_out_157_[0]),
		.chany_bottom_out_159_(sb_0__2__0_chany_bottom_out_159_[0]),
		.chany_bottom_out_161_(sb_0__2__0_chany_bottom_out_161_[0]),
		.chany_bottom_out_163_(sb_0__2__0_chany_bottom_out_163_[0]),
		.chany_bottom_out_165_(sb_0__2__0_chany_bottom_out_165_[0]),
		.chany_bottom_out_167_(sb_0__2__0_chany_bottom_out_167_[0]),
		.chany_bottom_out_169_(sb_0__2__0_chany_bottom_out_169_[0]),
		.chany_bottom_out_171_(sb_0__2__0_chany_bottom_out_171_[0]),
		.chany_bottom_out_173_(sb_0__2__0_chany_bottom_out_173_[0]),
		.chany_bottom_out_175_(sb_0__2__0_chany_bottom_out_175_[0]),
		.chany_bottom_out_177_(sb_0__2__0_chany_bottom_out_177_[0]),
		.chany_bottom_out_179_(sb_0__2__0_chany_bottom_out_179_[0]),
		.chany_bottom_out_181_(sb_0__2__0_chany_bottom_out_181_[0]),
		.chany_bottom_out_183_(sb_0__2__0_chany_bottom_out_183_[0]),
		.chany_bottom_out_185_(sb_0__2__0_chany_bottom_out_185_[0]),
		.chany_bottom_out_187_(sb_0__2__0_chany_bottom_out_187_[0]),
		.chany_bottom_out_189_(sb_0__2__0_chany_bottom_out_189_[0]),
		.chany_bottom_out_191_(sb_0__2__0_chany_bottom_out_191_[0]),
		.chany_bottom_out_193_(sb_0__2__0_chany_bottom_out_193_[0]),
		.chany_bottom_out_195_(sb_0__2__0_chany_bottom_out_195_[0]),
		.chany_bottom_out_197_(sb_0__2__0_chany_bottom_out_197_[0]),
		.chany_bottom_out_199_(sb_0__2__0_chany_bottom_out_199_[0]),
		.ccff_tail(sb_0__2__0_ccff_tail[0]));

	sb_1__0_ sb_1__0_ (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.chany_top_in_1_(cby_1__1__0_chany_out_1_[0]),
		.chany_top_in_3_(cby_1__1__0_chany_out_3_[0]),
		.chany_top_in_5_(cby_1__1__0_chany_out_5_[0]),
		.chany_top_in_7_(cby_1__1__0_chany_out_7_[0]),
		.chany_top_in_9_(cby_1__1__0_chany_out_9_[0]),
		.chany_top_in_11_(cby_1__1__0_chany_out_11_[0]),
		.chany_top_in_13_(cby_1__1__0_chany_out_13_[0]),
		.chany_top_in_15_(cby_1__1__0_chany_out_15_[0]),
		.chany_top_in_17_(cby_1__1__0_chany_out_17_[0]),
		.chany_top_in_19_(cby_1__1__0_chany_out_19_[0]),
		.chany_top_in_21_(cby_1__1__0_chany_out_21_[0]),
		.chany_top_in_23_(cby_1__1__0_chany_out_23_[0]),
		.chany_top_in_25_(cby_1__1__0_chany_out_25_[0]),
		.chany_top_in_27_(cby_1__1__0_chany_out_27_[0]),
		.chany_top_in_29_(cby_1__1__0_chany_out_29_[0]),
		.chany_top_in_31_(cby_1__1__0_chany_out_31_[0]),
		.chany_top_in_33_(cby_1__1__0_chany_out_33_[0]),
		.chany_top_in_35_(cby_1__1__0_chany_out_35_[0]),
		.chany_top_in_37_(cby_1__1__0_chany_out_37_[0]),
		.chany_top_in_39_(cby_1__1__0_chany_out_39_[0]),
		.chany_top_in_41_(cby_1__1__0_chany_out_41_[0]),
		.chany_top_in_43_(cby_1__1__0_chany_out_43_[0]),
		.chany_top_in_45_(cby_1__1__0_chany_out_45_[0]),
		.chany_top_in_47_(cby_1__1__0_chany_out_47_[0]),
		.chany_top_in_49_(cby_1__1__0_chany_out_49_[0]),
		.chany_top_in_51_(cby_1__1__0_chany_out_51_[0]),
		.chany_top_in_53_(cby_1__1__0_chany_out_53_[0]),
		.chany_top_in_55_(cby_1__1__0_chany_out_55_[0]),
		.chany_top_in_57_(cby_1__1__0_chany_out_57_[0]),
		.chany_top_in_59_(cby_1__1__0_chany_out_59_[0]),
		.chany_top_in_61_(cby_1__1__0_chany_out_61_[0]),
		.chany_top_in_63_(cby_1__1__0_chany_out_63_[0]),
		.chany_top_in_65_(cby_1__1__0_chany_out_65_[0]),
		.chany_top_in_67_(cby_1__1__0_chany_out_67_[0]),
		.chany_top_in_69_(cby_1__1__0_chany_out_69_[0]),
		.chany_top_in_71_(cby_1__1__0_chany_out_71_[0]),
		.chany_top_in_73_(cby_1__1__0_chany_out_73_[0]),
		.chany_top_in_75_(cby_1__1__0_chany_out_75_[0]),
		.chany_top_in_77_(cby_1__1__0_chany_out_77_[0]),
		.chany_top_in_79_(cby_1__1__0_chany_out_79_[0]),
		.chany_top_in_81_(cby_1__1__0_chany_out_81_[0]),
		.chany_top_in_83_(cby_1__1__0_chany_out_83_[0]),
		.chany_top_in_85_(cby_1__1__0_chany_out_85_[0]),
		.chany_top_in_87_(cby_1__1__0_chany_out_87_[0]),
		.chany_top_in_89_(cby_1__1__0_chany_out_89_[0]),
		.chany_top_in_91_(cby_1__1__0_chany_out_91_[0]),
		.chany_top_in_93_(cby_1__1__0_chany_out_93_[0]),
		.chany_top_in_95_(cby_1__1__0_chany_out_95_[0]),
		.chany_top_in_97_(cby_1__1__0_chany_out_97_[0]),
		.chany_top_in_99_(cby_1__1__0_chany_out_99_[0]),
		.chany_top_in_101_(cby_1__1__0_chany_out_101_[0]),
		.chany_top_in_103_(cby_1__1__0_chany_out_103_[0]),
		.chany_top_in_105_(cby_1__1__0_chany_out_105_[0]),
		.chany_top_in_107_(cby_1__1__0_chany_out_107_[0]),
		.chany_top_in_109_(cby_1__1__0_chany_out_109_[0]),
		.chany_top_in_111_(cby_1__1__0_chany_out_111_[0]),
		.chany_top_in_113_(cby_1__1__0_chany_out_113_[0]),
		.chany_top_in_115_(cby_1__1__0_chany_out_115_[0]),
		.chany_top_in_117_(cby_1__1__0_chany_out_117_[0]),
		.chany_top_in_119_(cby_1__1__0_chany_out_119_[0]),
		.chany_top_in_121_(cby_1__1__0_chany_out_121_[0]),
		.chany_top_in_123_(cby_1__1__0_chany_out_123_[0]),
		.chany_top_in_125_(cby_1__1__0_chany_out_125_[0]),
		.chany_top_in_127_(cby_1__1__0_chany_out_127_[0]),
		.chany_top_in_129_(cby_1__1__0_chany_out_129_[0]),
		.chany_top_in_131_(cby_1__1__0_chany_out_131_[0]),
		.chany_top_in_133_(cby_1__1__0_chany_out_133_[0]),
		.chany_top_in_135_(cby_1__1__0_chany_out_135_[0]),
		.chany_top_in_137_(cby_1__1__0_chany_out_137_[0]),
		.chany_top_in_139_(cby_1__1__0_chany_out_139_[0]),
		.chany_top_in_141_(cby_1__1__0_chany_out_141_[0]),
		.chany_top_in_143_(cby_1__1__0_chany_out_143_[0]),
		.chany_top_in_145_(cby_1__1__0_chany_out_145_[0]),
		.chany_top_in_147_(cby_1__1__0_chany_out_147_[0]),
		.chany_top_in_149_(cby_1__1__0_chany_out_149_[0]),
		.chany_top_in_151_(cby_1__1__0_chany_out_151_[0]),
		.chany_top_in_153_(cby_1__1__0_chany_out_153_[0]),
		.chany_top_in_155_(cby_1__1__0_chany_out_155_[0]),
		.chany_top_in_157_(cby_1__1__0_chany_out_157_[0]),
		.chany_top_in_159_(cby_1__1__0_chany_out_159_[0]),
		.chany_top_in_161_(cby_1__1__0_chany_out_161_[0]),
		.chany_top_in_163_(cby_1__1__0_chany_out_163_[0]),
		.chany_top_in_165_(cby_1__1__0_chany_out_165_[0]),
		.chany_top_in_167_(cby_1__1__0_chany_out_167_[0]),
		.chany_top_in_169_(cby_1__1__0_chany_out_169_[0]),
		.chany_top_in_171_(cby_1__1__0_chany_out_171_[0]),
		.chany_top_in_173_(cby_1__1__0_chany_out_173_[0]),
		.chany_top_in_175_(cby_1__1__0_chany_out_175_[0]),
		.chany_top_in_177_(cby_1__1__0_chany_out_177_[0]),
		.chany_top_in_179_(cby_1__1__0_chany_out_179_[0]),
		.chany_top_in_181_(cby_1__1__0_chany_out_181_[0]),
		.chany_top_in_183_(cby_1__1__0_chany_out_183_[0]),
		.chany_top_in_185_(cby_1__1__0_chany_out_185_[0]),
		.chany_top_in_187_(cby_1__1__0_chany_out_187_[0]),
		.chany_top_in_189_(cby_1__1__0_chany_out_189_[0]),
		.chany_top_in_191_(cby_1__1__0_chany_out_191_[0]),
		.chany_top_in_193_(cby_1__1__0_chany_out_193_[0]),
		.chany_top_in_195_(cby_1__1__0_chany_out_195_[0]),
		.chany_top_in_197_(cby_1__1__0_chany_out_197_[0]),
		.chany_top_in_199_(cby_1__1__0_chany_out_199_[0]),
		.top_left_grid_pin_44_(grid_clb_spypad_0_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_spypad_0_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_spypad_0_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_spypad_0_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_spypad_0_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_spypad_0_right_width_0_height_0__pin_49_lower[0]),
		.top_left_grid_pin_50_(grid_clb_spypad_0_right_width_0_height_0__pin_50_lower[0]),
		.top_left_grid_pin_51_(grid_clb_spypad_0_right_width_0_height_0__pin_51_lower[0]),
		.top_left_grid_pin_52_(grid_clb_spypad_0_right_width_0_height_0__pin_52_lower[0]),
		.top_left_grid_pin_53_(grid_clb_spypad_0_right_width_0_height_0__pin_53_lower[0]),
		.chanx_right_in_1_(cbx_1__0__1_chanx_out_1_[0]),
		.chanx_right_in_3_(cbx_1__0__1_chanx_out_3_[0]),
		.chanx_right_in_5_(cbx_1__0__1_chanx_out_5_[0]),
		.chanx_right_in_7_(cbx_1__0__1_chanx_out_7_[0]),
		.chanx_right_in_9_(cbx_1__0__1_chanx_out_9_[0]),
		.chanx_right_in_11_(cbx_1__0__1_chanx_out_11_[0]),
		.chanx_right_in_13_(cbx_1__0__1_chanx_out_13_[0]),
		.chanx_right_in_15_(cbx_1__0__1_chanx_out_15_[0]),
		.chanx_right_in_17_(cbx_1__0__1_chanx_out_17_[0]),
		.chanx_right_in_19_(cbx_1__0__1_chanx_out_19_[0]),
		.chanx_right_in_21_(cbx_1__0__1_chanx_out_21_[0]),
		.chanx_right_in_23_(cbx_1__0__1_chanx_out_23_[0]),
		.chanx_right_in_25_(cbx_1__0__1_chanx_out_25_[0]),
		.chanx_right_in_27_(cbx_1__0__1_chanx_out_27_[0]),
		.chanx_right_in_29_(cbx_1__0__1_chanx_out_29_[0]),
		.chanx_right_in_31_(cbx_1__0__1_chanx_out_31_[0]),
		.chanx_right_in_33_(cbx_1__0__1_chanx_out_33_[0]),
		.chanx_right_in_35_(cbx_1__0__1_chanx_out_35_[0]),
		.chanx_right_in_37_(cbx_1__0__1_chanx_out_37_[0]),
		.chanx_right_in_39_(cbx_1__0__1_chanx_out_39_[0]),
		.chanx_right_in_41_(cbx_1__0__1_chanx_out_41_[0]),
		.chanx_right_in_43_(cbx_1__0__1_chanx_out_43_[0]),
		.chanx_right_in_45_(cbx_1__0__1_chanx_out_45_[0]),
		.chanx_right_in_47_(cbx_1__0__1_chanx_out_47_[0]),
		.chanx_right_in_49_(cbx_1__0__1_chanx_out_49_[0]),
		.chanx_right_in_51_(cbx_1__0__1_chanx_out_51_[0]),
		.chanx_right_in_53_(cbx_1__0__1_chanx_out_53_[0]),
		.chanx_right_in_55_(cbx_1__0__1_chanx_out_55_[0]),
		.chanx_right_in_57_(cbx_1__0__1_chanx_out_57_[0]),
		.chanx_right_in_59_(cbx_1__0__1_chanx_out_59_[0]),
		.chanx_right_in_61_(cbx_1__0__1_chanx_out_61_[0]),
		.chanx_right_in_63_(cbx_1__0__1_chanx_out_63_[0]),
		.chanx_right_in_65_(cbx_1__0__1_chanx_out_65_[0]),
		.chanx_right_in_67_(cbx_1__0__1_chanx_out_67_[0]),
		.chanx_right_in_69_(cbx_1__0__1_chanx_out_69_[0]),
		.chanx_right_in_71_(cbx_1__0__1_chanx_out_71_[0]),
		.chanx_right_in_73_(cbx_1__0__1_chanx_out_73_[0]),
		.chanx_right_in_75_(cbx_1__0__1_chanx_out_75_[0]),
		.chanx_right_in_77_(cbx_1__0__1_chanx_out_77_[0]),
		.chanx_right_in_79_(cbx_1__0__1_chanx_out_79_[0]),
		.chanx_right_in_81_(cbx_1__0__1_chanx_out_81_[0]),
		.chanx_right_in_83_(cbx_1__0__1_chanx_out_83_[0]),
		.chanx_right_in_85_(cbx_1__0__1_chanx_out_85_[0]),
		.chanx_right_in_87_(cbx_1__0__1_chanx_out_87_[0]),
		.chanx_right_in_89_(cbx_1__0__1_chanx_out_89_[0]),
		.chanx_right_in_91_(cbx_1__0__1_chanx_out_91_[0]),
		.chanx_right_in_93_(cbx_1__0__1_chanx_out_93_[0]),
		.chanx_right_in_95_(cbx_1__0__1_chanx_out_95_[0]),
		.chanx_right_in_97_(cbx_1__0__1_chanx_out_97_[0]),
		.chanx_right_in_99_(cbx_1__0__1_chanx_out_99_[0]),
		.chanx_right_in_101_(cbx_1__0__1_chanx_out_101_[0]),
		.chanx_right_in_103_(cbx_1__0__1_chanx_out_103_[0]),
		.chanx_right_in_105_(cbx_1__0__1_chanx_out_105_[0]),
		.chanx_right_in_107_(cbx_1__0__1_chanx_out_107_[0]),
		.chanx_right_in_109_(cbx_1__0__1_chanx_out_109_[0]),
		.chanx_right_in_111_(cbx_1__0__1_chanx_out_111_[0]),
		.chanx_right_in_113_(cbx_1__0__1_chanx_out_113_[0]),
		.chanx_right_in_115_(cbx_1__0__1_chanx_out_115_[0]),
		.chanx_right_in_117_(cbx_1__0__1_chanx_out_117_[0]),
		.chanx_right_in_119_(cbx_1__0__1_chanx_out_119_[0]),
		.chanx_right_in_121_(cbx_1__0__1_chanx_out_121_[0]),
		.chanx_right_in_123_(cbx_1__0__1_chanx_out_123_[0]),
		.chanx_right_in_125_(cbx_1__0__1_chanx_out_125_[0]),
		.chanx_right_in_127_(cbx_1__0__1_chanx_out_127_[0]),
		.chanx_right_in_129_(cbx_1__0__1_chanx_out_129_[0]),
		.chanx_right_in_131_(cbx_1__0__1_chanx_out_131_[0]),
		.chanx_right_in_133_(cbx_1__0__1_chanx_out_133_[0]),
		.chanx_right_in_135_(cbx_1__0__1_chanx_out_135_[0]),
		.chanx_right_in_137_(cbx_1__0__1_chanx_out_137_[0]),
		.chanx_right_in_139_(cbx_1__0__1_chanx_out_139_[0]),
		.chanx_right_in_141_(cbx_1__0__1_chanx_out_141_[0]),
		.chanx_right_in_143_(cbx_1__0__1_chanx_out_143_[0]),
		.chanx_right_in_145_(cbx_1__0__1_chanx_out_145_[0]),
		.chanx_right_in_147_(cbx_1__0__1_chanx_out_147_[0]),
		.chanx_right_in_149_(cbx_1__0__1_chanx_out_149_[0]),
		.chanx_right_in_151_(cbx_1__0__1_chanx_out_151_[0]),
		.chanx_right_in_153_(cbx_1__0__1_chanx_out_153_[0]),
		.chanx_right_in_155_(cbx_1__0__1_chanx_out_155_[0]),
		.chanx_right_in_157_(cbx_1__0__1_chanx_out_157_[0]),
		.chanx_right_in_159_(cbx_1__0__1_chanx_out_159_[0]),
		.chanx_right_in_161_(cbx_1__0__1_chanx_out_161_[0]),
		.chanx_right_in_163_(cbx_1__0__1_chanx_out_163_[0]),
		.chanx_right_in_165_(cbx_1__0__1_chanx_out_165_[0]),
		.chanx_right_in_167_(cbx_1__0__1_chanx_out_167_[0]),
		.chanx_right_in_169_(cbx_1__0__1_chanx_out_169_[0]),
		.chanx_right_in_171_(cbx_1__0__1_chanx_out_171_[0]),
		.chanx_right_in_173_(cbx_1__0__1_chanx_out_173_[0]),
		.chanx_right_in_175_(cbx_1__0__1_chanx_out_175_[0]),
		.chanx_right_in_177_(cbx_1__0__1_chanx_out_177_[0]),
		.chanx_right_in_179_(cbx_1__0__1_chanx_out_179_[0]),
		.chanx_right_in_181_(cbx_1__0__1_chanx_out_181_[0]),
		.chanx_right_in_183_(cbx_1__0__1_chanx_out_183_[0]),
		.chanx_right_in_185_(cbx_1__0__1_chanx_out_185_[0]),
		.chanx_right_in_187_(cbx_1__0__1_chanx_out_187_[0]),
		.chanx_right_in_189_(cbx_1__0__1_chanx_out_189_[0]),
		.chanx_right_in_191_(cbx_1__0__1_chanx_out_191_[0]),
		.chanx_right_in_193_(cbx_1__0__1_chanx_out_193_[0]),
		.chanx_right_in_195_(cbx_1__0__1_chanx_out_195_[0]),
		.chanx_right_in_197_(cbx_1__0__1_chanx_out_197_[0]),
		.chanx_right_in_199_(cbx_1__0__1_chanx_out_199_[0]),
		.right_top_grid_pin_54_(grid_clb_1_bottom_width_0_height_0__pin_54_upper[0]),
		.right_top_grid_pin_55_(grid_clb_1_bottom_width_0_height_0__pin_55_upper[0]),
		.right_top_grid_pin_56_(grid_clb_1_bottom_width_0_height_0__pin_56_upper[0]),
		.right_top_grid_pin_57_(grid_clb_1_bottom_width_0_height_0__pin_57_upper[0]),
		.right_top_grid_pin_58_(grid_clb_1_bottom_width_0_height_0__pin_58_upper[0]),
		.right_top_grid_pin_59_(grid_clb_1_bottom_width_0_height_0__pin_59_upper[0]),
		.right_top_grid_pin_60_(grid_clb_1_bottom_width_0_height_0__pin_60_upper[0]),
		.right_top_grid_pin_61_(grid_clb_1_bottom_width_0_height_0__pin_61_upper[0]),
		.right_top_grid_pin_62_(grid_clb_1_bottom_width_0_height_0__pin_62_upper[0]),
		.right_top_grid_pin_63_(grid_clb_1_bottom_width_0_height_0__pin_63_upper[0]),
		.right_top_grid_pin_66_(grid_clb_1_bottom_width_0_height_0__pin_66_upper[0]),
		.right_top_grid_pin_67_(grid_clb_1_bottom_width_0_height_0__pin_67_upper[0]),
		.right_bottom_grid_pin_1_(grid_io_bottom_1_top_width_0_height_0__pin_1_upper[0]),
		.chanx_left_in_0_(cbx_1__0__0_chanx_out_0_[0]),
		.chanx_left_in_2_(cbx_1__0__0_chanx_out_2_[0]),
		.chanx_left_in_4_(cbx_1__0__0_chanx_out_4_[0]),
		.chanx_left_in_6_(cbx_1__0__0_chanx_out_6_[0]),
		.chanx_left_in_8_(cbx_1__0__0_chanx_out_8_[0]),
		.chanx_left_in_10_(cbx_1__0__0_chanx_out_10_[0]),
		.chanx_left_in_12_(cbx_1__0__0_chanx_out_12_[0]),
		.chanx_left_in_14_(cbx_1__0__0_chanx_out_14_[0]),
		.chanx_left_in_16_(cbx_1__0__0_chanx_out_16_[0]),
		.chanx_left_in_18_(cbx_1__0__0_chanx_out_18_[0]),
		.chanx_left_in_20_(cbx_1__0__0_chanx_out_20_[0]),
		.chanx_left_in_22_(cbx_1__0__0_chanx_out_22_[0]),
		.chanx_left_in_24_(cbx_1__0__0_chanx_out_24_[0]),
		.chanx_left_in_26_(cbx_1__0__0_chanx_out_26_[0]),
		.chanx_left_in_28_(cbx_1__0__0_chanx_out_28_[0]),
		.chanx_left_in_30_(cbx_1__0__0_chanx_out_30_[0]),
		.chanx_left_in_32_(cbx_1__0__0_chanx_out_32_[0]),
		.chanx_left_in_34_(cbx_1__0__0_chanx_out_34_[0]),
		.chanx_left_in_36_(cbx_1__0__0_chanx_out_36_[0]),
		.chanx_left_in_38_(cbx_1__0__0_chanx_out_38_[0]),
		.chanx_left_in_40_(cbx_1__0__0_chanx_out_40_[0]),
		.chanx_left_in_42_(cbx_1__0__0_chanx_out_42_[0]),
		.chanx_left_in_44_(cbx_1__0__0_chanx_out_44_[0]),
		.chanx_left_in_46_(cbx_1__0__0_chanx_out_46_[0]),
		.chanx_left_in_48_(cbx_1__0__0_chanx_out_48_[0]),
		.chanx_left_in_50_(cbx_1__0__0_chanx_out_50_[0]),
		.chanx_left_in_52_(cbx_1__0__0_chanx_out_52_[0]),
		.chanx_left_in_54_(cbx_1__0__0_chanx_out_54_[0]),
		.chanx_left_in_56_(cbx_1__0__0_chanx_out_56_[0]),
		.chanx_left_in_58_(cbx_1__0__0_chanx_out_58_[0]),
		.chanx_left_in_60_(cbx_1__0__0_chanx_out_60_[0]),
		.chanx_left_in_62_(cbx_1__0__0_chanx_out_62_[0]),
		.chanx_left_in_64_(cbx_1__0__0_chanx_out_64_[0]),
		.chanx_left_in_66_(cbx_1__0__0_chanx_out_66_[0]),
		.chanx_left_in_68_(cbx_1__0__0_chanx_out_68_[0]),
		.chanx_left_in_70_(cbx_1__0__0_chanx_out_70_[0]),
		.chanx_left_in_72_(cbx_1__0__0_chanx_out_72_[0]),
		.chanx_left_in_74_(cbx_1__0__0_chanx_out_74_[0]),
		.chanx_left_in_76_(cbx_1__0__0_chanx_out_76_[0]),
		.chanx_left_in_78_(cbx_1__0__0_chanx_out_78_[0]),
		.chanx_left_in_80_(cbx_1__0__0_chanx_out_80_[0]),
		.chanx_left_in_82_(cbx_1__0__0_chanx_out_82_[0]),
		.chanx_left_in_84_(cbx_1__0__0_chanx_out_84_[0]),
		.chanx_left_in_86_(cbx_1__0__0_chanx_out_86_[0]),
		.chanx_left_in_88_(cbx_1__0__0_chanx_out_88_[0]),
		.chanx_left_in_90_(cbx_1__0__0_chanx_out_90_[0]),
		.chanx_left_in_92_(cbx_1__0__0_chanx_out_92_[0]),
		.chanx_left_in_94_(cbx_1__0__0_chanx_out_94_[0]),
		.chanx_left_in_96_(cbx_1__0__0_chanx_out_96_[0]),
		.chanx_left_in_98_(cbx_1__0__0_chanx_out_98_[0]),
		.chanx_left_in_100_(cbx_1__0__0_chanx_out_100_[0]),
		.chanx_left_in_102_(cbx_1__0__0_chanx_out_102_[0]),
		.chanx_left_in_104_(cbx_1__0__0_chanx_out_104_[0]),
		.chanx_left_in_106_(cbx_1__0__0_chanx_out_106_[0]),
		.chanx_left_in_108_(cbx_1__0__0_chanx_out_108_[0]),
		.chanx_left_in_110_(cbx_1__0__0_chanx_out_110_[0]),
		.chanx_left_in_112_(cbx_1__0__0_chanx_out_112_[0]),
		.chanx_left_in_114_(cbx_1__0__0_chanx_out_114_[0]),
		.chanx_left_in_116_(cbx_1__0__0_chanx_out_116_[0]),
		.chanx_left_in_118_(cbx_1__0__0_chanx_out_118_[0]),
		.chanx_left_in_120_(cbx_1__0__0_chanx_out_120_[0]),
		.chanx_left_in_122_(cbx_1__0__0_chanx_out_122_[0]),
		.chanx_left_in_124_(cbx_1__0__0_chanx_out_124_[0]),
		.chanx_left_in_126_(cbx_1__0__0_chanx_out_126_[0]),
		.chanx_left_in_128_(cbx_1__0__0_chanx_out_128_[0]),
		.chanx_left_in_130_(cbx_1__0__0_chanx_out_130_[0]),
		.chanx_left_in_132_(cbx_1__0__0_chanx_out_132_[0]),
		.chanx_left_in_134_(cbx_1__0__0_chanx_out_134_[0]),
		.chanx_left_in_136_(cbx_1__0__0_chanx_out_136_[0]),
		.chanx_left_in_138_(cbx_1__0__0_chanx_out_138_[0]),
		.chanx_left_in_140_(cbx_1__0__0_chanx_out_140_[0]),
		.chanx_left_in_142_(cbx_1__0__0_chanx_out_142_[0]),
		.chanx_left_in_144_(cbx_1__0__0_chanx_out_144_[0]),
		.chanx_left_in_146_(cbx_1__0__0_chanx_out_146_[0]),
		.chanx_left_in_148_(cbx_1__0__0_chanx_out_148_[0]),
		.chanx_left_in_150_(cbx_1__0__0_chanx_out_150_[0]),
		.chanx_left_in_152_(cbx_1__0__0_chanx_out_152_[0]),
		.chanx_left_in_154_(cbx_1__0__0_chanx_out_154_[0]),
		.chanx_left_in_156_(cbx_1__0__0_chanx_out_156_[0]),
		.chanx_left_in_158_(cbx_1__0__0_chanx_out_158_[0]),
		.chanx_left_in_160_(cbx_1__0__0_chanx_out_160_[0]),
		.chanx_left_in_162_(cbx_1__0__0_chanx_out_162_[0]),
		.chanx_left_in_164_(cbx_1__0__0_chanx_out_164_[0]),
		.chanx_left_in_166_(cbx_1__0__0_chanx_out_166_[0]),
		.chanx_left_in_168_(cbx_1__0__0_chanx_out_168_[0]),
		.chanx_left_in_170_(cbx_1__0__0_chanx_out_170_[0]),
		.chanx_left_in_172_(cbx_1__0__0_chanx_out_172_[0]),
		.chanx_left_in_174_(cbx_1__0__0_chanx_out_174_[0]),
		.chanx_left_in_176_(cbx_1__0__0_chanx_out_176_[0]),
		.chanx_left_in_178_(cbx_1__0__0_chanx_out_178_[0]),
		.chanx_left_in_180_(cbx_1__0__0_chanx_out_180_[0]),
		.chanx_left_in_182_(cbx_1__0__0_chanx_out_182_[0]),
		.chanx_left_in_184_(cbx_1__0__0_chanx_out_184_[0]),
		.chanx_left_in_186_(cbx_1__0__0_chanx_out_186_[0]),
		.chanx_left_in_188_(cbx_1__0__0_chanx_out_188_[0]),
		.chanx_left_in_190_(cbx_1__0__0_chanx_out_190_[0]),
		.chanx_left_in_192_(cbx_1__0__0_chanx_out_192_[0]),
		.chanx_left_in_194_(cbx_1__0__0_chanx_out_194_[0]),
		.chanx_left_in_196_(cbx_1__0__0_chanx_out_196_[0]),
		.chanx_left_in_198_(cbx_1__0__0_chanx_out_198_[0]),
		.left_top_grid_pin_54_(grid_clb_spypad_0_bottom_width_0_height_0__pin_54_lower[0]),
		.left_top_grid_pin_55_(grid_clb_spypad_0_bottom_width_0_height_0__pin_55_lower[0]),
		.left_top_grid_pin_56_(grid_clb_spypad_0_bottom_width_0_height_0__pin_56_lower[0]),
		.left_top_grid_pin_57_(grid_clb_spypad_0_bottom_width_0_height_0__pin_57_lower[0]),
		.left_top_grid_pin_58_(grid_clb_spypad_0_bottom_width_0_height_0__pin_58_lower[0]),
		.left_top_grid_pin_59_(grid_clb_spypad_0_bottom_width_0_height_0__pin_59_lower[0]),
		.left_top_grid_pin_60_(grid_clb_spypad_0_bottom_width_0_height_0__pin_60_lower[0]),
		.left_top_grid_pin_61_(grid_clb_spypad_0_bottom_width_0_height_0__pin_61_lower[0]),
		.left_top_grid_pin_62_(grid_clb_spypad_0_bottom_width_0_height_0__pin_62_lower[0]),
		.left_top_grid_pin_63_(grid_clb_spypad_0_bottom_width_0_height_0__pin_63_lower[0]),
		.left_top_grid_pin_66_(grid_clb_spypad_0_bottom_width_0_height_0__pin_66_lower[0]),
		.left_top_grid_pin_67_(grid_clb_spypad_0_bottom_width_0_height_0__pin_67_lower[0]),
		.left_bottom_grid_pin_1_(grid_io_bottom_0_top_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_io_left_0_ccff_tail[0]),
		.chany_top_out_0_(sb_1__0__0_chany_top_out_0_[0]),
		.chany_top_out_2_(sb_1__0__0_chany_top_out_2_[0]),
		.chany_top_out_4_(sb_1__0__0_chany_top_out_4_[0]),
		.chany_top_out_6_(sb_1__0__0_chany_top_out_6_[0]),
		.chany_top_out_8_(sb_1__0__0_chany_top_out_8_[0]),
		.chany_top_out_10_(sb_1__0__0_chany_top_out_10_[0]),
		.chany_top_out_12_(sb_1__0__0_chany_top_out_12_[0]),
		.chany_top_out_14_(sb_1__0__0_chany_top_out_14_[0]),
		.chany_top_out_16_(sb_1__0__0_chany_top_out_16_[0]),
		.chany_top_out_18_(sb_1__0__0_chany_top_out_18_[0]),
		.chany_top_out_20_(sb_1__0__0_chany_top_out_20_[0]),
		.chany_top_out_22_(sb_1__0__0_chany_top_out_22_[0]),
		.chany_top_out_24_(sb_1__0__0_chany_top_out_24_[0]),
		.chany_top_out_26_(sb_1__0__0_chany_top_out_26_[0]),
		.chany_top_out_28_(sb_1__0__0_chany_top_out_28_[0]),
		.chany_top_out_30_(sb_1__0__0_chany_top_out_30_[0]),
		.chany_top_out_32_(sb_1__0__0_chany_top_out_32_[0]),
		.chany_top_out_34_(sb_1__0__0_chany_top_out_34_[0]),
		.chany_top_out_36_(sb_1__0__0_chany_top_out_36_[0]),
		.chany_top_out_38_(sb_1__0__0_chany_top_out_38_[0]),
		.chany_top_out_40_(sb_1__0__0_chany_top_out_40_[0]),
		.chany_top_out_42_(sb_1__0__0_chany_top_out_42_[0]),
		.chany_top_out_44_(sb_1__0__0_chany_top_out_44_[0]),
		.chany_top_out_46_(sb_1__0__0_chany_top_out_46_[0]),
		.chany_top_out_48_(sb_1__0__0_chany_top_out_48_[0]),
		.chany_top_out_50_(sb_1__0__0_chany_top_out_50_[0]),
		.chany_top_out_52_(sb_1__0__0_chany_top_out_52_[0]),
		.chany_top_out_54_(sb_1__0__0_chany_top_out_54_[0]),
		.chany_top_out_56_(sb_1__0__0_chany_top_out_56_[0]),
		.chany_top_out_58_(sb_1__0__0_chany_top_out_58_[0]),
		.chany_top_out_60_(sb_1__0__0_chany_top_out_60_[0]),
		.chany_top_out_62_(sb_1__0__0_chany_top_out_62_[0]),
		.chany_top_out_64_(sb_1__0__0_chany_top_out_64_[0]),
		.chany_top_out_66_(sb_1__0__0_chany_top_out_66_[0]),
		.chany_top_out_68_(sb_1__0__0_chany_top_out_68_[0]),
		.chany_top_out_70_(sb_1__0__0_chany_top_out_70_[0]),
		.chany_top_out_72_(sb_1__0__0_chany_top_out_72_[0]),
		.chany_top_out_74_(sb_1__0__0_chany_top_out_74_[0]),
		.chany_top_out_76_(sb_1__0__0_chany_top_out_76_[0]),
		.chany_top_out_78_(sb_1__0__0_chany_top_out_78_[0]),
		.chany_top_out_80_(sb_1__0__0_chany_top_out_80_[0]),
		.chany_top_out_82_(sb_1__0__0_chany_top_out_82_[0]),
		.chany_top_out_84_(sb_1__0__0_chany_top_out_84_[0]),
		.chany_top_out_86_(sb_1__0__0_chany_top_out_86_[0]),
		.chany_top_out_88_(sb_1__0__0_chany_top_out_88_[0]),
		.chany_top_out_90_(sb_1__0__0_chany_top_out_90_[0]),
		.chany_top_out_92_(sb_1__0__0_chany_top_out_92_[0]),
		.chany_top_out_94_(sb_1__0__0_chany_top_out_94_[0]),
		.chany_top_out_96_(sb_1__0__0_chany_top_out_96_[0]),
		.chany_top_out_98_(sb_1__0__0_chany_top_out_98_[0]),
		.chany_top_out_100_(sb_1__0__0_chany_top_out_100_[0]),
		.chany_top_out_102_(sb_1__0__0_chany_top_out_102_[0]),
		.chany_top_out_104_(sb_1__0__0_chany_top_out_104_[0]),
		.chany_top_out_106_(sb_1__0__0_chany_top_out_106_[0]),
		.chany_top_out_108_(sb_1__0__0_chany_top_out_108_[0]),
		.chany_top_out_110_(sb_1__0__0_chany_top_out_110_[0]),
		.chany_top_out_112_(sb_1__0__0_chany_top_out_112_[0]),
		.chany_top_out_114_(sb_1__0__0_chany_top_out_114_[0]),
		.chany_top_out_116_(sb_1__0__0_chany_top_out_116_[0]),
		.chany_top_out_118_(sb_1__0__0_chany_top_out_118_[0]),
		.chany_top_out_120_(sb_1__0__0_chany_top_out_120_[0]),
		.chany_top_out_122_(sb_1__0__0_chany_top_out_122_[0]),
		.chany_top_out_124_(sb_1__0__0_chany_top_out_124_[0]),
		.chany_top_out_126_(sb_1__0__0_chany_top_out_126_[0]),
		.chany_top_out_128_(sb_1__0__0_chany_top_out_128_[0]),
		.chany_top_out_130_(sb_1__0__0_chany_top_out_130_[0]),
		.chany_top_out_132_(sb_1__0__0_chany_top_out_132_[0]),
		.chany_top_out_134_(sb_1__0__0_chany_top_out_134_[0]),
		.chany_top_out_136_(sb_1__0__0_chany_top_out_136_[0]),
		.chany_top_out_138_(sb_1__0__0_chany_top_out_138_[0]),
		.chany_top_out_140_(sb_1__0__0_chany_top_out_140_[0]),
		.chany_top_out_142_(sb_1__0__0_chany_top_out_142_[0]),
		.chany_top_out_144_(sb_1__0__0_chany_top_out_144_[0]),
		.chany_top_out_146_(sb_1__0__0_chany_top_out_146_[0]),
		.chany_top_out_148_(sb_1__0__0_chany_top_out_148_[0]),
		.chany_top_out_150_(sb_1__0__0_chany_top_out_150_[0]),
		.chany_top_out_152_(sb_1__0__0_chany_top_out_152_[0]),
		.chany_top_out_154_(sb_1__0__0_chany_top_out_154_[0]),
		.chany_top_out_156_(sb_1__0__0_chany_top_out_156_[0]),
		.chany_top_out_158_(sb_1__0__0_chany_top_out_158_[0]),
		.chany_top_out_160_(sb_1__0__0_chany_top_out_160_[0]),
		.chany_top_out_162_(sb_1__0__0_chany_top_out_162_[0]),
		.chany_top_out_164_(sb_1__0__0_chany_top_out_164_[0]),
		.chany_top_out_166_(sb_1__0__0_chany_top_out_166_[0]),
		.chany_top_out_168_(sb_1__0__0_chany_top_out_168_[0]),
		.chany_top_out_170_(sb_1__0__0_chany_top_out_170_[0]),
		.chany_top_out_172_(sb_1__0__0_chany_top_out_172_[0]),
		.chany_top_out_174_(sb_1__0__0_chany_top_out_174_[0]),
		.chany_top_out_176_(sb_1__0__0_chany_top_out_176_[0]),
		.chany_top_out_178_(sb_1__0__0_chany_top_out_178_[0]),
		.chany_top_out_180_(sb_1__0__0_chany_top_out_180_[0]),
		.chany_top_out_182_(sb_1__0__0_chany_top_out_182_[0]),
		.chany_top_out_184_(sb_1__0__0_chany_top_out_184_[0]),
		.chany_top_out_186_(sb_1__0__0_chany_top_out_186_[0]),
		.chany_top_out_188_(sb_1__0__0_chany_top_out_188_[0]),
		.chany_top_out_190_(sb_1__0__0_chany_top_out_190_[0]),
		.chany_top_out_192_(sb_1__0__0_chany_top_out_192_[0]),
		.chany_top_out_194_(sb_1__0__0_chany_top_out_194_[0]),
		.chany_top_out_196_(sb_1__0__0_chany_top_out_196_[0]),
		.chany_top_out_198_(sb_1__0__0_chany_top_out_198_[0]),
		.chanx_right_out_0_(sb_1__0__0_chanx_right_out_0_[0]),
		.chanx_right_out_2_(sb_1__0__0_chanx_right_out_2_[0]),
		.chanx_right_out_4_(sb_1__0__0_chanx_right_out_4_[0]),
		.chanx_right_out_6_(sb_1__0__0_chanx_right_out_6_[0]),
		.chanx_right_out_8_(sb_1__0__0_chanx_right_out_8_[0]),
		.chanx_right_out_10_(sb_1__0__0_chanx_right_out_10_[0]),
		.chanx_right_out_12_(sb_1__0__0_chanx_right_out_12_[0]),
		.chanx_right_out_14_(sb_1__0__0_chanx_right_out_14_[0]),
		.chanx_right_out_16_(sb_1__0__0_chanx_right_out_16_[0]),
		.chanx_right_out_18_(sb_1__0__0_chanx_right_out_18_[0]),
		.chanx_right_out_20_(sb_1__0__0_chanx_right_out_20_[0]),
		.chanx_right_out_22_(sb_1__0__0_chanx_right_out_22_[0]),
		.chanx_right_out_24_(sb_1__0__0_chanx_right_out_24_[0]),
		.chanx_right_out_26_(sb_1__0__0_chanx_right_out_26_[0]),
		.chanx_right_out_28_(sb_1__0__0_chanx_right_out_28_[0]),
		.chanx_right_out_30_(sb_1__0__0_chanx_right_out_30_[0]),
		.chanx_right_out_32_(sb_1__0__0_chanx_right_out_32_[0]),
		.chanx_right_out_34_(sb_1__0__0_chanx_right_out_34_[0]),
		.chanx_right_out_36_(sb_1__0__0_chanx_right_out_36_[0]),
		.chanx_right_out_38_(sb_1__0__0_chanx_right_out_38_[0]),
		.chanx_right_out_40_(sb_1__0__0_chanx_right_out_40_[0]),
		.chanx_right_out_42_(sb_1__0__0_chanx_right_out_42_[0]),
		.chanx_right_out_44_(sb_1__0__0_chanx_right_out_44_[0]),
		.chanx_right_out_46_(sb_1__0__0_chanx_right_out_46_[0]),
		.chanx_right_out_48_(sb_1__0__0_chanx_right_out_48_[0]),
		.chanx_right_out_50_(sb_1__0__0_chanx_right_out_50_[0]),
		.chanx_right_out_52_(sb_1__0__0_chanx_right_out_52_[0]),
		.chanx_right_out_54_(sb_1__0__0_chanx_right_out_54_[0]),
		.chanx_right_out_56_(sb_1__0__0_chanx_right_out_56_[0]),
		.chanx_right_out_58_(sb_1__0__0_chanx_right_out_58_[0]),
		.chanx_right_out_60_(sb_1__0__0_chanx_right_out_60_[0]),
		.chanx_right_out_62_(sb_1__0__0_chanx_right_out_62_[0]),
		.chanx_right_out_64_(sb_1__0__0_chanx_right_out_64_[0]),
		.chanx_right_out_66_(sb_1__0__0_chanx_right_out_66_[0]),
		.chanx_right_out_68_(sb_1__0__0_chanx_right_out_68_[0]),
		.chanx_right_out_70_(sb_1__0__0_chanx_right_out_70_[0]),
		.chanx_right_out_72_(sb_1__0__0_chanx_right_out_72_[0]),
		.chanx_right_out_74_(sb_1__0__0_chanx_right_out_74_[0]),
		.chanx_right_out_76_(sb_1__0__0_chanx_right_out_76_[0]),
		.chanx_right_out_78_(sb_1__0__0_chanx_right_out_78_[0]),
		.chanx_right_out_80_(sb_1__0__0_chanx_right_out_80_[0]),
		.chanx_right_out_82_(sb_1__0__0_chanx_right_out_82_[0]),
		.chanx_right_out_84_(sb_1__0__0_chanx_right_out_84_[0]),
		.chanx_right_out_86_(sb_1__0__0_chanx_right_out_86_[0]),
		.chanx_right_out_88_(sb_1__0__0_chanx_right_out_88_[0]),
		.chanx_right_out_90_(sb_1__0__0_chanx_right_out_90_[0]),
		.chanx_right_out_92_(sb_1__0__0_chanx_right_out_92_[0]),
		.chanx_right_out_94_(sb_1__0__0_chanx_right_out_94_[0]),
		.chanx_right_out_96_(sb_1__0__0_chanx_right_out_96_[0]),
		.chanx_right_out_98_(sb_1__0__0_chanx_right_out_98_[0]),
		.chanx_right_out_100_(sb_1__0__0_chanx_right_out_100_[0]),
		.chanx_right_out_102_(sb_1__0__0_chanx_right_out_102_[0]),
		.chanx_right_out_104_(sb_1__0__0_chanx_right_out_104_[0]),
		.chanx_right_out_106_(sb_1__0__0_chanx_right_out_106_[0]),
		.chanx_right_out_108_(sb_1__0__0_chanx_right_out_108_[0]),
		.chanx_right_out_110_(sb_1__0__0_chanx_right_out_110_[0]),
		.chanx_right_out_112_(sb_1__0__0_chanx_right_out_112_[0]),
		.chanx_right_out_114_(sb_1__0__0_chanx_right_out_114_[0]),
		.chanx_right_out_116_(sb_1__0__0_chanx_right_out_116_[0]),
		.chanx_right_out_118_(sb_1__0__0_chanx_right_out_118_[0]),
		.chanx_right_out_120_(sb_1__0__0_chanx_right_out_120_[0]),
		.chanx_right_out_122_(sb_1__0__0_chanx_right_out_122_[0]),
		.chanx_right_out_124_(sb_1__0__0_chanx_right_out_124_[0]),
		.chanx_right_out_126_(sb_1__0__0_chanx_right_out_126_[0]),
		.chanx_right_out_128_(sb_1__0__0_chanx_right_out_128_[0]),
		.chanx_right_out_130_(sb_1__0__0_chanx_right_out_130_[0]),
		.chanx_right_out_132_(sb_1__0__0_chanx_right_out_132_[0]),
		.chanx_right_out_134_(sb_1__0__0_chanx_right_out_134_[0]),
		.chanx_right_out_136_(sb_1__0__0_chanx_right_out_136_[0]),
		.chanx_right_out_138_(sb_1__0__0_chanx_right_out_138_[0]),
		.chanx_right_out_140_(sb_1__0__0_chanx_right_out_140_[0]),
		.chanx_right_out_142_(sb_1__0__0_chanx_right_out_142_[0]),
		.chanx_right_out_144_(sb_1__0__0_chanx_right_out_144_[0]),
		.chanx_right_out_146_(sb_1__0__0_chanx_right_out_146_[0]),
		.chanx_right_out_148_(sb_1__0__0_chanx_right_out_148_[0]),
		.chanx_right_out_150_(sb_1__0__0_chanx_right_out_150_[0]),
		.chanx_right_out_152_(sb_1__0__0_chanx_right_out_152_[0]),
		.chanx_right_out_154_(sb_1__0__0_chanx_right_out_154_[0]),
		.chanx_right_out_156_(sb_1__0__0_chanx_right_out_156_[0]),
		.chanx_right_out_158_(sb_1__0__0_chanx_right_out_158_[0]),
		.chanx_right_out_160_(sb_1__0__0_chanx_right_out_160_[0]),
		.chanx_right_out_162_(sb_1__0__0_chanx_right_out_162_[0]),
		.chanx_right_out_164_(sb_1__0__0_chanx_right_out_164_[0]),
		.chanx_right_out_166_(sb_1__0__0_chanx_right_out_166_[0]),
		.chanx_right_out_168_(sb_1__0__0_chanx_right_out_168_[0]),
		.chanx_right_out_170_(sb_1__0__0_chanx_right_out_170_[0]),
		.chanx_right_out_172_(sb_1__0__0_chanx_right_out_172_[0]),
		.chanx_right_out_174_(sb_1__0__0_chanx_right_out_174_[0]),
		.chanx_right_out_176_(sb_1__0__0_chanx_right_out_176_[0]),
		.chanx_right_out_178_(sb_1__0__0_chanx_right_out_178_[0]),
		.chanx_right_out_180_(sb_1__0__0_chanx_right_out_180_[0]),
		.chanx_right_out_182_(sb_1__0__0_chanx_right_out_182_[0]),
		.chanx_right_out_184_(sb_1__0__0_chanx_right_out_184_[0]),
		.chanx_right_out_186_(sb_1__0__0_chanx_right_out_186_[0]),
		.chanx_right_out_188_(sb_1__0__0_chanx_right_out_188_[0]),
		.chanx_right_out_190_(sb_1__0__0_chanx_right_out_190_[0]),
		.chanx_right_out_192_(sb_1__0__0_chanx_right_out_192_[0]),
		.chanx_right_out_194_(sb_1__0__0_chanx_right_out_194_[0]),
		.chanx_right_out_196_(sb_1__0__0_chanx_right_out_196_[0]),
		.chanx_right_out_198_(sb_1__0__0_chanx_right_out_198_[0]),
		.chanx_left_out_1_(sb_1__0__0_chanx_left_out_1_[0]),
		.chanx_left_out_3_(sb_1__0__0_chanx_left_out_3_[0]),
		.chanx_left_out_5_(sb_1__0__0_chanx_left_out_5_[0]),
		.chanx_left_out_7_(sb_1__0__0_chanx_left_out_7_[0]),
		.chanx_left_out_9_(sb_1__0__0_chanx_left_out_9_[0]),
		.chanx_left_out_11_(sb_1__0__0_chanx_left_out_11_[0]),
		.chanx_left_out_13_(sb_1__0__0_chanx_left_out_13_[0]),
		.chanx_left_out_15_(sb_1__0__0_chanx_left_out_15_[0]),
		.chanx_left_out_17_(sb_1__0__0_chanx_left_out_17_[0]),
		.chanx_left_out_19_(sb_1__0__0_chanx_left_out_19_[0]),
		.chanx_left_out_21_(sb_1__0__0_chanx_left_out_21_[0]),
		.chanx_left_out_23_(sb_1__0__0_chanx_left_out_23_[0]),
		.chanx_left_out_25_(sb_1__0__0_chanx_left_out_25_[0]),
		.chanx_left_out_27_(sb_1__0__0_chanx_left_out_27_[0]),
		.chanx_left_out_29_(sb_1__0__0_chanx_left_out_29_[0]),
		.chanx_left_out_31_(sb_1__0__0_chanx_left_out_31_[0]),
		.chanx_left_out_33_(sb_1__0__0_chanx_left_out_33_[0]),
		.chanx_left_out_35_(sb_1__0__0_chanx_left_out_35_[0]),
		.chanx_left_out_37_(sb_1__0__0_chanx_left_out_37_[0]),
		.chanx_left_out_39_(sb_1__0__0_chanx_left_out_39_[0]),
		.chanx_left_out_41_(sb_1__0__0_chanx_left_out_41_[0]),
		.chanx_left_out_43_(sb_1__0__0_chanx_left_out_43_[0]),
		.chanx_left_out_45_(sb_1__0__0_chanx_left_out_45_[0]),
		.chanx_left_out_47_(sb_1__0__0_chanx_left_out_47_[0]),
		.chanx_left_out_49_(sb_1__0__0_chanx_left_out_49_[0]),
		.chanx_left_out_51_(sb_1__0__0_chanx_left_out_51_[0]),
		.chanx_left_out_53_(sb_1__0__0_chanx_left_out_53_[0]),
		.chanx_left_out_55_(sb_1__0__0_chanx_left_out_55_[0]),
		.chanx_left_out_57_(sb_1__0__0_chanx_left_out_57_[0]),
		.chanx_left_out_59_(sb_1__0__0_chanx_left_out_59_[0]),
		.chanx_left_out_61_(sb_1__0__0_chanx_left_out_61_[0]),
		.chanx_left_out_63_(sb_1__0__0_chanx_left_out_63_[0]),
		.chanx_left_out_65_(sb_1__0__0_chanx_left_out_65_[0]),
		.chanx_left_out_67_(sb_1__0__0_chanx_left_out_67_[0]),
		.chanx_left_out_69_(sb_1__0__0_chanx_left_out_69_[0]),
		.chanx_left_out_71_(sb_1__0__0_chanx_left_out_71_[0]),
		.chanx_left_out_73_(sb_1__0__0_chanx_left_out_73_[0]),
		.chanx_left_out_75_(sb_1__0__0_chanx_left_out_75_[0]),
		.chanx_left_out_77_(sb_1__0__0_chanx_left_out_77_[0]),
		.chanx_left_out_79_(sb_1__0__0_chanx_left_out_79_[0]),
		.chanx_left_out_81_(sb_1__0__0_chanx_left_out_81_[0]),
		.chanx_left_out_83_(sb_1__0__0_chanx_left_out_83_[0]),
		.chanx_left_out_85_(sb_1__0__0_chanx_left_out_85_[0]),
		.chanx_left_out_87_(sb_1__0__0_chanx_left_out_87_[0]),
		.chanx_left_out_89_(sb_1__0__0_chanx_left_out_89_[0]),
		.chanx_left_out_91_(sb_1__0__0_chanx_left_out_91_[0]),
		.chanx_left_out_93_(sb_1__0__0_chanx_left_out_93_[0]),
		.chanx_left_out_95_(sb_1__0__0_chanx_left_out_95_[0]),
		.chanx_left_out_97_(sb_1__0__0_chanx_left_out_97_[0]),
		.chanx_left_out_99_(sb_1__0__0_chanx_left_out_99_[0]),
		.chanx_left_out_101_(sb_1__0__0_chanx_left_out_101_[0]),
		.chanx_left_out_103_(sb_1__0__0_chanx_left_out_103_[0]),
		.chanx_left_out_105_(sb_1__0__0_chanx_left_out_105_[0]),
		.chanx_left_out_107_(sb_1__0__0_chanx_left_out_107_[0]),
		.chanx_left_out_109_(sb_1__0__0_chanx_left_out_109_[0]),
		.chanx_left_out_111_(sb_1__0__0_chanx_left_out_111_[0]),
		.chanx_left_out_113_(sb_1__0__0_chanx_left_out_113_[0]),
		.chanx_left_out_115_(sb_1__0__0_chanx_left_out_115_[0]),
		.chanx_left_out_117_(sb_1__0__0_chanx_left_out_117_[0]),
		.chanx_left_out_119_(sb_1__0__0_chanx_left_out_119_[0]),
		.chanx_left_out_121_(sb_1__0__0_chanx_left_out_121_[0]),
		.chanx_left_out_123_(sb_1__0__0_chanx_left_out_123_[0]),
		.chanx_left_out_125_(sb_1__0__0_chanx_left_out_125_[0]),
		.chanx_left_out_127_(sb_1__0__0_chanx_left_out_127_[0]),
		.chanx_left_out_129_(sb_1__0__0_chanx_left_out_129_[0]),
		.chanx_left_out_131_(sb_1__0__0_chanx_left_out_131_[0]),
		.chanx_left_out_133_(sb_1__0__0_chanx_left_out_133_[0]),
		.chanx_left_out_135_(sb_1__0__0_chanx_left_out_135_[0]),
		.chanx_left_out_137_(sb_1__0__0_chanx_left_out_137_[0]),
		.chanx_left_out_139_(sb_1__0__0_chanx_left_out_139_[0]),
		.chanx_left_out_141_(sb_1__0__0_chanx_left_out_141_[0]),
		.chanx_left_out_143_(sb_1__0__0_chanx_left_out_143_[0]),
		.chanx_left_out_145_(sb_1__0__0_chanx_left_out_145_[0]),
		.chanx_left_out_147_(sb_1__0__0_chanx_left_out_147_[0]),
		.chanx_left_out_149_(sb_1__0__0_chanx_left_out_149_[0]),
		.chanx_left_out_151_(sb_1__0__0_chanx_left_out_151_[0]),
		.chanx_left_out_153_(sb_1__0__0_chanx_left_out_153_[0]),
		.chanx_left_out_155_(sb_1__0__0_chanx_left_out_155_[0]),
		.chanx_left_out_157_(sb_1__0__0_chanx_left_out_157_[0]),
		.chanx_left_out_159_(sb_1__0__0_chanx_left_out_159_[0]),
		.chanx_left_out_161_(sb_1__0__0_chanx_left_out_161_[0]),
		.chanx_left_out_163_(sb_1__0__0_chanx_left_out_163_[0]),
		.chanx_left_out_165_(sb_1__0__0_chanx_left_out_165_[0]),
		.chanx_left_out_167_(sb_1__0__0_chanx_left_out_167_[0]),
		.chanx_left_out_169_(sb_1__0__0_chanx_left_out_169_[0]),
		.chanx_left_out_171_(sb_1__0__0_chanx_left_out_171_[0]),
		.chanx_left_out_173_(sb_1__0__0_chanx_left_out_173_[0]),
		.chanx_left_out_175_(sb_1__0__0_chanx_left_out_175_[0]),
		.chanx_left_out_177_(sb_1__0__0_chanx_left_out_177_[0]),
		.chanx_left_out_179_(sb_1__0__0_chanx_left_out_179_[0]),
		.chanx_left_out_181_(sb_1__0__0_chanx_left_out_181_[0]),
		.chanx_left_out_183_(sb_1__0__0_chanx_left_out_183_[0]),
		.chanx_left_out_185_(sb_1__0__0_chanx_left_out_185_[0]),
		.chanx_left_out_187_(sb_1__0__0_chanx_left_out_187_[0]),
		.chanx_left_out_189_(sb_1__0__0_chanx_left_out_189_[0]),
		.chanx_left_out_191_(sb_1__0__0_chanx_left_out_191_[0]),
		.chanx_left_out_193_(sb_1__0__0_chanx_left_out_193_[0]),
		.chanx_left_out_195_(sb_1__0__0_chanx_left_out_195_[0]),
		.chanx_left_out_197_(sb_1__0__0_chanx_left_out_197_[0]),
		.chanx_left_out_199_(sb_1__0__0_chanx_left_out_199_[0]),
		.ccff_tail(sb_1__0__0_ccff_tail[0]));

	sb_1__1_ sb_1__1_ (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.chany_top_in_1_(cby_1__1__1_chany_out_1_[0]),
		.chany_top_in_3_(cby_1__1__1_chany_out_3_[0]),
		.chany_top_in_5_(cby_1__1__1_chany_out_5_[0]),
		.chany_top_in_7_(cby_1__1__1_chany_out_7_[0]),
		.chany_top_in_9_(cby_1__1__1_chany_out_9_[0]),
		.chany_top_in_11_(cby_1__1__1_chany_out_11_[0]),
		.chany_top_in_13_(cby_1__1__1_chany_out_13_[0]),
		.chany_top_in_15_(cby_1__1__1_chany_out_15_[0]),
		.chany_top_in_17_(cby_1__1__1_chany_out_17_[0]),
		.chany_top_in_19_(cby_1__1__1_chany_out_19_[0]),
		.chany_top_in_21_(cby_1__1__1_chany_out_21_[0]),
		.chany_top_in_23_(cby_1__1__1_chany_out_23_[0]),
		.chany_top_in_25_(cby_1__1__1_chany_out_25_[0]),
		.chany_top_in_27_(cby_1__1__1_chany_out_27_[0]),
		.chany_top_in_29_(cby_1__1__1_chany_out_29_[0]),
		.chany_top_in_31_(cby_1__1__1_chany_out_31_[0]),
		.chany_top_in_33_(cby_1__1__1_chany_out_33_[0]),
		.chany_top_in_35_(cby_1__1__1_chany_out_35_[0]),
		.chany_top_in_37_(cby_1__1__1_chany_out_37_[0]),
		.chany_top_in_39_(cby_1__1__1_chany_out_39_[0]),
		.chany_top_in_41_(cby_1__1__1_chany_out_41_[0]),
		.chany_top_in_43_(cby_1__1__1_chany_out_43_[0]),
		.chany_top_in_45_(cby_1__1__1_chany_out_45_[0]),
		.chany_top_in_47_(cby_1__1__1_chany_out_47_[0]),
		.chany_top_in_49_(cby_1__1__1_chany_out_49_[0]),
		.chany_top_in_51_(cby_1__1__1_chany_out_51_[0]),
		.chany_top_in_53_(cby_1__1__1_chany_out_53_[0]),
		.chany_top_in_55_(cby_1__1__1_chany_out_55_[0]),
		.chany_top_in_57_(cby_1__1__1_chany_out_57_[0]),
		.chany_top_in_59_(cby_1__1__1_chany_out_59_[0]),
		.chany_top_in_61_(cby_1__1__1_chany_out_61_[0]),
		.chany_top_in_63_(cby_1__1__1_chany_out_63_[0]),
		.chany_top_in_65_(cby_1__1__1_chany_out_65_[0]),
		.chany_top_in_67_(cby_1__1__1_chany_out_67_[0]),
		.chany_top_in_69_(cby_1__1__1_chany_out_69_[0]),
		.chany_top_in_71_(cby_1__1__1_chany_out_71_[0]),
		.chany_top_in_73_(cby_1__1__1_chany_out_73_[0]),
		.chany_top_in_75_(cby_1__1__1_chany_out_75_[0]),
		.chany_top_in_77_(cby_1__1__1_chany_out_77_[0]),
		.chany_top_in_79_(cby_1__1__1_chany_out_79_[0]),
		.chany_top_in_81_(cby_1__1__1_chany_out_81_[0]),
		.chany_top_in_83_(cby_1__1__1_chany_out_83_[0]),
		.chany_top_in_85_(cby_1__1__1_chany_out_85_[0]),
		.chany_top_in_87_(cby_1__1__1_chany_out_87_[0]),
		.chany_top_in_89_(cby_1__1__1_chany_out_89_[0]),
		.chany_top_in_91_(cby_1__1__1_chany_out_91_[0]),
		.chany_top_in_93_(cby_1__1__1_chany_out_93_[0]),
		.chany_top_in_95_(cby_1__1__1_chany_out_95_[0]),
		.chany_top_in_97_(cby_1__1__1_chany_out_97_[0]),
		.chany_top_in_99_(cby_1__1__1_chany_out_99_[0]),
		.chany_top_in_101_(cby_1__1__1_chany_out_101_[0]),
		.chany_top_in_103_(cby_1__1__1_chany_out_103_[0]),
		.chany_top_in_105_(cby_1__1__1_chany_out_105_[0]),
		.chany_top_in_107_(cby_1__1__1_chany_out_107_[0]),
		.chany_top_in_109_(cby_1__1__1_chany_out_109_[0]),
		.chany_top_in_111_(cby_1__1__1_chany_out_111_[0]),
		.chany_top_in_113_(cby_1__1__1_chany_out_113_[0]),
		.chany_top_in_115_(cby_1__1__1_chany_out_115_[0]),
		.chany_top_in_117_(cby_1__1__1_chany_out_117_[0]),
		.chany_top_in_119_(cby_1__1__1_chany_out_119_[0]),
		.chany_top_in_121_(cby_1__1__1_chany_out_121_[0]),
		.chany_top_in_123_(cby_1__1__1_chany_out_123_[0]),
		.chany_top_in_125_(cby_1__1__1_chany_out_125_[0]),
		.chany_top_in_127_(cby_1__1__1_chany_out_127_[0]),
		.chany_top_in_129_(cby_1__1__1_chany_out_129_[0]),
		.chany_top_in_131_(cby_1__1__1_chany_out_131_[0]),
		.chany_top_in_133_(cby_1__1__1_chany_out_133_[0]),
		.chany_top_in_135_(cby_1__1__1_chany_out_135_[0]),
		.chany_top_in_137_(cby_1__1__1_chany_out_137_[0]),
		.chany_top_in_139_(cby_1__1__1_chany_out_139_[0]),
		.chany_top_in_141_(cby_1__1__1_chany_out_141_[0]),
		.chany_top_in_143_(cby_1__1__1_chany_out_143_[0]),
		.chany_top_in_145_(cby_1__1__1_chany_out_145_[0]),
		.chany_top_in_147_(cby_1__1__1_chany_out_147_[0]),
		.chany_top_in_149_(cby_1__1__1_chany_out_149_[0]),
		.chany_top_in_151_(cby_1__1__1_chany_out_151_[0]),
		.chany_top_in_153_(cby_1__1__1_chany_out_153_[0]),
		.chany_top_in_155_(cby_1__1__1_chany_out_155_[0]),
		.chany_top_in_157_(cby_1__1__1_chany_out_157_[0]),
		.chany_top_in_159_(cby_1__1__1_chany_out_159_[0]),
		.chany_top_in_161_(cby_1__1__1_chany_out_161_[0]),
		.chany_top_in_163_(cby_1__1__1_chany_out_163_[0]),
		.chany_top_in_165_(cby_1__1__1_chany_out_165_[0]),
		.chany_top_in_167_(cby_1__1__1_chany_out_167_[0]),
		.chany_top_in_169_(cby_1__1__1_chany_out_169_[0]),
		.chany_top_in_171_(cby_1__1__1_chany_out_171_[0]),
		.chany_top_in_173_(cby_1__1__1_chany_out_173_[0]),
		.chany_top_in_175_(cby_1__1__1_chany_out_175_[0]),
		.chany_top_in_177_(cby_1__1__1_chany_out_177_[0]),
		.chany_top_in_179_(cby_1__1__1_chany_out_179_[0]),
		.chany_top_in_181_(cby_1__1__1_chany_out_181_[0]),
		.chany_top_in_183_(cby_1__1__1_chany_out_183_[0]),
		.chany_top_in_185_(cby_1__1__1_chany_out_185_[0]),
		.chany_top_in_187_(cby_1__1__1_chany_out_187_[0]),
		.chany_top_in_189_(cby_1__1__1_chany_out_189_[0]),
		.chany_top_in_191_(cby_1__1__1_chany_out_191_[0]),
		.chany_top_in_193_(cby_1__1__1_chany_out_193_[0]),
		.chany_top_in_195_(cby_1__1__1_chany_out_195_[0]),
		.chany_top_in_197_(cby_1__1__1_chany_out_197_[0]),
		.chany_top_in_199_(cby_1__1__1_chany_out_199_[0]),
		.top_left_grid_pin_44_(grid_clb_0_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_0_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_0_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_0_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_0_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_0_right_width_0_height_0__pin_49_lower[0]),
		.top_left_grid_pin_50_(grid_clb_0_right_width_0_height_0__pin_50_lower[0]),
		.top_left_grid_pin_51_(grid_clb_0_right_width_0_height_0__pin_51_lower[0]),
		.top_left_grid_pin_52_(grid_clb_0_right_width_0_height_0__pin_52_lower[0]),
		.top_left_grid_pin_53_(grid_clb_0_right_width_0_height_0__pin_53_lower[0]),
		.chanx_right_in_1_(cbx_1__1__1_chanx_out_1_[0]),
		.chanx_right_in_3_(cbx_1__1__1_chanx_out_3_[0]),
		.chanx_right_in_5_(cbx_1__1__1_chanx_out_5_[0]),
		.chanx_right_in_7_(cbx_1__1__1_chanx_out_7_[0]),
		.chanx_right_in_9_(cbx_1__1__1_chanx_out_9_[0]),
		.chanx_right_in_11_(cbx_1__1__1_chanx_out_11_[0]),
		.chanx_right_in_13_(cbx_1__1__1_chanx_out_13_[0]),
		.chanx_right_in_15_(cbx_1__1__1_chanx_out_15_[0]),
		.chanx_right_in_17_(cbx_1__1__1_chanx_out_17_[0]),
		.chanx_right_in_19_(cbx_1__1__1_chanx_out_19_[0]),
		.chanx_right_in_21_(cbx_1__1__1_chanx_out_21_[0]),
		.chanx_right_in_23_(cbx_1__1__1_chanx_out_23_[0]),
		.chanx_right_in_25_(cbx_1__1__1_chanx_out_25_[0]),
		.chanx_right_in_27_(cbx_1__1__1_chanx_out_27_[0]),
		.chanx_right_in_29_(cbx_1__1__1_chanx_out_29_[0]),
		.chanx_right_in_31_(cbx_1__1__1_chanx_out_31_[0]),
		.chanx_right_in_33_(cbx_1__1__1_chanx_out_33_[0]),
		.chanx_right_in_35_(cbx_1__1__1_chanx_out_35_[0]),
		.chanx_right_in_37_(cbx_1__1__1_chanx_out_37_[0]),
		.chanx_right_in_39_(cbx_1__1__1_chanx_out_39_[0]),
		.chanx_right_in_41_(cbx_1__1__1_chanx_out_41_[0]),
		.chanx_right_in_43_(cbx_1__1__1_chanx_out_43_[0]),
		.chanx_right_in_45_(cbx_1__1__1_chanx_out_45_[0]),
		.chanx_right_in_47_(cbx_1__1__1_chanx_out_47_[0]),
		.chanx_right_in_49_(cbx_1__1__1_chanx_out_49_[0]),
		.chanx_right_in_51_(cbx_1__1__1_chanx_out_51_[0]),
		.chanx_right_in_53_(cbx_1__1__1_chanx_out_53_[0]),
		.chanx_right_in_55_(cbx_1__1__1_chanx_out_55_[0]),
		.chanx_right_in_57_(cbx_1__1__1_chanx_out_57_[0]),
		.chanx_right_in_59_(cbx_1__1__1_chanx_out_59_[0]),
		.chanx_right_in_61_(cbx_1__1__1_chanx_out_61_[0]),
		.chanx_right_in_63_(cbx_1__1__1_chanx_out_63_[0]),
		.chanx_right_in_65_(cbx_1__1__1_chanx_out_65_[0]),
		.chanx_right_in_67_(cbx_1__1__1_chanx_out_67_[0]),
		.chanx_right_in_69_(cbx_1__1__1_chanx_out_69_[0]),
		.chanx_right_in_71_(cbx_1__1__1_chanx_out_71_[0]),
		.chanx_right_in_73_(cbx_1__1__1_chanx_out_73_[0]),
		.chanx_right_in_75_(cbx_1__1__1_chanx_out_75_[0]),
		.chanx_right_in_77_(cbx_1__1__1_chanx_out_77_[0]),
		.chanx_right_in_79_(cbx_1__1__1_chanx_out_79_[0]),
		.chanx_right_in_81_(cbx_1__1__1_chanx_out_81_[0]),
		.chanx_right_in_83_(cbx_1__1__1_chanx_out_83_[0]),
		.chanx_right_in_85_(cbx_1__1__1_chanx_out_85_[0]),
		.chanx_right_in_87_(cbx_1__1__1_chanx_out_87_[0]),
		.chanx_right_in_89_(cbx_1__1__1_chanx_out_89_[0]),
		.chanx_right_in_91_(cbx_1__1__1_chanx_out_91_[0]),
		.chanx_right_in_93_(cbx_1__1__1_chanx_out_93_[0]),
		.chanx_right_in_95_(cbx_1__1__1_chanx_out_95_[0]),
		.chanx_right_in_97_(cbx_1__1__1_chanx_out_97_[0]),
		.chanx_right_in_99_(cbx_1__1__1_chanx_out_99_[0]),
		.chanx_right_in_101_(cbx_1__1__1_chanx_out_101_[0]),
		.chanx_right_in_103_(cbx_1__1__1_chanx_out_103_[0]),
		.chanx_right_in_105_(cbx_1__1__1_chanx_out_105_[0]),
		.chanx_right_in_107_(cbx_1__1__1_chanx_out_107_[0]),
		.chanx_right_in_109_(cbx_1__1__1_chanx_out_109_[0]),
		.chanx_right_in_111_(cbx_1__1__1_chanx_out_111_[0]),
		.chanx_right_in_113_(cbx_1__1__1_chanx_out_113_[0]),
		.chanx_right_in_115_(cbx_1__1__1_chanx_out_115_[0]),
		.chanx_right_in_117_(cbx_1__1__1_chanx_out_117_[0]),
		.chanx_right_in_119_(cbx_1__1__1_chanx_out_119_[0]),
		.chanx_right_in_121_(cbx_1__1__1_chanx_out_121_[0]),
		.chanx_right_in_123_(cbx_1__1__1_chanx_out_123_[0]),
		.chanx_right_in_125_(cbx_1__1__1_chanx_out_125_[0]),
		.chanx_right_in_127_(cbx_1__1__1_chanx_out_127_[0]),
		.chanx_right_in_129_(cbx_1__1__1_chanx_out_129_[0]),
		.chanx_right_in_131_(cbx_1__1__1_chanx_out_131_[0]),
		.chanx_right_in_133_(cbx_1__1__1_chanx_out_133_[0]),
		.chanx_right_in_135_(cbx_1__1__1_chanx_out_135_[0]),
		.chanx_right_in_137_(cbx_1__1__1_chanx_out_137_[0]),
		.chanx_right_in_139_(cbx_1__1__1_chanx_out_139_[0]),
		.chanx_right_in_141_(cbx_1__1__1_chanx_out_141_[0]),
		.chanx_right_in_143_(cbx_1__1__1_chanx_out_143_[0]),
		.chanx_right_in_145_(cbx_1__1__1_chanx_out_145_[0]),
		.chanx_right_in_147_(cbx_1__1__1_chanx_out_147_[0]),
		.chanx_right_in_149_(cbx_1__1__1_chanx_out_149_[0]),
		.chanx_right_in_151_(cbx_1__1__1_chanx_out_151_[0]),
		.chanx_right_in_153_(cbx_1__1__1_chanx_out_153_[0]),
		.chanx_right_in_155_(cbx_1__1__1_chanx_out_155_[0]),
		.chanx_right_in_157_(cbx_1__1__1_chanx_out_157_[0]),
		.chanx_right_in_159_(cbx_1__1__1_chanx_out_159_[0]),
		.chanx_right_in_161_(cbx_1__1__1_chanx_out_161_[0]),
		.chanx_right_in_163_(cbx_1__1__1_chanx_out_163_[0]),
		.chanx_right_in_165_(cbx_1__1__1_chanx_out_165_[0]),
		.chanx_right_in_167_(cbx_1__1__1_chanx_out_167_[0]),
		.chanx_right_in_169_(cbx_1__1__1_chanx_out_169_[0]),
		.chanx_right_in_171_(cbx_1__1__1_chanx_out_171_[0]),
		.chanx_right_in_173_(cbx_1__1__1_chanx_out_173_[0]),
		.chanx_right_in_175_(cbx_1__1__1_chanx_out_175_[0]),
		.chanx_right_in_177_(cbx_1__1__1_chanx_out_177_[0]),
		.chanx_right_in_179_(cbx_1__1__1_chanx_out_179_[0]),
		.chanx_right_in_181_(cbx_1__1__1_chanx_out_181_[0]),
		.chanx_right_in_183_(cbx_1__1__1_chanx_out_183_[0]),
		.chanx_right_in_185_(cbx_1__1__1_chanx_out_185_[0]),
		.chanx_right_in_187_(cbx_1__1__1_chanx_out_187_[0]),
		.chanx_right_in_189_(cbx_1__1__1_chanx_out_189_[0]),
		.chanx_right_in_191_(cbx_1__1__1_chanx_out_191_[0]),
		.chanx_right_in_193_(cbx_1__1__1_chanx_out_193_[0]),
		.chanx_right_in_195_(cbx_1__1__1_chanx_out_195_[0]),
		.chanx_right_in_197_(cbx_1__1__1_chanx_out_197_[0]),
		.chanx_right_in_199_(cbx_1__1__1_chanx_out_199_[0]),
		.right_top_grid_pin_54_(grid_clb_2_bottom_width_0_height_0__pin_54_upper[0]),
		.right_top_grid_pin_55_(grid_clb_2_bottom_width_0_height_0__pin_55_upper[0]),
		.right_top_grid_pin_56_(grid_clb_2_bottom_width_0_height_0__pin_56_upper[0]),
		.right_top_grid_pin_57_(grid_clb_2_bottom_width_0_height_0__pin_57_upper[0]),
		.right_top_grid_pin_58_(grid_clb_2_bottom_width_0_height_0__pin_58_upper[0]),
		.right_top_grid_pin_59_(grid_clb_2_bottom_width_0_height_0__pin_59_upper[0]),
		.right_top_grid_pin_60_(grid_clb_2_bottom_width_0_height_0__pin_60_upper[0]),
		.right_top_grid_pin_61_(grid_clb_2_bottom_width_0_height_0__pin_61_upper[0]),
		.right_top_grid_pin_62_(grid_clb_2_bottom_width_0_height_0__pin_62_upper[0]),
		.right_top_grid_pin_63_(grid_clb_2_bottom_width_0_height_0__pin_63_upper[0]),
		.right_top_grid_pin_66_(grid_clb_2_bottom_width_0_height_0__pin_66_upper[0]),
		.right_top_grid_pin_67_(grid_clb_2_bottom_width_0_height_0__pin_67_upper[0]),
		.chany_bottom_in_0_(cby_1__1__0_chany_out_0_[0]),
		.chany_bottom_in_2_(cby_1__1__0_chany_out_2_[0]),
		.chany_bottom_in_4_(cby_1__1__0_chany_out_4_[0]),
		.chany_bottom_in_6_(cby_1__1__0_chany_out_6_[0]),
		.chany_bottom_in_8_(cby_1__1__0_chany_out_8_[0]),
		.chany_bottom_in_10_(cby_1__1__0_chany_out_10_[0]),
		.chany_bottom_in_12_(cby_1__1__0_chany_out_12_[0]),
		.chany_bottom_in_14_(cby_1__1__0_chany_out_14_[0]),
		.chany_bottom_in_16_(cby_1__1__0_chany_out_16_[0]),
		.chany_bottom_in_18_(cby_1__1__0_chany_out_18_[0]),
		.chany_bottom_in_20_(cby_1__1__0_chany_out_20_[0]),
		.chany_bottom_in_22_(cby_1__1__0_chany_out_22_[0]),
		.chany_bottom_in_24_(cby_1__1__0_chany_out_24_[0]),
		.chany_bottom_in_26_(cby_1__1__0_chany_out_26_[0]),
		.chany_bottom_in_28_(cby_1__1__0_chany_out_28_[0]),
		.chany_bottom_in_30_(cby_1__1__0_chany_out_30_[0]),
		.chany_bottom_in_32_(cby_1__1__0_chany_out_32_[0]),
		.chany_bottom_in_34_(cby_1__1__0_chany_out_34_[0]),
		.chany_bottom_in_36_(cby_1__1__0_chany_out_36_[0]),
		.chany_bottom_in_38_(cby_1__1__0_chany_out_38_[0]),
		.chany_bottom_in_40_(cby_1__1__0_chany_out_40_[0]),
		.chany_bottom_in_42_(cby_1__1__0_chany_out_42_[0]),
		.chany_bottom_in_44_(cby_1__1__0_chany_out_44_[0]),
		.chany_bottom_in_46_(cby_1__1__0_chany_out_46_[0]),
		.chany_bottom_in_48_(cby_1__1__0_chany_out_48_[0]),
		.chany_bottom_in_50_(cby_1__1__0_chany_out_50_[0]),
		.chany_bottom_in_52_(cby_1__1__0_chany_out_52_[0]),
		.chany_bottom_in_54_(cby_1__1__0_chany_out_54_[0]),
		.chany_bottom_in_56_(cby_1__1__0_chany_out_56_[0]),
		.chany_bottom_in_58_(cby_1__1__0_chany_out_58_[0]),
		.chany_bottom_in_60_(cby_1__1__0_chany_out_60_[0]),
		.chany_bottom_in_62_(cby_1__1__0_chany_out_62_[0]),
		.chany_bottom_in_64_(cby_1__1__0_chany_out_64_[0]),
		.chany_bottom_in_66_(cby_1__1__0_chany_out_66_[0]),
		.chany_bottom_in_68_(cby_1__1__0_chany_out_68_[0]),
		.chany_bottom_in_70_(cby_1__1__0_chany_out_70_[0]),
		.chany_bottom_in_72_(cby_1__1__0_chany_out_72_[0]),
		.chany_bottom_in_74_(cby_1__1__0_chany_out_74_[0]),
		.chany_bottom_in_76_(cby_1__1__0_chany_out_76_[0]),
		.chany_bottom_in_78_(cby_1__1__0_chany_out_78_[0]),
		.chany_bottom_in_80_(cby_1__1__0_chany_out_80_[0]),
		.chany_bottom_in_82_(cby_1__1__0_chany_out_82_[0]),
		.chany_bottom_in_84_(cby_1__1__0_chany_out_84_[0]),
		.chany_bottom_in_86_(cby_1__1__0_chany_out_86_[0]),
		.chany_bottom_in_88_(cby_1__1__0_chany_out_88_[0]),
		.chany_bottom_in_90_(cby_1__1__0_chany_out_90_[0]),
		.chany_bottom_in_92_(cby_1__1__0_chany_out_92_[0]),
		.chany_bottom_in_94_(cby_1__1__0_chany_out_94_[0]),
		.chany_bottom_in_96_(cby_1__1__0_chany_out_96_[0]),
		.chany_bottom_in_98_(cby_1__1__0_chany_out_98_[0]),
		.chany_bottom_in_100_(cby_1__1__0_chany_out_100_[0]),
		.chany_bottom_in_102_(cby_1__1__0_chany_out_102_[0]),
		.chany_bottom_in_104_(cby_1__1__0_chany_out_104_[0]),
		.chany_bottom_in_106_(cby_1__1__0_chany_out_106_[0]),
		.chany_bottom_in_108_(cby_1__1__0_chany_out_108_[0]),
		.chany_bottom_in_110_(cby_1__1__0_chany_out_110_[0]),
		.chany_bottom_in_112_(cby_1__1__0_chany_out_112_[0]),
		.chany_bottom_in_114_(cby_1__1__0_chany_out_114_[0]),
		.chany_bottom_in_116_(cby_1__1__0_chany_out_116_[0]),
		.chany_bottom_in_118_(cby_1__1__0_chany_out_118_[0]),
		.chany_bottom_in_120_(cby_1__1__0_chany_out_120_[0]),
		.chany_bottom_in_122_(cby_1__1__0_chany_out_122_[0]),
		.chany_bottom_in_124_(cby_1__1__0_chany_out_124_[0]),
		.chany_bottom_in_126_(cby_1__1__0_chany_out_126_[0]),
		.chany_bottom_in_128_(cby_1__1__0_chany_out_128_[0]),
		.chany_bottom_in_130_(cby_1__1__0_chany_out_130_[0]),
		.chany_bottom_in_132_(cby_1__1__0_chany_out_132_[0]),
		.chany_bottom_in_134_(cby_1__1__0_chany_out_134_[0]),
		.chany_bottom_in_136_(cby_1__1__0_chany_out_136_[0]),
		.chany_bottom_in_138_(cby_1__1__0_chany_out_138_[0]),
		.chany_bottom_in_140_(cby_1__1__0_chany_out_140_[0]),
		.chany_bottom_in_142_(cby_1__1__0_chany_out_142_[0]),
		.chany_bottom_in_144_(cby_1__1__0_chany_out_144_[0]),
		.chany_bottom_in_146_(cby_1__1__0_chany_out_146_[0]),
		.chany_bottom_in_148_(cby_1__1__0_chany_out_148_[0]),
		.chany_bottom_in_150_(cby_1__1__0_chany_out_150_[0]),
		.chany_bottom_in_152_(cby_1__1__0_chany_out_152_[0]),
		.chany_bottom_in_154_(cby_1__1__0_chany_out_154_[0]),
		.chany_bottom_in_156_(cby_1__1__0_chany_out_156_[0]),
		.chany_bottom_in_158_(cby_1__1__0_chany_out_158_[0]),
		.chany_bottom_in_160_(cby_1__1__0_chany_out_160_[0]),
		.chany_bottom_in_162_(cby_1__1__0_chany_out_162_[0]),
		.chany_bottom_in_164_(cby_1__1__0_chany_out_164_[0]),
		.chany_bottom_in_166_(cby_1__1__0_chany_out_166_[0]),
		.chany_bottom_in_168_(cby_1__1__0_chany_out_168_[0]),
		.chany_bottom_in_170_(cby_1__1__0_chany_out_170_[0]),
		.chany_bottom_in_172_(cby_1__1__0_chany_out_172_[0]),
		.chany_bottom_in_174_(cby_1__1__0_chany_out_174_[0]),
		.chany_bottom_in_176_(cby_1__1__0_chany_out_176_[0]),
		.chany_bottom_in_178_(cby_1__1__0_chany_out_178_[0]),
		.chany_bottom_in_180_(cby_1__1__0_chany_out_180_[0]),
		.chany_bottom_in_182_(cby_1__1__0_chany_out_182_[0]),
		.chany_bottom_in_184_(cby_1__1__0_chany_out_184_[0]),
		.chany_bottom_in_186_(cby_1__1__0_chany_out_186_[0]),
		.chany_bottom_in_188_(cby_1__1__0_chany_out_188_[0]),
		.chany_bottom_in_190_(cby_1__1__0_chany_out_190_[0]),
		.chany_bottom_in_192_(cby_1__1__0_chany_out_192_[0]),
		.chany_bottom_in_194_(cby_1__1__0_chany_out_194_[0]),
		.chany_bottom_in_196_(cby_1__1__0_chany_out_196_[0]),
		.chany_bottom_in_198_(cby_1__1__0_chany_out_198_[0]),
		.bottom_left_grid_pin_44_(grid_clb_spypad_0_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_spypad_0_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_spypad_0_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_spypad_0_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_spypad_0_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_spypad_0_right_width_0_height_0__pin_49_upper[0]),
		.bottom_left_grid_pin_50_(grid_clb_spypad_0_right_width_0_height_0__pin_50_upper[0]),
		.bottom_left_grid_pin_51_(grid_clb_spypad_0_right_width_0_height_0__pin_51_upper[0]),
		.bottom_left_grid_pin_52_(grid_clb_spypad_0_right_width_0_height_0__pin_52_upper[0]),
		.bottom_left_grid_pin_53_(grid_clb_spypad_0_right_width_0_height_0__pin_53_upper[0]),
		.chanx_left_in_0_(cbx_1__1__0_chanx_out_0_[0]),
		.chanx_left_in_2_(cbx_1__1__0_chanx_out_2_[0]),
		.chanx_left_in_4_(cbx_1__1__0_chanx_out_4_[0]),
		.chanx_left_in_6_(cbx_1__1__0_chanx_out_6_[0]),
		.chanx_left_in_8_(cbx_1__1__0_chanx_out_8_[0]),
		.chanx_left_in_10_(cbx_1__1__0_chanx_out_10_[0]),
		.chanx_left_in_12_(cbx_1__1__0_chanx_out_12_[0]),
		.chanx_left_in_14_(cbx_1__1__0_chanx_out_14_[0]),
		.chanx_left_in_16_(cbx_1__1__0_chanx_out_16_[0]),
		.chanx_left_in_18_(cbx_1__1__0_chanx_out_18_[0]),
		.chanx_left_in_20_(cbx_1__1__0_chanx_out_20_[0]),
		.chanx_left_in_22_(cbx_1__1__0_chanx_out_22_[0]),
		.chanx_left_in_24_(cbx_1__1__0_chanx_out_24_[0]),
		.chanx_left_in_26_(cbx_1__1__0_chanx_out_26_[0]),
		.chanx_left_in_28_(cbx_1__1__0_chanx_out_28_[0]),
		.chanx_left_in_30_(cbx_1__1__0_chanx_out_30_[0]),
		.chanx_left_in_32_(cbx_1__1__0_chanx_out_32_[0]),
		.chanx_left_in_34_(cbx_1__1__0_chanx_out_34_[0]),
		.chanx_left_in_36_(cbx_1__1__0_chanx_out_36_[0]),
		.chanx_left_in_38_(cbx_1__1__0_chanx_out_38_[0]),
		.chanx_left_in_40_(cbx_1__1__0_chanx_out_40_[0]),
		.chanx_left_in_42_(cbx_1__1__0_chanx_out_42_[0]),
		.chanx_left_in_44_(cbx_1__1__0_chanx_out_44_[0]),
		.chanx_left_in_46_(cbx_1__1__0_chanx_out_46_[0]),
		.chanx_left_in_48_(cbx_1__1__0_chanx_out_48_[0]),
		.chanx_left_in_50_(cbx_1__1__0_chanx_out_50_[0]),
		.chanx_left_in_52_(cbx_1__1__0_chanx_out_52_[0]),
		.chanx_left_in_54_(cbx_1__1__0_chanx_out_54_[0]),
		.chanx_left_in_56_(cbx_1__1__0_chanx_out_56_[0]),
		.chanx_left_in_58_(cbx_1__1__0_chanx_out_58_[0]),
		.chanx_left_in_60_(cbx_1__1__0_chanx_out_60_[0]),
		.chanx_left_in_62_(cbx_1__1__0_chanx_out_62_[0]),
		.chanx_left_in_64_(cbx_1__1__0_chanx_out_64_[0]),
		.chanx_left_in_66_(cbx_1__1__0_chanx_out_66_[0]),
		.chanx_left_in_68_(cbx_1__1__0_chanx_out_68_[0]),
		.chanx_left_in_70_(cbx_1__1__0_chanx_out_70_[0]),
		.chanx_left_in_72_(cbx_1__1__0_chanx_out_72_[0]),
		.chanx_left_in_74_(cbx_1__1__0_chanx_out_74_[0]),
		.chanx_left_in_76_(cbx_1__1__0_chanx_out_76_[0]),
		.chanx_left_in_78_(cbx_1__1__0_chanx_out_78_[0]),
		.chanx_left_in_80_(cbx_1__1__0_chanx_out_80_[0]),
		.chanx_left_in_82_(cbx_1__1__0_chanx_out_82_[0]),
		.chanx_left_in_84_(cbx_1__1__0_chanx_out_84_[0]),
		.chanx_left_in_86_(cbx_1__1__0_chanx_out_86_[0]),
		.chanx_left_in_88_(cbx_1__1__0_chanx_out_88_[0]),
		.chanx_left_in_90_(cbx_1__1__0_chanx_out_90_[0]),
		.chanx_left_in_92_(cbx_1__1__0_chanx_out_92_[0]),
		.chanx_left_in_94_(cbx_1__1__0_chanx_out_94_[0]),
		.chanx_left_in_96_(cbx_1__1__0_chanx_out_96_[0]),
		.chanx_left_in_98_(cbx_1__1__0_chanx_out_98_[0]),
		.chanx_left_in_100_(cbx_1__1__0_chanx_out_100_[0]),
		.chanx_left_in_102_(cbx_1__1__0_chanx_out_102_[0]),
		.chanx_left_in_104_(cbx_1__1__0_chanx_out_104_[0]),
		.chanx_left_in_106_(cbx_1__1__0_chanx_out_106_[0]),
		.chanx_left_in_108_(cbx_1__1__0_chanx_out_108_[0]),
		.chanx_left_in_110_(cbx_1__1__0_chanx_out_110_[0]),
		.chanx_left_in_112_(cbx_1__1__0_chanx_out_112_[0]),
		.chanx_left_in_114_(cbx_1__1__0_chanx_out_114_[0]),
		.chanx_left_in_116_(cbx_1__1__0_chanx_out_116_[0]),
		.chanx_left_in_118_(cbx_1__1__0_chanx_out_118_[0]),
		.chanx_left_in_120_(cbx_1__1__0_chanx_out_120_[0]),
		.chanx_left_in_122_(cbx_1__1__0_chanx_out_122_[0]),
		.chanx_left_in_124_(cbx_1__1__0_chanx_out_124_[0]),
		.chanx_left_in_126_(cbx_1__1__0_chanx_out_126_[0]),
		.chanx_left_in_128_(cbx_1__1__0_chanx_out_128_[0]),
		.chanx_left_in_130_(cbx_1__1__0_chanx_out_130_[0]),
		.chanx_left_in_132_(cbx_1__1__0_chanx_out_132_[0]),
		.chanx_left_in_134_(cbx_1__1__0_chanx_out_134_[0]),
		.chanx_left_in_136_(cbx_1__1__0_chanx_out_136_[0]),
		.chanx_left_in_138_(cbx_1__1__0_chanx_out_138_[0]),
		.chanx_left_in_140_(cbx_1__1__0_chanx_out_140_[0]),
		.chanx_left_in_142_(cbx_1__1__0_chanx_out_142_[0]),
		.chanx_left_in_144_(cbx_1__1__0_chanx_out_144_[0]),
		.chanx_left_in_146_(cbx_1__1__0_chanx_out_146_[0]),
		.chanx_left_in_148_(cbx_1__1__0_chanx_out_148_[0]),
		.chanx_left_in_150_(cbx_1__1__0_chanx_out_150_[0]),
		.chanx_left_in_152_(cbx_1__1__0_chanx_out_152_[0]),
		.chanx_left_in_154_(cbx_1__1__0_chanx_out_154_[0]),
		.chanx_left_in_156_(cbx_1__1__0_chanx_out_156_[0]),
		.chanx_left_in_158_(cbx_1__1__0_chanx_out_158_[0]),
		.chanx_left_in_160_(cbx_1__1__0_chanx_out_160_[0]),
		.chanx_left_in_162_(cbx_1__1__0_chanx_out_162_[0]),
		.chanx_left_in_164_(cbx_1__1__0_chanx_out_164_[0]),
		.chanx_left_in_166_(cbx_1__1__0_chanx_out_166_[0]),
		.chanx_left_in_168_(cbx_1__1__0_chanx_out_168_[0]),
		.chanx_left_in_170_(cbx_1__1__0_chanx_out_170_[0]),
		.chanx_left_in_172_(cbx_1__1__0_chanx_out_172_[0]),
		.chanx_left_in_174_(cbx_1__1__0_chanx_out_174_[0]),
		.chanx_left_in_176_(cbx_1__1__0_chanx_out_176_[0]),
		.chanx_left_in_178_(cbx_1__1__0_chanx_out_178_[0]),
		.chanx_left_in_180_(cbx_1__1__0_chanx_out_180_[0]),
		.chanx_left_in_182_(cbx_1__1__0_chanx_out_182_[0]),
		.chanx_left_in_184_(cbx_1__1__0_chanx_out_184_[0]),
		.chanx_left_in_186_(cbx_1__1__0_chanx_out_186_[0]),
		.chanx_left_in_188_(cbx_1__1__0_chanx_out_188_[0]),
		.chanx_left_in_190_(cbx_1__1__0_chanx_out_190_[0]),
		.chanx_left_in_192_(cbx_1__1__0_chanx_out_192_[0]),
		.chanx_left_in_194_(cbx_1__1__0_chanx_out_194_[0]),
		.chanx_left_in_196_(cbx_1__1__0_chanx_out_196_[0]),
		.chanx_left_in_198_(cbx_1__1__0_chanx_out_198_[0]),
		.left_top_grid_pin_54_(grid_clb_0_bottom_width_0_height_0__pin_54_lower[0]),
		.left_top_grid_pin_55_(grid_clb_0_bottom_width_0_height_0__pin_55_lower[0]),
		.left_top_grid_pin_56_(grid_clb_0_bottom_width_0_height_0__pin_56_lower[0]),
		.left_top_grid_pin_57_(grid_clb_0_bottom_width_0_height_0__pin_57_lower[0]),
		.left_top_grid_pin_58_(grid_clb_0_bottom_width_0_height_0__pin_58_lower[0]),
		.left_top_grid_pin_59_(grid_clb_0_bottom_width_0_height_0__pin_59_lower[0]),
		.left_top_grid_pin_60_(grid_clb_0_bottom_width_0_height_0__pin_60_lower[0]),
		.left_top_grid_pin_61_(grid_clb_0_bottom_width_0_height_0__pin_61_lower[0]),
		.left_top_grid_pin_62_(grid_clb_0_bottom_width_0_height_0__pin_62_lower[0]),
		.left_top_grid_pin_63_(grid_clb_0_bottom_width_0_height_0__pin_63_lower[0]),
		.left_top_grid_pin_66_(grid_clb_0_bottom_width_0_height_0__pin_66_lower[0]),
		.left_top_grid_pin_67_(grid_clb_0_bottom_width_0_height_0__pin_67_lower[0]),
		.ccff_head(grid_clb_2_ccff_tail[0]),
		.chany_top_out_0_(sb_1__1__0_chany_top_out_0_[0]),
		.chany_top_out_2_(sb_1__1__0_chany_top_out_2_[0]),
		.chany_top_out_4_(sb_1__1__0_chany_top_out_4_[0]),
		.chany_top_out_6_(sb_1__1__0_chany_top_out_6_[0]),
		.chany_top_out_8_(sb_1__1__0_chany_top_out_8_[0]),
		.chany_top_out_10_(sb_1__1__0_chany_top_out_10_[0]),
		.chany_top_out_12_(sb_1__1__0_chany_top_out_12_[0]),
		.chany_top_out_14_(sb_1__1__0_chany_top_out_14_[0]),
		.chany_top_out_16_(sb_1__1__0_chany_top_out_16_[0]),
		.chany_top_out_18_(sb_1__1__0_chany_top_out_18_[0]),
		.chany_top_out_20_(sb_1__1__0_chany_top_out_20_[0]),
		.chany_top_out_22_(sb_1__1__0_chany_top_out_22_[0]),
		.chany_top_out_24_(sb_1__1__0_chany_top_out_24_[0]),
		.chany_top_out_26_(sb_1__1__0_chany_top_out_26_[0]),
		.chany_top_out_28_(sb_1__1__0_chany_top_out_28_[0]),
		.chany_top_out_30_(sb_1__1__0_chany_top_out_30_[0]),
		.chany_top_out_32_(sb_1__1__0_chany_top_out_32_[0]),
		.chany_top_out_34_(sb_1__1__0_chany_top_out_34_[0]),
		.chany_top_out_36_(sb_1__1__0_chany_top_out_36_[0]),
		.chany_top_out_38_(sb_1__1__0_chany_top_out_38_[0]),
		.chany_top_out_40_(sb_1__1__0_chany_top_out_40_[0]),
		.chany_top_out_42_(sb_1__1__0_chany_top_out_42_[0]),
		.chany_top_out_44_(sb_1__1__0_chany_top_out_44_[0]),
		.chany_top_out_46_(sb_1__1__0_chany_top_out_46_[0]),
		.chany_top_out_48_(sb_1__1__0_chany_top_out_48_[0]),
		.chany_top_out_50_(sb_1__1__0_chany_top_out_50_[0]),
		.chany_top_out_52_(sb_1__1__0_chany_top_out_52_[0]),
		.chany_top_out_54_(sb_1__1__0_chany_top_out_54_[0]),
		.chany_top_out_56_(sb_1__1__0_chany_top_out_56_[0]),
		.chany_top_out_58_(sb_1__1__0_chany_top_out_58_[0]),
		.chany_top_out_60_(sb_1__1__0_chany_top_out_60_[0]),
		.chany_top_out_62_(sb_1__1__0_chany_top_out_62_[0]),
		.chany_top_out_64_(sb_1__1__0_chany_top_out_64_[0]),
		.chany_top_out_66_(sb_1__1__0_chany_top_out_66_[0]),
		.chany_top_out_68_(sb_1__1__0_chany_top_out_68_[0]),
		.chany_top_out_70_(sb_1__1__0_chany_top_out_70_[0]),
		.chany_top_out_72_(sb_1__1__0_chany_top_out_72_[0]),
		.chany_top_out_74_(sb_1__1__0_chany_top_out_74_[0]),
		.chany_top_out_76_(sb_1__1__0_chany_top_out_76_[0]),
		.chany_top_out_78_(sb_1__1__0_chany_top_out_78_[0]),
		.chany_top_out_80_(sb_1__1__0_chany_top_out_80_[0]),
		.chany_top_out_82_(sb_1__1__0_chany_top_out_82_[0]),
		.chany_top_out_84_(sb_1__1__0_chany_top_out_84_[0]),
		.chany_top_out_86_(sb_1__1__0_chany_top_out_86_[0]),
		.chany_top_out_88_(sb_1__1__0_chany_top_out_88_[0]),
		.chany_top_out_90_(sb_1__1__0_chany_top_out_90_[0]),
		.chany_top_out_92_(sb_1__1__0_chany_top_out_92_[0]),
		.chany_top_out_94_(sb_1__1__0_chany_top_out_94_[0]),
		.chany_top_out_96_(sb_1__1__0_chany_top_out_96_[0]),
		.chany_top_out_98_(sb_1__1__0_chany_top_out_98_[0]),
		.chany_top_out_100_(sb_1__1__0_chany_top_out_100_[0]),
		.chany_top_out_102_(sb_1__1__0_chany_top_out_102_[0]),
		.chany_top_out_104_(sb_1__1__0_chany_top_out_104_[0]),
		.chany_top_out_106_(sb_1__1__0_chany_top_out_106_[0]),
		.chany_top_out_108_(sb_1__1__0_chany_top_out_108_[0]),
		.chany_top_out_110_(sb_1__1__0_chany_top_out_110_[0]),
		.chany_top_out_112_(sb_1__1__0_chany_top_out_112_[0]),
		.chany_top_out_114_(sb_1__1__0_chany_top_out_114_[0]),
		.chany_top_out_116_(sb_1__1__0_chany_top_out_116_[0]),
		.chany_top_out_118_(sb_1__1__0_chany_top_out_118_[0]),
		.chany_top_out_120_(sb_1__1__0_chany_top_out_120_[0]),
		.chany_top_out_122_(sb_1__1__0_chany_top_out_122_[0]),
		.chany_top_out_124_(sb_1__1__0_chany_top_out_124_[0]),
		.chany_top_out_126_(sb_1__1__0_chany_top_out_126_[0]),
		.chany_top_out_128_(sb_1__1__0_chany_top_out_128_[0]),
		.chany_top_out_130_(sb_1__1__0_chany_top_out_130_[0]),
		.chany_top_out_132_(sb_1__1__0_chany_top_out_132_[0]),
		.chany_top_out_134_(sb_1__1__0_chany_top_out_134_[0]),
		.chany_top_out_136_(sb_1__1__0_chany_top_out_136_[0]),
		.chany_top_out_138_(sb_1__1__0_chany_top_out_138_[0]),
		.chany_top_out_140_(sb_1__1__0_chany_top_out_140_[0]),
		.chany_top_out_142_(sb_1__1__0_chany_top_out_142_[0]),
		.chany_top_out_144_(sb_1__1__0_chany_top_out_144_[0]),
		.chany_top_out_146_(sb_1__1__0_chany_top_out_146_[0]),
		.chany_top_out_148_(sb_1__1__0_chany_top_out_148_[0]),
		.chany_top_out_150_(sb_1__1__0_chany_top_out_150_[0]),
		.chany_top_out_152_(sb_1__1__0_chany_top_out_152_[0]),
		.chany_top_out_154_(sb_1__1__0_chany_top_out_154_[0]),
		.chany_top_out_156_(sb_1__1__0_chany_top_out_156_[0]),
		.chany_top_out_158_(sb_1__1__0_chany_top_out_158_[0]),
		.chany_top_out_160_(sb_1__1__0_chany_top_out_160_[0]),
		.chany_top_out_162_(sb_1__1__0_chany_top_out_162_[0]),
		.chany_top_out_164_(sb_1__1__0_chany_top_out_164_[0]),
		.chany_top_out_166_(sb_1__1__0_chany_top_out_166_[0]),
		.chany_top_out_168_(sb_1__1__0_chany_top_out_168_[0]),
		.chany_top_out_170_(sb_1__1__0_chany_top_out_170_[0]),
		.chany_top_out_172_(sb_1__1__0_chany_top_out_172_[0]),
		.chany_top_out_174_(sb_1__1__0_chany_top_out_174_[0]),
		.chany_top_out_176_(sb_1__1__0_chany_top_out_176_[0]),
		.chany_top_out_178_(sb_1__1__0_chany_top_out_178_[0]),
		.chany_top_out_180_(sb_1__1__0_chany_top_out_180_[0]),
		.chany_top_out_182_(sb_1__1__0_chany_top_out_182_[0]),
		.chany_top_out_184_(sb_1__1__0_chany_top_out_184_[0]),
		.chany_top_out_186_(sb_1__1__0_chany_top_out_186_[0]),
		.chany_top_out_188_(sb_1__1__0_chany_top_out_188_[0]),
		.chany_top_out_190_(sb_1__1__0_chany_top_out_190_[0]),
		.chany_top_out_192_(sb_1__1__0_chany_top_out_192_[0]),
		.chany_top_out_194_(sb_1__1__0_chany_top_out_194_[0]),
		.chany_top_out_196_(sb_1__1__0_chany_top_out_196_[0]),
		.chany_top_out_198_(sb_1__1__0_chany_top_out_198_[0]),
		.chanx_right_out_0_(sb_1__1__0_chanx_right_out_0_[0]),
		.chanx_right_out_2_(sb_1__1__0_chanx_right_out_2_[0]),
		.chanx_right_out_4_(sb_1__1__0_chanx_right_out_4_[0]),
		.chanx_right_out_6_(sb_1__1__0_chanx_right_out_6_[0]),
		.chanx_right_out_8_(sb_1__1__0_chanx_right_out_8_[0]),
		.chanx_right_out_10_(sb_1__1__0_chanx_right_out_10_[0]),
		.chanx_right_out_12_(sb_1__1__0_chanx_right_out_12_[0]),
		.chanx_right_out_14_(sb_1__1__0_chanx_right_out_14_[0]),
		.chanx_right_out_16_(sb_1__1__0_chanx_right_out_16_[0]),
		.chanx_right_out_18_(sb_1__1__0_chanx_right_out_18_[0]),
		.chanx_right_out_20_(sb_1__1__0_chanx_right_out_20_[0]),
		.chanx_right_out_22_(sb_1__1__0_chanx_right_out_22_[0]),
		.chanx_right_out_24_(sb_1__1__0_chanx_right_out_24_[0]),
		.chanx_right_out_26_(sb_1__1__0_chanx_right_out_26_[0]),
		.chanx_right_out_28_(sb_1__1__0_chanx_right_out_28_[0]),
		.chanx_right_out_30_(sb_1__1__0_chanx_right_out_30_[0]),
		.chanx_right_out_32_(sb_1__1__0_chanx_right_out_32_[0]),
		.chanx_right_out_34_(sb_1__1__0_chanx_right_out_34_[0]),
		.chanx_right_out_36_(sb_1__1__0_chanx_right_out_36_[0]),
		.chanx_right_out_38_(sb_1__1__0_chanx_right_out_38_[0]),
		.chanx_right_out_40_(sb_1__1__0_chanx_right_out_40_[0]),
		.chanx_right_out_42_(sb_1__1__0_chanx_right_out_42_[0]),
		.chanx_right_out_44_(sb_1__1__0_chanx_right_out_44_[0]),
		.chanx_right_out_46_(sb_1__1__0_chanx_right_out_46_[0]),
		.chanx_right_out_48_(sb_1__1__0_chanx_right_out_48_[0]),
		.chanx_right_out_50_(sb_1__1__0_chanx_right_out_50_[0]),
		.chanx_right_out_52_(sb_1__1__0_chanx_right_out_52_[0]),
		.chanx_right_out_54_(sb_1__1__0_chanx_right_out_54_[0]),
		.chanx_right_out_56_(sb_1__1__0_chanx_right_out_56_[0]),
		.chanx_right_out_58_(sb_1__1__0_chanx_right_out_58_[0]),
		.chanx_right_out_60_(sb_1__1__0_chanx_right_out_60_[0]),
		.chanx_right_out_62_(sb_1__1__0_chanx_right_out_62_[0]),
		.chanx_right_out_64_(sb_1__1__0_chanx_right_out_64_[0]),
		.chanx_right_out_66_(sb_1__1__0_chanx_right_out_66_[0]),
		.chanx_right_out_68_(sb_1__1__0_chanx_right_out_68_[0]),
		.chanx_right_out_70_(sb_1__1__0_chanx_right_out_70_[0]),
		.chanx_right_out_72_(sb_1__1__0_chanx_right_out_72_[0]),
		.chanx_right_out_74_(sb_1__1__0_chanx_right_out_74_[0]),
		.chanx_right_out_76_(sb_1__1__0_chanx_right_out_76_[0]),
		.chanx_right_out_78_(sb_1__1__0_chanx_right_out_78_[0]),
		.chanx_right_out_80_(sb_1__1__0_chanx_right_out_80_[0]),
		.chanx_right_out_82_(sb_1__1__0_chanx_right_out_82_[0]),
		.chanx_right_out_84_(sb_1__1__0_chanx_right_out_84_[0]),
		.chanx_right_out_86_(sb_1__1__0_chanx_right_out_86_[0]),
		.chanx_right_out_88_(sb_1__1__0_chanx_right_out_88_[0]),
		.chanx_right_out_90_(sb_1__1__0_chanx_right_out_90_[0]),
		.chanx_right_out_92_(sb_1__1__0_chanx_right_out_92_[0]),
		.chanx_right_out_94_(sb_1__1__0_chanx_right_out_94_[0]),
		.chanx_right_out_96_(sb_1__1__0_chanx_right_out_96_[0]),
		.chanx_right_out_98_(sb_1__1__0_chanx_right_out_98_[0]),
		.chanx_right_out_100_(sb_1__1__0_chanx_right_out_100_[0]),
		.chanx_right_out_102_(sb_1__1__0_chanx_right_out_102_[0]),
		.chanx_right_out_104_(sb_1__1__0_chanx_right_out_104_[0]),
		.chanx_right_out_106_(sb_1__1__0_chanx_right_out_106_[0]),
		.chanx_right_out_108_(sb_1__1__0_chanx_right_out_108_[0]),
		.chanx_right_out_110_(sb_1__1__0_chanx_right_out_110_[0]),
		.chanx_right_out_112_(sb_1__1__0_chanx_right_out_112_[0]),
		.chanx_right_out_114_(sb_1__1__0_chanx_right_out_114_[0]),
		.chanx_right_out_116_(sb_1__1__0_chanx_right_out_116_[0]),
		.chanx_right_out_118_(sb_1__1__0_chanx_right_out_118_[0]),
		.chanx_right_out_120_(sb_1__1__0_chanx_right_out_120_[0]),
		.chanx_right_out_122_(sb_1__1__0_chanx_right_out_122_[0]),
		.chanx_right_out_124_(sb_1__1__0_chanx_right_out_124_[0]),
		.chanx_right_out_126_(sb_1__1__0_chanx_right_out_126_[0]),
		.chanx_right_out_128_(sb_1__1__0_chanx_right_out_128_[0]),
		.chanx_right_out_130_(sb_1__1__0_chanx_right_out_130_[0]),
		.chanx_right_out_132_(sb_1__1__0_chanx_right_out_132_[0]),
		.chanx_right_out_134_(sb_1__1__0_chanx_right_out_134_[0]),
		.chanx_right_out_136_(sb_1__1__0_chanx_right_out_136_[0]),
		.chanx_right_out_138_(sb_1__1__0_chanx_right_out_138_[0]),
		.chanx_right_out_140_(sb_1__1__0_chanx_right_out_140_[0]),
		.chanx_right_out_142_(sb_1__1__0_chanx_right_out_142_[0]),
		.chanx_right_out_144_(sb_1__1__0_chanx_right_out_144_[0]),
		.chanx_right_out_146_(sb_1__1__0_chanx_right_out_146_[0]),
		.chanx_right_out_148_(sb_1__1__0_chanx_right_out_148_[0]),
		.chanx_right_out_150_(sb_1__1__0_chanx_right_out_150_[0]),
		.chanx_right_out_152_(sb_1__1__0_chanx_right_out_152_[0]),
		.chanx_right_out_154_(sb_1__1__0_chanx_right_out_154_[0]),
		.chanx_right_out_156_(sb_1__1__0_chanx_right_out_156_[0]),
		.chanx_right_out_158_(sb_1__1__0_chanx_right_out_158_[0]),
		.chanx_right_out_160_(sb_1__1__0_chanx_right_out_160_[0]),
		.chanx_right_out_162_(sb_1__1__0_chanx_right_out_162_[0]),
		.chanx_right_out_164_(sb_1__1__0_chanx_right_out_164_[0]),
		.chanx_right_out_166_(sb_1__1__0_chanx_right_out_166_[0]),
		.chanx_right_out_168_(sb_1__1__0_chanx_right_out_168_[0]),
		.chanx_right_out_170_(sb_1__1__0_chanx_right_out_170_[0]),
		.chanx_right_out_172_(sb_1__1__0_chanx_right_out_172_[0]),
		.chanx_right_out_174_(sb_1__1__0_chanx_right_out_174_[0]),
		.chanx_right_out_176_(sb_1__1__0_chanx_right_out_176_[0]),
		.chanx_right_out_178_(sb_1__1__0_chanx_right_out_178_[0]),
		.chanx_right_out_180_(sb_1__1__0_chanx_right_out_180_[0]),
		.chanx_right_out_182_(sb_1__1__0_chanx_right_out_182_[0]),
		.chanx_right_out_184_(sb_1__1__0_chanx_right_out_184_[0]),
		.chanx_right_out_186_(sb_1__1__0_chanx_right_out_186_[0]),
		.chanx_right_out_188_(sb_1__1__0_chanx_right_out_188_[0]),
		.chanx_right_out_190_(sb_1__1__0_chanx_right_out_190_[0]),
		.chanx_right_out_192_(sb_1__1__0_chanx_right_out_192_[0]),
		.chanx_right_out_194_(sb_1__1__0_chanx_right_out_194_[0]),
		.chanx_right_out_196_(sb_1__1__0_chanx_right_out_196_[0]),
		.chanx_right_out_198_(sb_1__1__0_chanx_right_out_198_[0]),
		.chany_bottom_out_1_(sb_1__1__0_chany_bottom_out_1_[0]),
		.chany_bottom_out_3_(sb_1__1__0_chany_bottom_out_3_[0]),
		.chany_bottom_out_5_(sb_1__1__0_chany_bottom_out_5_[0]),
		.chany_bottom_out_7_(sb_1__1__0_chany_bottom_out_7_[0]),
		.chany_bottom_out_9_(sb_1__1__0_chany_bottom_out_9_[0]),
		.chany_bottom_out_11_(sb_1__1__0_chany_bottom_out_11_[0]),
		.chany_bottom_out_13_(sb_1__1__0_chany_bottom_out_13_[0]),
		.chany_bottom_out_15_(sb_1__1__0_chany_bottom_out_15_[0]),
		.chany_bottom_out_17_(sb_1__1__0_chany_bottom_out_17_[0]),
		.chany_bottom_out_19_(sb_1__1__0_chany_bottom_out_19_[0]),
		.chany_bottom_out_21_(sb_1__1__0_chany_bottom_out_21_[0]),
		.chany_bottom_out_23_(sb_1__1__0_chany_bottom_out_23_[0]),
		.chany_bottom_out_25_(sb_1__1__0_chany_bottom_out_25_[0]),
		.chany_bottom_out_27_(sb_1__1__0_chany_bottom_out_27_[0]),
		.chany_bottom_out_29_(sb_1__1__0_chany_bottom_out_29_[0]),
		.chany_bottom_out_31_(sb_1__1__0_chany_bottom_out_31_[0]),
		.chany_bottom_out_33_(sb_1__1__0_chany_bottom_out_33_[0]),
		.chany_bottom_out_35_(sb_1__1__0_chany_bottom_out_35_[0]),
		.chany_bottom_out_37_(sb_1__1__0_chany_bottom_out_37_[0]),
		.chany_bottom_out_39_(sb_1__1__0_chany_bottom_out_39_[0]),
		.chany_bottom_out_41_(sb_1__1__0_chany_bottom_out_41_[0]),
		.chany_bottom_out_43_(sb_1__1__0_chany_bottom_out_43_[0]),
		.chany_bottom_out_45_(sb_1__1__0_chany_bottom_out_45_[0]),
		.chany_bottom_out_47_(sb_1__1__0_chany_bottom_out_47_[0]),
		.chany_bottom_out_49_(sb_1__1__0_chany_bottom_out_49_[0]),
		.chany_bottom_out_51_(sb_1__1__0_chany_bottom_out_51_[0]),
		.chany_bottom_out_53_(sb_1__1__0_chany_bottom_out_53_[0]),
		.chany_bottom_out_55_(sb_1__1__0_chany_bottom_out_55_[0]),
		.chany_bottom_out_57_(sb_1__1__0_chany_bottom_out_57_[0]),
		.chany_bottom_out_59_(sb_1__1__0_chany_bottom_out_59_[0]),
		.chany_bottom_out_61_(sb_1__1__0_chany_bottom_out_61_[0]),
		.chany_bottom_out_63_(sb_1__1__0_chany_bottom_out_63_[0]),
		.chany_bottom_out_65_(sb_1__1__0_chany_bottom_out_65_[0]),
		.chany_bottom_out_67_(sb_1__1__0_chany_bottom_out_67_[0]),
		.chany_bottom_out_69_(sb_1__1__0_chany_bottom_out_69_[0]),
		.chany_bottom_out_71_(sb_1__1__0_chany_bottom_out_71_[0]),
		.chany_bottom_out_73_(sb_1__1__0_chany_bottom_out_73_[0]),
		.chany_bottom_out_75_(sb_1__1__0_chany_bottom_out_75_[0]),
		.chany_bottom_out_77_(sb_1__1__0_chany_bottom_out_77_[0]),
		.chany_bottom_out_79_(sb_1__1__0_chany_bottom_out_79_[0]),
		.chany_bottom_out_81_(sb_1__1__0_chany_bottom_out_81_[0]),
		.chany_bottom_out_83_(sb_1__1__0_chany_bottom_out_83_[0]),
		.chany_bottom_out_85_(sb_1__1__0_chany_bottom_out_85_[0]),
		.chany_bottom_out_87_(sb_1__1__0_chany_bottom_out_87_[0]),
		.chany_bottom_out_89_(sb_1__1__0_chany_bottom_out_89_[0]),
		.chany_bottom_out_91_(sb_1__1__0_chany_bottom_out_91_[0]),
		.chany_bottom_out_93_(sb_1__1__0_chany_bottom_out_93_[0]),
		.chany_bottom_out_95_(sb_1__1__0_chany_bottom_out_95_[0]),
		.chany_bottom_out_97_(sb_1__1__0_chany_bottom_out_97_[0]),
		.chany_bottom_out_99_(sb_1__1__0_chany_bottom_out_99_[0]),
		.chany_bottom_out_101_(sb_1__1__0_chany_bottom_out_101_[0]),
		.chany_bottom_out_103_(sb_1__1__0_chany_bottom_out_103_[0]),
		.chany_bottom_out_105_(sb_1__1__0_chany_bottom_out_105_[0]),
		.chany_bottom_out_107_(sb_1__1__0_chany_bottom_out_107_[0]),
		.chany_bottom_out_109_(sb_1__1__0_chany_bottom_out_109_[0]),
		.chany_bottom_out_111_(sb_1__1__0_chany_bottom_out_111_[0]),
		.chany_bottom_out_113_(sb_1__1__0_chany_bottom_out_113_[0]),
		.chany_bottom_out_115_(sb_1__1__0_chany_bottom_out_115_[0]),
		.chany_bottom_out_117_(sb_1__1__0_chany_bottom_out_117_[0]),
		.chany_bottom_out_119_(sb_1__1__0_chany_bottom_out_119_[0]),
		.chany_bottom_out_121_(sb_1__1__0_chany_bottom_out_121_[0]),
		.chany_bottom_out_123_(sb_1__1__0_chany_bottom_out_123_[0]),
		.chany_bottom_out_125_(sb_1__1__0_chany_bottom_out_125_[0]),
		.chany_bottom_out_127_(sb_1__1__0_chany_bottom_out_127_[0]),
		.chany_bottom_out_129_(sb_1__1__0_chany_bottom_out_129_[0]),
		.chany_bottom_out_131_(sb_1__1__0_chany_bottom_out_131_[0]),
		.chany_bottom_out_133_(sb_1__1__0_chany_bottom_out_133_[0]),
		.chany_bottom_out_135_(sb_1__1__0_chany_bottom_out_135_[0]),
		.chany_bottom_out_137_(sb_1__1__0_chany_bottom_out_137_[0]),
		.chany_bottom_out_139_(sb_1__1__0_chany_bottom_out_139_[0]),
		.chany_bottom_out_141_(sb_1__1__0_chany_bottom_out_141_[0]),
		.chany_bottom_out_143_(sb_1__1__0_chany_bottom_out_143_[0]),
		.chany_bottom_out_145_(sb_1__1__0_chany_bottom_out_145_[0]),
		.chany_bottom_out_147_(sb_1__1__0_chany_bottom_out_147_[0]),
		.chany_bottom_out_149_(sb_1__1__0_chany_bottom_out_149_[0]),
		.chany_bottom_out_151_(sb_1__1__0_chany_bottom_out_151_[0]),
		.chany_bottom_out_153_(sb_1__1__0_chany_bottom_out_153_[0]),
		.chany_bottom_out_155_(sb_1__1__0_chany_bottom_out_155_[0]),
		.chany_bottom_out_157_(sb_1__1__0_chany_bottom_out_157_[0]),
		.chany_bottom_out_159_(sb_1__1__0_chany_bottom_out_159_[0]),
		.chany_bottom_out_161_(sb_1__1__0_chany_bottom_out_161_[0]),
		.chany_bottom_out_163_(sb_1__1__0_chany_bottom_out_163_[0]),
		.chany_bottom_out_165_(sb_1__1__0_chany_bottom_out_165_[0]),
		.chany_bottom_out_167_(sb_1__1__0_chany_bottom_out_167_[0]),
		.chany_bottom_out_169_(sb_1__1__0_chany_bottom_out_169_[0]),
		.chany_bottom_out_171_(sb_1__1__0_chany_bottom_out_171_[0]),
		.chany_bottom_out_173_(sb_1__1__0_chany_bottom_out_173_[0]),
		.chany_bottom_out_175_(sb_1__1__0_chany_bottom_out_175_[0]),
		.chany_bottom_out_177_(sb_1__1__0_chany_bottom_out_177_[0]),
		.chany_bottom_out_179_(sb_1__1__0_chany_bottom_out_179_[0]),
		.chany_bottom_out_181_(sb_1__1__0_chany_bottom_out_181_[0]),
		.chany_bottom_out_183_(sb_1__1__0_chany_bottom_out_183_[0]),
		.chany_bottom_out_185_(sb_1__1__0_chany_bottom_out_185_[0]),
		.chany_bottom_out_187_(sb_1__1__0_chany_bottom_out_187_[0]),
		.chany_bottom_out_189_(sb_1__1__0_chany_bottom_out_189_[0]),
		.chany_bottom_out_191_(sb_1__1__0_chany_bottom_out_191_[0]),
		.chany_bottom_out_193_(sb_1__1__0_chany_bottom_out_193_[0]),
		.chany_bottom_out_195_(sb_1__1__0_chany_bottom_out_195_[0]),
		.chany_bottom_out_197_(sb_1__1__0_chany_bottom_out_197_[0]),
		.chany_bottom_out_199_(sb_1__1__0_chany_bottom_out_199_[0]),
		.chanx_left_out_1_(sb_1__1__0_chanx_left_out_1_[0]),
		.chanx_left_out_3_(sb_1__1__0_chanx_left_out_3_[0]),
		.chanx_left_out_5_(sb_1__1__0_chanx_left_out_5_[0]),
		.chanx_left_out_7_(sb_1__1__0_chanx_left_out_7_[0]),
		.chanx_left_out_9_(sb_1__1__0_chanx_left_out_9_[0]),
		.chanx_left_out_11_(sb_1__1__0_chanx_left_out_11_[0]),
		.chanx_left_out_13_(sb_1__1__0_chanx_left_out_13_[0]),
		.chanx_left_out_15_(sb_1__1__0_chanx_left_out_15_[0]),
		.chanx_left_out_17_(sb_1__1__0_chanx_left_out_17_[0]),
		.chanx_left_out_19_(sb_1__1__0_chanx_left_out_19_[0]),
		.chanx_left_out_21_(sb_1__1__0_chanx_left_out_21_[0]),
		.chanx_left_out_23_(sb_1__1__0_chanx_left_out_23_[0]),
		.chanx_left_out_25_(sb_1__1__0_chanx_left_out_25_[0]),
		.chanx_left_out_27_(sb_1__1__0_chanx_left_out_27_[0]),
		.chanx_left_out_29_(sb_1__1__0_chanx_left_out_29_[0]),
		.chanx_left_out_31_(sb_1__1__0_chanx_left_out_31_[0]),
		.chanx_left_out_33_(sb_1__1__0_chanx_left_out_33_[0]),
		.chanx_left_out_35_(sb_1__1__0_chanx_left_out_35_[0]),
		.chanx_left_out_37_(sb_1__1__0_chanx_left_out_37_[0]),
		.chanx_left_out_39_(sb_1__1__0_chanx_left_out_39_[0]),
		.chanx_left_out_41_(sb_1__1__0_chanx_left_out_41_[0]),
		.chanx_left_out_43_(sb_1__1__0_chanx_left_out_43_[0]),
		.chanx_left_out_45_(sb_1__1__0_chanx_left_out_45_[0]),
		.chanx_left_out_47_(sb_1__1__0_chanx_left_out_47_[0]),
		.chanx_left_out_49_(sb_1__1__0_chanx_left_out_49_[0]),
		.chanx_left_out_51_(sb_1__1__0_chanx_left_out_51_[0]),
		.chanx_left_out_53_(sb_1__1__0_chanx_left_out_53_[0]),
		.chanx_left_out_55_(sb_1__1__0_chanx_left_out_55_[0]),
		.chanx_left_out_57_(sb_1__1__0_chanx_left_out_57_[0]),
		.chanx_left_out_59_(sb_1__1__0_chanx_left_out_59_[0]),
		.chanx_left_out_61_(sb_1__1__0_chanx_left_out_61_[0]),
		.chanx_left_out_63_(sb_1__1__0_chanx_left_out_63_[0]),
		.chanx_left_out_65_(sb_1__1__0_chanx_left_out_65_[0]),
		.chanx_left_out_67_(sb_1__1__0_chanx_left_out_67_[0]),
		.chanx_left_out_69_(sb_1__1__0_chanx_left_out_69_[0]),
		.chanx_left_out_71_(sb_1__1__0_chanx_left_out_71_[0]),
		.chanx_left_out_73_(sb_1__1__0_chanx_left_out_73_[0]),
		.chanx_left_out_75_(sb_1__1__0_chanx_left_out_75_[0]),
		.chanx_left_out_77_(sb_1__1__0_chanx_left_out_77_[0]),
		.chanx_left_out_79_(sb_1__1__0_chanx_left_out_79_[0]),
		.chanx_left_out_81_(sb_1__1__0_chanx_left_out_81_[0]),
		.chanx_left_out_83_(sb_1__1__0_chanx_left_out_83_[0]),
		.chanx_left_out_85_(sb_1__1__0_chanx_left_out_85_[0]),
		.chanx_left_out_87_(sb_1__1__0_chanx_left_out_87_[0]),
		.chanx_left_out_89_(sb_1__1__0_chanx_left_out_89_[0]),
		.chanx_left_out_91_(sb_1__1__0_chanx_left_out_91_[0]),
		.chanx_left_out_93_(sb_1__1__0_chanx_left_out_93_[0]),
		.chanx_left_out_95_(sb_1__1__0_chanx_left_out_95_[0]),
		.chanx_left_out_97_(sb_1__1__0_chanx_left_out_97_[0]),
		.chanx_left_out_99_(sb_1__1__0_chanx_left_out_99_[0]),
		.chanx_left_out_101_(sb_1__1__0_chanx_left_out_101_[0]),
		.chanx_left_out_103_(sb_1__1__0_chanx_left_out_103_[0]),
		.chanx_left_out_105_(sb_1__1__0_chanx_left_out_105_[0]),
		.chanx_left_out_107_(sb_1__1__0_chanx_left_out_107_[0]),
		.chanx_left_out_109_(sb_1__1__0_chanx_left_out_109_[0]),
		.chanx_left_out_111_(sb_1__1__0_chanx_left_out_111_[0]),
		.chanx_left_out_113_(sb_1__1__0_chanx_left_out_113_[0]),
		.chanx_left_out_115_(sb_1__1__0_chanx_left_out_115_[0]),
		.chanx_left_out_117_(sb_1__1__0_chanx_left_out_117_[0]),
		.chanx_left_out_119_(sb_1__1__0_chanx_left_out_119_[0]),
		.chanx_left_out_121_(sb_1__1__0_chanx_left_out_121_[0]),
		.chanx_left_out_123_(sb_1__1__0_chanx_left_out_123_[0]),
		.chanx_left_out_125_(sb_1__1__0_chanx_left_out_125_[0]),
		.chanx_left_out_127_(sb_1__1__0_chanx_left_out_127_[0]),
		.chanx_left_out_129_(sb_1__1__0_chanx_left_out_129_[0]),
		.chanx_left_out_131_(sb_1__1__0_chanx_left_out_131_[0]),
		.chanx_left_out_133_(sb_1__1__0_chanx_left_out_133_[0]),
		.chanx_left_out_135_(sb_1__1__0_chanx_left_out_135_[0]),
		.chanx_left_out_137_(sb_1__1__0_chanx_left_out_137_[0]),
		.chanx_left_out_139_(sb_1__1__0_chanx_left_out_139_[0]),
		.chanx_left_out_141_(sb_1__1__0_chanx_left_out_141_[0]),
		.chanx_left_out_143_(sb_1__1__0_chanx_left_out_143_[0]),
		.chanx_left_out_145_(sb_1__1__0_chanx_left_out_145_[0]),
		.chanx_left_out_147_(sb_1__1__0_chanx_left_out_147_[0]),
		.chanx_left_out_149_(sb_1__1__0_chanx_left_out_149_[0]),
		.chanx_left_out_151_(sb_1__1__0_chanx_left_out_151_[0]),
		.chanx_left_out_153_(sb_1__1__0_chanx_left_out_153_[0]),
		.chanx_left_out_155_(sb_1__1__0_chanx_left_out_155_[0]),
		.chanx_left_out_157_(sb_1__1__0_chanx_left_out_157_[0]),
		.chanx_left_out_159_(sb_1__1__0_chanx_left_out_159_[0]),
		.chanx_left_out_161_(sb_1__1__0_chanx_left_out_161_[0]),
		.chanx_left_out_163_(sb_1__1__0_chanx_left_out_163_[0]),
		.chanx_left_out_165_(sb_1__1__0_chanx_left_out_165_[0]),
		.chanx_left_out_167_(sb_1__1__0_chanx_left_out_167_[0]),
		.chanx_left_out_169_(sb_1__1__0_chanx_left_out_169_[0]),
		.chanx_left_out_171_(sb_1__1__0_chanx_left_out_171_[0]),
		.chanx_left_out_173_(sb_1__1__0_chanx_left_out_173_[0]),
		.chanx_left_out_175_(sb_1__1__0_chanx_left_out_175_[0]),
		.chanx_left_out_177_(sb_1__1__0_chanx_left_out_177_[0]),
		.chanx_left_out_179_(sb_1__1__0_chanx_left_out_179_[0]),
		.chanx_left_out_181_(sb_1__1__0_chanx_left_out_181_[0]),
		.chanx_left_out_183_(sb_1__1__0_chanx_left_out_183_[0]),
		.chanx_left_out_185_(sb_1__1__0_chanx_left_out_185_[0]),
		.chanx_left_out_187_(sb_1__1__0_chanx_left_out_187_[0]),
		.chanx_left_out_189_(sb_1__1__0_chanx_left_out_189_[0]),
		.chanx_left_out_191_(sb_1__1__0_chanx_left_out_191_[0]),
		.chanx_left_out_193_(sb_1__1__0_chanx_left_out_193_[0]),
		.chanx_left_out_195_(sb_1__1__0_chanx_left_out_195_[0]),
		.chanx_left_out_197_(sb_1__1__0_chanx_left_out_197_[0]),
		.chanx_left_out_199_(sb_1__1__0_chanx_left_out_199_[0]),
		.ccff_tail(sb_1__1__0_ccff_tail[0]));

	sb_1__2_ sb_1__2_ (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.chanx_right_in_1_(cbx_1__2__1_chanx_out_1_[0]),
		.chanx_right_in_3_(cbx_1__2__1_chanx_out_3_[0]),
		.chanx_right_in_5_(cbx_1__2__1_chanx_out_5_[0]),
		.chanx_right_in_7_(cbx_1__2__1_chanx_out_7_[0]),
		.chanx_right_in_9_(cbx_1__2__1_chanx_out_9_[0]),
		.chanx_right_in_11_(cbx_1__2__1_chanx_out_11_[0]),
		.chanx_right_in_13_(cbx_1__2__1_chanx_out_13_[0]),
		.chanx_right_in_15_(cbx_1__2__1_chanx_out_15_[0]),
		.chanx_right_in_17_(cbx_1__2__1_chanx_out_17_[0]),
		.chanx_right_in_19_(cbx_1__2__1_chanx_out_19_[0]),
		.chanx_right_in_21_(cbx_1__2__1_chanx_out_21_[0]),
		.chanx_right_in_23_(cbx_1__2__1_chanx_out_23_[0]),
		.chanx_right_in_25_(cbx_1__2__1_chanx_out_25_[0]),
		.chanx_right_in_27_(cbx_1__2__1_chanx_out_27_[0]),
		.chanx_right_in_29_(cbx_1__2__1_chanx_out_29_[0]),
		.chanx_right_in_31_(cbx_1__2__1_chanx_out_31_[0]),
		.chanx_right_in_33_(cbx_1__2__1_chanx_out_33_[0]),
		.chanx_right_in_35_(cbx_1__2__1_chanx_out_35_[0]),
		.chanx_right_in_37_(cbx_1__2__1_chanx_out_37_[0]),
		.chanx_right_in_39_(cbx_1__2__1_chanx_out_39_[0]),
		.chanx_right_in_41_(cbx_1__2__1_chanx_out_41_[0]),
		.chanx_right_in_43_(cbx_1__2__1_chanx_out_43_[0]),
		.chanx_right_in_45_(cbx_1__2__1_chanx_out_45_[0]),
		.chanx_right_in_47_(cbx_1__2__1_chanx_out_47_[0]),
		.chanx_right_in_49_(cbx_1__2__1_chanx_out_49_[0]),
		.chanx_right_in_51_(cbx_1__2__1_chanx_out_51_[0]),
		.chanx_right_in_53_(cbx_1__2__1_chanx_out_53_[0]),
		.chanx_right_in_55_(cbx_1__2__1_chanx_out_55_[0]),
		.chanx_right_in_57_(cbx_1__2__1_chanx_out_57_[0]),
		.chanx_right_in_59_(cbx_1__2__1_chanx_out_59_[0]),
		.chanx_right_in_61_(cbx_1__2__1_chanx_out_61_[0]),
		.chanx_right_in_63_(cbx_1__2__1_chanx_out_63_[0]),
		.chanx_right_in_65_(cbx_1__2__1_chanx_out_65_[0]),
		.chanx_right_in_67_(cbx_1__2__1_chanx_out_67_[0]),
		.chanx_right_in_69_(cbx_1__2__1_chanx_out_69_[0]),
		.chanx_right_in_71_(cbx_1__2__1_chanx_out_71_[0]),
		.chanx_right_in_73_(cbx_1__2__1_chanx_out_73_[0]),
		.chanx_right_in_75_(cbx_1__2__1_chanx_out_75_[0]),
		.chanx_right_in_77_(cbx_1__2__1_chanx_out_77_[0]),
		.chanx_right_in_79_(cbx_1__2__1_chanx_out_79_[0]),
		.chanx_right_in_81_(cbx_1__2__1_chanx_out_81_[0]),
		.chanx_right_in_83_(cbx_1__2__1_chanx_out_83_[0]),
		.chanx_right_in_85_(cbx_1__2__1_chanx_out_85_[0]),
		.chanx_right_in_87_(cbx_1__2__1_chanx_out_87_[0]),
		.chanx_right_in_89_(cbx_1__2__1_chanx_out_89_[0]),
		.chanx_right_in_91_(cbx_1__2__1_chanx_out_91_[0]),
		.chanx_right_in_93_(cbx_1__2__1_chanx_out_93_[0]),
		.chanx_right_in_95_(cbx_1__2__1_chanx_out_95_[0]),
		.chanx_right_in_97_(cbx_1__2__1_chanx_out_97_[0]),
		.chanx_right_in_99_(cbx_1__2__1_chanx_out_99_[0]),
		.chanx_right_in_101_(cbx_1__2__1_chanx_out_101_[0]),
		.chanx_right_in_103_(cbx_1__2__1_chanx_out_103_[0]),
		.chanx_right_in_105_(cbx_1__2__1_chanx_out_105_[0]),
		.chanx_right_in_107_(cbx_1__2__1_chanx_out_107_[0]),
		.chanx_right_in_109_(cbx_1__2__1_chanx_out_109_[0]),
		.chanx_right_in_111_(cbx_1__2__1_chanx_out_111_[0]),
		.chanx_right_in_113_(cbx_1__2__1_chanx_out_113_[0]),
		.chanx_right_in_115_(cbx_1__2__1_chanx_out_115_[0]),
		.chanx_right_in_117_(cbx_1__2__1_chanx_out_117_[0]),
		.chanx_right_in_119_(cbx_1__2__1_chanx_out_119_[0]),
		.chanx_right_in_121_(cbx_1__2__1_chanx_out_121_[0]),
		.chanx_right_in_123_(cbx_1__2__1_chanx_out_123_[0]),
		.chanx_right_in_125_(cbx_1__2__1_chanx_out_125_[0]),
		.chanx_right_in_127_(cbx_1__2__1_chanx_out_127_[0]),
		.chanx_right_in_129_(cbx_1__2__1_chanx_out_129_[0]),
		.chanx_right_in_131_(cbx_1__2__1_chanx_out_131_[0]),
		.chanx_right_in_133_(cbx_1__2__1_chanx_out_133_[0]),
		.chanx_right_in_135_(cbx_1__2__1_chanx_out_135_[0]),
		.chanx_right_in_137_(cbx_1__2__1_chanx_out_137_[0]),
		.chanx_right_in_139_(cbx_1__2__1_chanx_out_139_[0]),
		.chanx_right_in_141_(cbx_1__2__1_chanx_out_141_[0]),
		.chanx_right_in_143_(cbx_1__2__1_chanx_out_143_[0]),
		.chanx_right_in_145_(cbx_1__2__1_chanx_out_145_[0]),
		.chanx_right_in_147_(cbx_1__2__1_chanx_out_147_[0]),
		.chanx_right_in_149_(cbx_1__2__1_chanx_out_149_[0]),
		.chanx_right_in_151_(cbx_1__2__1_chanx_out_151_[0]),
		.chanx_right_in_153_(cbx_1__2__1_chanx_out_153_[0]),
		.chanx_right_in_155_(cbx_1__2__1_chanx_out_155_[0]),
		.chanx_right_in_157_(cbx_1__2__1_chanx_out_157_[0]),
		.chanx_right_in_159_(cbx_1__2__1_chanx_out_159_[0]),
		.chanx_right_in_161_(cbx_1__2__1_chanx_out_161_[0]),
		.chanx_right_in_163_(cbx_1__2__1_chanx_out_163_[0]),
		.chanx_right_in_165_(cbx_1__2__1_chanx_out_165_[0]),
		.chanx_right_in_167_(cbx_1__2__1_chanx_out_167_[0]),
		.chanx_right_in_169_(cbx_1__2__1_chanx_out_169_[0]),
		.chanx_right_in_171_(cbx_1__2__1_chanx_out_171_[0]),
		.chanx_right_in_173_(cbx_1__2__1_chanx_out_173_[0]),
		.chanx_right_in_175_(cbx_1__2__1_chanx_out_175_[0]),
		.chanx_right_in_177_(cbx_1__2__1_chanx_out_177_[0]),
		.chanx_right_in_179_(cbx_1__2__1_chanx_out_179_[0]),
		.chanx_right_in_181_(cbx_1__2__1_chanx_out_181_[0]),
		.chanx_right_in_183_(cbx_1__2__1_chanx_out_183_[0]),
		.chanx_right_in_185_(cbx_1__2__1_chanx_out_185_[0]),
		.chanx_right_in_187_(cbx_1__2__1_chanx_out_187_[0]),
		.chanx_right_in_189_(cbx_1__2__1_chanx_out_189_[0]),
		.chanx_right_in_191_(cbx_1__2__1_chanx_out_191_[0]),
		.chanx_right_in_193_(cbx_1__2__1_chanx_out_193_[0]),
		.chanx_right_in_195_(cbx_1__2__1_chanx_out_195_[0]),
		.chanx_right_in_197_(cbx_1__2__1_chanx_out_197_[0]),
		.chanx_right_in_199_(cbx_1__2__1_chanx_out_199_[0]),
		.right_top_grid_pin_1_(grid_io_top_1_bottom_width_0_height_0__pin_1_upper[0]),
		.chany_bottom_in_0_(cby_1__1__1_chany_out_0_[0]),
		.chany_bottom_in_2_(cby_1__1__1_chany_out_2_[0]),
		.chany_bottom_in_4_(cby_1__1__1_chany_out_4_[0]),
		.chany_bottom_in_6_(cby_1__1__1_chany_out_6_[0]),
		.chany_bottom_in_8_(cby_1__1__1_chany_out_8_[0]),
		.chany_bottom_in_10_(cby_1__1__1_chany_out_10_[0]),
		.chany_bottom_in_12_(cby_1__1__1_chany_out_12_[0]),
		.chany_bottom_in_14_(cby_1__1__1_chany_out_14_[0]),
		.chany_bottom_in_16_(cby_1__1__1_chany_out_16_[0]),
		.chany_bottom_in_18_(cby_1__1__1_chany_out_18_[0]),
		.chany_bottom_in_20_(cby_1__1__1_chany_out_20_[0]),
		.chany_bottom_in_22_(cby_1__1__1_chany_out_22_[0]),
		.chany_bottom_in_24_(cby_1__1__1_chany_out_24_[0]),
		.chany_bottom_in_26_(cby_1__1__1_chany_out_26_[0]),
		.chany_bottom_in_28_(cby_1__1__1_chany_out_28_[0]),
		.chany_bottom_in_30_(cby_1__1__1_chany_out_30_[0]),
		.chany_bottom_in_32_(cby_1__1__1_chany_out_32_[0]),
		.chany_bottom_in_34_(cby_1__1__1_chany_out_34_[0]),
		.chany_bottom_in_36_(cby_1__1__1_chany_out_36_[0]),
		.chany_bottom_in_38_(cby_1__1__1_chany_out_38_[0]),
		.chany_bottom_in_40_(cby_1__1__1_chany_out_40_[0]),
		.chany_bottom_in_42_(cby_1__1__1_chany_out_42_[0]),
		.chany_bottom_in_44_(cby_1__1__1_chany_out_44_[0]),
		.chany_bottom_in_46_(cby_1__1__1_chany_out_46_[0]),
		.chany_bottom_in_48_(cby_1__1__1_chany_out_48_[0]),
		.chany_bottom_in_50_(cby_1__1__1_chany_out_50_[0]),
		.chany_bottom_in_52_(cby_1__1__1_chany_out_52_[0]),
		.chany_bottom_in_54_(cby_1__1__1_chany_out_54_[0]),
		.chany_bottom_in_56_(cby_1__1__1_chany_out_56_[0]),
		.chany_bottom_in_58_(cby_1__1__1_chany_out_58_[0]),
		.chany_bottom_in_60_(cby_1__1__1_chany_out_60_[0]),
		.chany_bottom_in_62_(cby_1__1__1_chany_out_62_[0]),
		.chany_bottom_in_64_(cby_1__1__1_chany_out_64_[0]),
		.chany_bottom_in_66_(cby_1__1__1_chany_out_66_[0]),
		.chany_bottom_in_68_(cby_1__1__1_chany_out_68_[0]),
		.chany_bottom_in_70_(cby_1__1__1_chany_out_70_[0]),
		.chany_bottom_in_72_(cby_1__1__1_chany_out_72_[0]),
		.chany_bottom_in_74_(cby_1__1__1_chany_out_74_[0]),
		.chany_bottom_in_76_(cby_1__1__1_chany_out_76_[0]),
		.chany_bottom_in_78_(cby_1__1__1_chany_out_78_[0]),
		.chany_bottom_in_80_(cby_1__1__1_chany_out_80_[0]),
		.chany_bottom_in_82_(cby_1__1__1_chany_out_82_[0]),
		.chany_bottom_in_84_(cby_1__1__1_chany_out_84_[0]),
		.chany_bottom_in_86_(cby_1__1__1_chany_out_86_[0]),
		.chany_bottom_in_88_(cby_1__1__1_chany_out_88_[0]),
		.chany_bottom_in_90_(cby_1__1__1_chany_out_90_[0]),
		.chany_bottom_in_92_(cby_1__1__1_chany_out_92_[0]),
		.chany_bottom_in_94_(cby_1__1__1_chany_out_94_[0]),
		.chany_bottom_in_96_(cby_1__1__1_chany_out_96_[0]),
		.chany_bottom_in_98_(cby_1__1__1_chany_out_98_[0]),
		.chany_bottom_in_100_(cby_1__1__1_chany_out_100_[0]),
		.chany_bottom_in_102_(cby_1__1__1_chany_out_102_[0]),
		.chany_bottom_in_104_(cby_1__1__1_chany_out_104_[0]),
		.chany_bottom_in_106_(cby_1__1__1_chany_out_106_[0]),
		.chany_bottom_in_108_(cby_1__1__1_chany_out_108_[0]),
		.chany_bottom_in_110_(cby_1__1__1_chany_out_110_[0]),
		.chany_bottom_in_112_(cby_1__1__1_chany_out_112_[0]),
		.chany_bottom_in_114_(cby_1__1__1_chany_out_114_[0]),
		.chany_bottom_in_116_(cby_1__1__1_chany_out_116_[0]),
		.chany_bottom_in_118_(cby_1__1__1_chany_out_118_[0]),
		.chany_bottom_in_120_(cby_1__1__1_chany_out_120_[0]),
		.chany_bottom_in_122_(cby_1__1__1_chany_out_122_[0]),
		.chany_bottom_in_124_(cby_1__1__1_chany_out_124_[0]),
		.chany_bottom_in_126_(cby_1__1__1_chany_out_126_[0]),
		.chany_bottom_in_128_(cby_1__1__1_chany_out_128_[0]),
		.chany_bottom_in_130_(cby_1__1__1_chany_out_130_[0]),
		.chany_bottom_in_132_(cby_1__1__1_chany_out_132_[0]),
		.chany_bottom_in_134_(cby_1__1__1_chany_out_134_[0]),
		.chany_bottom_in_136_(cby_1__1__1_chany_out_136_[0]),
		.chany_bottom_in_138_(cby_1__1__1_chany_out_138_[0]),
		.chany_bottom_in_140_(cby_1__1__1_chany_out_140_[0]),
		.chany_bottom_in_142_(cby_1__1__1_chany_out_142_[0]),
		.chany_bottom_in_144_(cby_1__1__1_chany_out_144_[0]),
		.chany_bottom_in_146_(cby_1__1__1_chany_out_146_[0]),
		.chany_bottom_in_148_(cby_1__1__1_chany_out_148_[0]),
		.chany_bottom_in_150_(cby_1__1__1_chany_out_150_[0]),
		.chany_bottom_in_152_(cby_1__1__1_chany_out_152_[0]),
		.chany_bottom_in_154_(cby_1__1__1_chany_out_154_[0]),
		.chany_bottom_in_156_(cby_1__1__1_chany_out_156_[0]),
		.chany_bottom_in_158_(cby_1__1__1_chany_out_158_[0]),
		.chany_bottom_in_160_(cby_1__1__1_chany_out_160_[0]),
		.chany_bottom_in_162_(cby_1__1__1_chany_out_162_[0]),
		.chany_bottom_in_164_(cby_1__1__1_chany_out_164_[0]),
		.chany_bottom_in_166_(cby_1__1__1_chany_out_166_[0]),
		.chany_bottom_in_168_(cby_1__1__1_chany_out_168_[0]),
		.chany_bottom_in_170_(cby_1__1__1_chany_out_170_[0]),
		.chany_bottom_in_172_(cby_1__1__1_chany_out_172_[0]),
		.chany_bottom_in_174_(cby_1__1__1_chany_out_174_[0]),
		.chany_bottom_in_176_(cby_1__1__1_chany_out_176_[0]),
		.chany_bottom_in_178_(cby_1__1__1_chany_out_178_[0]),
		.chany_bottom_in_180_(cby_1__1__1_chany_out_180_[0]),
		.chany_bottom_in_182_(cby_1__1__1_chany_out_182_[0]),
		.chany_bottom_in_184_(cby_1__1__1_chany_out_184_[0]),
		.chany_bottom_in_186_(cby_1__1__1_chany_out_186_[0]),
		.chany_bottom_in_188_(cby_1__1__1_chany_out_188_[0]),
		.chany_bottom_in_190_(cby_1__1__1_chany_out_190_[0]),
		.chany_bottom_in_192_(cby_1__1__1_chany_out_192_[0]),
		.chany_bottom_in_194_(cby_1__1__1_chany_out_194_[0]),
		.chany_bottom_in_196_(cby_1__1__1_chany_out_196_[0]),
		.chany_bottom_in_198_(cby_1__1__1_chany_out_198_[0]),
		.bottom_left_grid_pin_44_(grid_clb_0_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_0_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_0_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_0_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_0_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_0_right_width_0_height_0__pin_49_upper[0]),
		.bottom_left_grid_pin_50_(grid_clb_0_right_width_0_height_0__pin_50_upper[0]),
		.bottom_left_grid_pin_51_(grid_clb_0_right_width_0_height_0__pin_51_upper[0]),
		.bottom_left_grid_pin_52_(grid_clb_0_right_width_0_height_0__pin_52_upper[0]),
		.bottom_left_grid_pin_53_(grid_clb_0_right_width_0_height_0__pin_53_upper[0]),
		.chanx_left_in_0_(cbx_1__2__0_chanx_out_0_[0]),
		.chanx_left_in_2_(cbx_1__2__0_chanx_out_2_[0]),
		.chanx_left_in_4_(cbx_1__2__0_chanx_out_4_[0]),
		.chanx_left_in_6_(cbx_1__2__0_chanx_out_6_[0]),
		.chanx_left_in_8_(cbx_1__2__0_chanx_out_8_[0]),
		.chanx_left_in_10_(cbx_1__2__0_chanx_out_10_[0]),
		.chanx_left_in_12_(cbx_1__2__0_chanx_out_12_[0]),
		.chanx_left_in_14_(cbx_1__2__0_chanx_out_14_[0]),
		.chanx_left_in_16_(cbx_1__2__0_chanx_out_16_[0]),
		.chanx_left_in_18_(cbx_1__2__0_chanx_out_18_[0]),
		.chanx_left_in_20_(cbx_1__2__0_chanx_out_20_[0]),
		.chanx_left_in_22_(cbx_1__2__0_chanx_out_22_[0]),
		.chanx_left_in_24_(cbx_1__2__0_chanx_out_24_[0]),
		.chanx_left_in_26_(cbx_1__2__0_chanx_out_26_[0]),
		.chanx_left_in_28_(cbx_1__2__0_chanx_out_28_[0]),
		.chanx_left_in_30_(cbx_1__2__0_chanx_out_30_[0]),
		.chanx_left_in_32_(cbx_1__2__0_chanx_out_32_[0]),
		.chanx_left_in_34_(cbx_1__2__0_chanx_out_34_[0]),
		.chanx_left_in_36_(cbx_1__2__0_chanx_out_36_[0]),
		.chanx_left_in_38_(cbx_1__2__0_chanx_out_38_[0]),
		.chanx_left_in_40_(cbx_1__2__0_chanx_out_40_[0]),
		.chanx_left_in_42_(cbx_1__2__0_chanx_out_42_[0]),
		.chanx_left_in_44_(cbx_1__2__0_chanx_out_44_[0]),
		.chanx_left_in_46_(cbx_1__2__0_chanx_out_46_[0]),
		.chanx_left_in_48_(cbx_1__2__0_chanx_out_48_[0]),
		.chanx_left_in_50_(cbx_1__2__0_chanx_out_50_[0]),
		.chanx_left_in_52_(cbx_1__2__0_chanx_out_52_[0]),
		.chanx_left_in_54_(cbx_1__2__0_chanx_out_54_[0]),
		.chanx_left_in_56_(cbx_1__2__0_chanx_out_56_[0]),
		.chanx_left_in_58_(cbx_1__2__0_chanx_out_58_[0]),
		.chanx_left_in_60_(cbx_1__2__0_chanx_out_60_[0]),
		.chanx_left_in_62_(cbx_1__2__0_chanx_out_62_[0]),
		.chanx_left_in_64_(cbx_1__2__0_chanx_out_64_[0]),
		.chanx_left_in_66_(cbx_1__2__0_chanx_out_66_[0]),
		.chanx_left_in_68_(cbx_1__2__0_chanx_out_68_[0]),
		.chanx_left_in_70_(cbx_1__2__0_chanx_out_70_[0]),
		.chanx_left_in_72_(cbx_1__2__0_chanx_out_72_[0]),
		.chanx_left_in_74_(cbx_1__2__0_chanx_out_74_[0]),
		.chanx_left_in_76_(cbx_1__2__0_chanx_out_76_[0]),
		.chanx_left_in_78_(cbx_1__2__0_chanx_out_78_[0]),
		.chanx_left_in_80_(cbx_1__2__0_chanx_out_80_[0]),
		.chanx_left_in_82_(cbx_1__2__0_chanx_out_82_[0]),
		.chanx_left_in_84_(cbx_1__2__0_chanx_out_84_[0]),
		.chanx_left_in_86_(cbx_1__2__0_chanx_out_86_[0]),
		.chanx_left_in_88_(cbx_1__2__0_chanx_out_88_[0]),
		.chanx_left_in_90_(cbx_1__2__0_chanx_out_90_[0]),
		.chanx_left_in_92_(cbx_1__2__0_chanx_out_92_[0]),
		.chanx_left_in_94_(cbx_1__2__0_chanx_out_94_[0]),
		.chanx_left_in_96_(cbx_1__2__0_chanx_out_96_[0]),
		.chanx_left_in_98_(cbx_1__2__0_chanx_out_98_[0]),
		.chanx_left_in_100_(cbx_1__2__0_chanx_out_100_[0]),
		.chanx_left_in_102_(cbx_1__2__0_chanx_out_102_[0]),
		.chanx_left_in_104_(cbx_1__2__0_chanx_out_104_[0]),
		.chanx_left_in_106_(cbx_1__2__0_chanx_out_106_[0]),
		.chanx_left_in_108_(cbx_1__2__0_chanx_out_108_[0]),
		.chanx_left_in_110_(cbx_1__2__0_chanx_out_110_[0]),
		.chanx_left_in_112_(cbx_1__2__0_chanx_out_112_[0]),
		.chanx_left_in_114_(cbx_1__2__0_chanx_out_114_[0]),
		.chanx_left_in_116_(cbx_1__2__0_chanx_out_116_[0]),
		.chanx_left_in_118_(cbx_1__2__0_chanx_out_118_[0]),
		.chanx_left_in_120_(cbx_1__2__0_chanx_out_120_[0]),
		.chanx_left_in_122_(cbx_1__2__0_chanx_out_122_[0]),
		.chanx_left_in_124_(cbx_1__2__0_chanx_out_124_[0]),
		.chanx_left_in_126_(cbx_1__2__0_chanx_out_126_[0]),
		.chanx_left_in_128_(cbx_1__2__0_chanx_out_128_[0]),
		.chanx_left_in_130_(cbx_1__2__0_chanx_out_130_[0]),
		.chanx_left_in_132_(cbx_1__2__0_chanx_out_132_[0]),
		.chanx_left_in_134_(cbx_1__2__0_chanx_out_134_[0]),
		.chanx_left_in_136_(cbx_1__2__0_chanx_out_136_[0]),
		.chanx_left_in_138_(cbx_1__2__0_chanx_out_138_[0]),
		.chanx_left_in_140_(cbx_1__2__0_chanx_out_140_[0]),
		.chanx_left_in_142_(cbx_1__2__0_chanx_out_142_[0]),
		.chanx_left_in_144_(cbx_1__2__0_chanx_out_144_[0]),
		.chanx_left_in_146_(cbx_1__2__0_chanx_out_146_[0]),
		.chanx_left_in_148_(cbx_1__2__0_chanx_out_148_[0]),
		.chanx_left_in_150_(cbx_1__2__0_chanx_out_150_[0]),
		.chanx_left_in_152_(cbx_1__2__0_chanx_out_152_[0]),
		.chanx_left_in_154_(cbx_1__2__0_chanx_out_154_[0]),
		.chanx_left_in_156_(cbx_1__2__0_chanx_out_156_[0]),
		.chanx_left_in_158_(cbx_1__2__0_chanx_out_158_[0]),
		.chanx_left_in_160_(cbx_1__2__0_chanx_out_160_[0]),
		.chanx_left_in_162_(cbx_1__2__0_chanx_out_162_[0]),
		.chanx_left_in_164_(cbx_1__2__0_chanx_out_164_[0]),
		.chanx_left_in_166_(cbx_1__2__0_chanx_out_166_[0]),
		.chanx_left_in_168_(cbx_1__2__0_chanx_out_168_[0]),
		.chanx_left_in_170_(cbx_1__2__0_chanx_out_170_[0]),
		.chanx_left_in_172_(cbx_1__2__0_chanx_out_172_[0]),
		.chanx_left_in_174_(cbx_1__2__0_chanx_out_174_[0]),
		.chanx_left_in_176_(cbx_1__2__0_chanx_out_176_[0]),
		.chanx_left_in_178_(cbx_1__2__0_chanx_out_178_[0]),
		.chanx_left_in_180_(cbx_1__2__0_chanx_out_180_[0]),
		.chanx_left_in_182_(cbx_1__2__0_chanx_out_182_[0]),
		.chanx_left_in_184_(cbx_1__2__0_chanx_out_184_[0]),
		.chanx_left_in_186_(cbx_1__2__0_chanx_out_186_[0]),
		.chanx_left_in_188_(cbx_1__2__0_chanx_out_188_[0]),
		.chanx_left_in_190_(cbx_1__2__0_chanx_out_190_[0]),
		.chanx_left_in_192_(cbx_1__2__0_chanx_out_192_[0]),
		.chanx_left_in_194_(cbx_1__2__0_chanx_out_194_[0]),
		.chanx_left_in_196_(cbx_1__2__0_chanx_out_196_[0]),
		.chanx_left_in_198_(cbx_1__2__0_chanx_out_198_[0]),
		.left_top_grid_pin_1_(grid_io_top_0_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_io_top_1_ccff_tail[0]),
		.chanx_right_out_0_(sb_1__2__0_chanx_right_out_0_[0]),
		.chanx_right_out_2_(sb_1__2__0_chanx_right_out_2_[0]),
		.chanx_right_out_4_(sb_1__2__0_chanx_right_out_4_[0]),
		.chanx_right_out_6_(sb_1__2__0_chanx_right_out_6_[0]),
		.chanx_right_out_8_(sb_1__2__0_chanx_right_out_8_[0]),
		.chanx_right_out_10_(sb_1__2__0_chanx_right_out_10_[0]),
		.chanx_right_out_12_(sb_1__2__0_chanx_right_out_12_[0]),
		.chanx_right_out_14_(sb_1__2__0_chanx_right_out_14_[0]),
		.chanx_right_out_16_(sb_1__2__0_chanx_right_out_16_[0]),
		.chanx_right_out_18_(sb_1__2__0_chanx_right_out_18_[0]),
		.chanx_right_out_20_(sb_1__2__0_chanx_right_out_20_[0]),
		.chanx_right_out_22_(sb_1__2__0_chanx_right_out_22_[0]),
		.chanx_right_out_24_(sb_1__2__0_chanx_right_out_24_[0]),
		.chanx_right_out_26_(sb_1__2__0_chanx_right_out_26_[0]),
		.chanx_right_out_28_(sb_1__2__0_chanx_right_out_28_[0]),
		.chanx_right_out_30_(sb_1__2__0_chanx_right_out_30_[0]),
		.chanx_right_out_32_(sb_1__2__0_chanx_right_out_32_[0]),
		.chanx_right_out_34_(sb_1__2__0_chanx_right_out_34_[0]),
		.chanx_right_out_36_(sb_1__2__0_chanx_right_out_36_[0]),
		.chanx_right_out_38_(sb_1__2__0_chanx_right_out_38_[0]),
		.chanx_right_out_40_(sb_1__2__0_chanx_right_out_40_[0]),
		.chanx_right_out_42_(sb_1__2__0_chanx_right_out_42_[0]),
		.chanx_right_out_44_(sb_1__2__0_chanx_right_out_44_[0]),
		.chanx_right_out_46_(sb_1__2__0_chanx_right_out_46_[0]),
		.chanx_right_out_48_(sb_1__2__0_chanx_right_out_48_[0]),
		.chanx_right_out_50_(sb_1__2__0_chanx_right_out_50_[0]),
		.chanx_right_out_52_(sb_1__2__0_chanx_right_out_52_[0]),
		.chanx_right_out_54_(sb_1__2__0_chanx_right_out_54_[0]),
		.chanx_right_out_56_(sb_1__2__0_chanx_right_out_56_[0]),
		.chanx_right_out_58_(sb_1__2__0_chanx_right_out_58_[0]),
		.chanx_right_out_60_(sb_1__2__0_chanx_right_out_60_[0]),
		.chanx_right_out_62_(sb_1__2__0_chanx_right_out_62_[0]),
		.chanx_right_out_64_(sb_1__2__0_chanx_right_out_64_[0]),
		.chanx_right_out_66_(sb_1__2__0_chanx_right_out_66_[0]),
		.chanx_right_out_68_(sb_1__2__0_chanx_right_out_68_[0]),
		.chanx_right_out_70_(sb_1__2__0_chanx_right_out_70_[0]),
		.chanx_right_out_72_(sb_1__2__0_chanx_right_out_72_[0]),
		.chanx_right_out_74_(sb_1__2__0_chanx_right_out_74_[0]),
		.chanx_right_out_76_(sb_1__2__0_chanx_right_out_76_[0]),
		.chanx_right_out_78_(sb_1__2__0_chanx_right_out_78_[0]),
		.chanx_right_out_80_(sb_1__2__0_chanx_right_out_80_[0]),
		.chanx_right_out_82_(sb_1__2__0_chanx_right_out_82_[0]),
		.chanx_right_out_84_(sb_1__2__0_chanx_right_out_84_[0]),
		.chanx_right_out_86_(sb_1__2__0_chanx_right_out_86_[0]),
		.chanx_right_out_88_(sb_1__2__0_chanx_right_out_88_[0]),
		.chanx_right_out_90_(sb_1__2__0_chanx_right_out_90_[0]),
		.chanx_right_out_92_(sb_1__2__0_chanx_right_out_92_[0]),
		.chanx_right_out_94_(sb_1__2__0_chanx_right_out_94_[0]),
		.chanx_right_out_96_(sb_1__2__0_chanx_right_out_96_[0]),
		.chanx_right_out_98_(sb_1__2__0_chanx_right_out_98_[0]),
		.chanx_right_out_100_(sb_1__2__0_chanx_right_out_100_[0]),
		.chanx_right_out_102_(sb_1__2__0_chanx_right_out_102_[0]),
		.chanx_right_out_104_(sb_1__2__0_chanx_right_out_104_[0]),
		.chanx_right_out_106_(sb_1__2__0_chanx_right_out_106_[0]),
		.chanx_right_out_108_(sb_1__2__0_chanx_right_out_108_[0]),
		.chanx_right_out_110_(sb_1__2__0_chanx_right_out_110_[0]),
		.chanx_right_out_112_(sb_1__2__0_chanx_right_out_112_[0]),
		.chanx_right_out_114_(sb_1__2__0_chanx_right_out_114_[0]),
		.chanx_right_out_116_(sb_1__2__0_chanx_right_out_116_[0]),
		.chanx_right_out_118_(sb_1__2__0_chanx_right_out_118_[0]),
		.chanx_right_out_120_(sb_1__2__0_chanx_right_out_120_[0]),
		.chanx_right_out_122_(sb_1__2__0_chanx_right_out_122_[0]),
		.chanx_right_out_124_(sb_1__2__0_chanx_right_out_124_[0]),
		.chanx_right_out_126_(sb_1__2__0_chanx_right_out_126_[0]),
		.chanx_right_out_128_(sb_1__2__0_chanx_right_out_128_[0]),
		.chanx_right_out_130_(sb_1__2__0_chanx_right_out_130_[0]),
		.chanx_right_out_132_(sb_1__2__0_chanx_right_out_132_[0]),
		.chanx_right_out_134_(sb_1__2__0_chanx_right_out_134_[0]),
		.chanx_right_out_136_(sb_1__2__0_chanx_right_out_136_[0]),
		.chanx_right_out_138_(sb_1__2__0_chanx_right_out_138_[0]),
		.chanx_right_out_140_(sb_1__2__0_chanx_right_out_140_[0]),
		.chanx_right_out_142_(sb_1__2__0_chanx_right_out_142_[0]),
		.chanx_right_out_144_(sb_1__2__0_chanx_right_out_144_[0]),
		.chanx_right_out_146_(sb_1__2__0_chanx_right_out_146_[0]),
		.chanx_right_out_148_(sb_1__2__0_chanx_right_out_148_[0]),
		.chanx_right_out_150_(sb_1__2__0_chanx_right_out_150_[0]),
		.chanx_right_out_152_(sb_1__2__0_chanx_right_out_152_[0]),
		.chanx_right_out_154_(sb_1__2__0_chanx_right_out_154_[0]),
		.chanx_right_out_156_(sb_1__2__0_chanx_right_out_156_[0]),
		.chanx_right_out_158_(sb_1__2__0_chanx_right_out_158_[0]),
		.chanx_right_out_160_(sb_1__2__0_chanx_right_out_160_[0]),
		.chanx_right_out_162_(sb_1__2__0_chanx_right_out_162_[0]),
		.chanx_right_out_164_(sb_1__2__0_chanx_right_out_164_[0]),
		.chanx_right_out_166_(sb_1__2__0_chanx_right_out_166_[0]),
		.chanx_right_out_168_(sb_1__2__0_chanx_right_out_168_[0]),
		.chanx_right_out_170_(sb_1__2__0_chanx_right_out_170_[0]),
		.chanx_right_out_172_(sb_1__2__0_chanx_right_out_172_[0]),
		.chanx_right_out_174_(sb_1__2__0_chanx_right_out_174_[0]),
		.chanx_right_out_176_(sb_1__2__0_chanx_right_out_176_[0]),
		.chanx_right_out_178_(sb_1__2__0_chanx_right_out_178_[0]),
		.chanx_right_out_180_(sb_1__2__0_chanx_right_out_180_[0]),
		.chanx_right_out_182_(sb_1__2__0_chanx_right_out_182_[0]),
		.chanx_right_out_184_(sb_1__2__0_chanx_right_out_184_[0]),
		.chanx_right_out_186_(sb_1__2__0_chanx_right_out_186_[0]),
		.chanx_right_out_188_(sb_1__2__0_chanx_right_out_188_[0]),
		.chanx_right_out_190_(sb_1__2__0_chanx_right_out_190_[0]),
		.chanx_right_out_192_(sb_1__2__0_chanx_right_out_192_[0]),
		.chanx_right_out_194_(sb_1__2__0_chanx_right_out_194_[0]),
		.chanx_right_out_196_(sb_1__2__0_chanx_right_out_196_[0]),
		.chanx_right_out_198_(sb_1__2__0_chanx_right_out_198_[0]),
		.chany_bottom_out_1_(sb_1__2__0_chany_bottom_out_1_[0]),
		.chany_bottom_out_3_(sb_1__2__0_chany_bottom_out_3_[0]),
		.chany_bottom_out_5_(sb_1__2__0_chany_bottom_out_5_[0]),
		.chany_bottom_out_7_(sb_1__2__0_chany_bottom_out_7_[0]),
		.chany_bottom_out_9_(sb_1__2__0_chany_bottom_out_9_[0]),
		.chany_bottom_out_11_(sb_1__2__0_chany_bottom_out_11_[0]),
		.chany_bottom_out_13_(sb_1__2__0_chany_bottom_out_13_[0]),
		.chany_bottom_out_15_(sb_1__2__0_chany_bottom_out_15_[0]),
		.chany_bottom_out_17_(sb_1__2__0_chany_bottom_out_17_[0]),
		.chany_bottom_out_19_(sb_1__2__0_chany_bottom_out_19_[0]),
		.chany_bottom_out_21_(sb_1__2__0_chany_bottom_out_21_[0]),
		.chany_bottom_out_23_(sb_1__2__0_chany_bottom_out_23_[0]),
		.chany_bottom_out_25_(sb_1__2__0_chany_bottom_out_25_[0]),
		.chany_bottom_out_27_(sb_1__2__0_chany_bottom_out_27_[0]),
		.chany_bottom_out_29_(sb_1__2__0_chany_bottom_out_29_[0]),
		.chany_bottom_out_31_(sb_1__2__0_chany_bottom_out_31_[0]),
		.chany_bottom_out_33_(sb_1__2__0_chany_bottom_out_33_[0]),
		.chany_bottom_out_35_(sb_1__2__0_chany_bottom_out_35_[0]),
		.chany_bottom_out_37_(sb_1__2__0_chany_bottom_out_37_[0]),
		.chany_bottom_out_39_(sb_1__2__0_chany_bottom_out_39_[0]),
		.chany_bottom_out_41_(sb_1__2__0_chany_bottom_out_41_[0]),
		.chany_bottom_out_43_(sb_1__2__0_chany_bottom_out_43_[0]),
		.chany_bottom_out_45_(sb_1__2__0_chany_bottom_out_45_[0]),
		.chany_bottom_out_47_(sb_1__2__0_chany_bottom_out_47_[0]),
		.chany_bottom_out_49_(sb_1__2__0_chany_bottom_out_49_[0]),
		.chany_bottom_out_51_(sb_1__2__0_chany_bottom_out_51_[0]),
		.chany_bottom_out_53_(sb_1__2__0_chany_bottom_out_53_[0]),
		.chany_bottom_out_55_(sb_1__2__0_chany_bottom_out_55_[0]),
		.chany_bottom_out_57_(sb_1__2__0_chany_bottom_out_57_[0]),
		.chany_bottom_out_59_(sb_1__2__0_chany_bottom_out_59_[0]),
		.chany_bottom_out_61_(sb_1__2__0_chany_bottom_out_61_[0]),
		.chany_bottom_out_63_(sb_1__2__0_chany_bottom_out_63_[0]),
		.chany_bottom_out_65_(sb_1__2__0_chany_bottom_out_65_[0]),
		.chany_bottom_out_67_(sb_1__2__0_chany_bottom_out_67_[0]),
		.chany_bottom_out_69_(sb_1__2__0_chany_bottom_out_69_[0]),
		.chany_bottom_out_71_(sb_1__2__0_chany_bottom_out_71_[0]),
		.chany_bottom_out_73_(sb_1__2__0_chany_bottom_out_73_[0]),
		.chany_bottom_out_75_(sb_1__2__0_chany_bottom_out_75_[0]),
		.chany_bottom_out_77_(sb_1__2__0_chany_bottom_out_77_[0]),
		.chany_bottom_out_79_(sb_1__2__0_chany_bottom_out_79_[0]),
		.chany_bottom_out_81_(sb_1__2__0_chany_bottom_out_81_[0]),
		.chany_bottom_out_83_(sb_1__2__0_chany_bottom_out_83_[0]),
		.chany_bottom_out_85_(sb_1__2__0_chany_bottom_out_85_[0]),
		.chany_bottom_out_87_(sb_1__2__0_chany_bottom_out_87_[0]),
		.chany_bottom_out_89_(sb_1__2__0_chany_bottom_out_89_[0]),
		.chany_bottom_out_91_(sb_1__2__0_chany_bottom_out_91_[0]),
		.chany_bottom_out_93_(sb_1__2__0_chany_bottom_out_93_[0]),
		.chany_bottom_out_95_(sb_1__2__0_chany_bottom_out_95_[0]),
		.chany_bottom_out_97_(sb_1__2__0_chany_bottom_out_97_[0]),
		.chany_bottom_out_99_(sb_1__2__0_chany_bottom_out_99_[0]),
		.chany_bottom_out_101_(sb_1__2__0_chany_bottom_out_101_[0]),
		.chany_bottom_out_103_(sb_1__2__0_chany_bottom_out_103_[0]),
		.chany_bottom_out_105_(sb_1__2__0_chany_bottom_out_105_[0]),
		.chany_bottom_out_107_(sb_1__2__0_chany_bottom_out_107_[0]),
		.chany_bottom_out_109_(sb_1__2__0_chany_bottom_out_109_[0]),
		.chany_bottom_out_111_(sb_1__2__0_chany_bottom_out_111_[0]),
		.chany_bottom_out_113_(sb_1__2__0_chany_bottom_out_113_[0]),
		.chany_bottom_out_115_(sb_1__2__0_chany_bottom_out_115_[0]),
		.chany_bottom_out_117_(sb_1__2__0_chany_bottom_out_117_[0]),
		.chany_bottom_out_119_(sb_1__2__0_chany_bottom_out_119_[0]),
		.chany_bottom_out_121_(sb_1__2__0_chany_bottom_out_121_[0]),
		.chany_bottom_out_123_(sb_1__2__0_chany_bottom_out_123_[0]),
		.chany_bottom_out_125_(sb_1__2__0_chany_bottom_out_125_[0]),
		.chany_bottom_out_127_(sb_1__2__0_chany_bottom_out_127_[0]),
		.chany_bottom_out_129_(sb_1__2__0_chany_bottom_out_129_[0]),
		.chany_bottom_out_131_(sb_1__2__0_chany_bottom_out_131_[0]),
		.chany_bottom_out_133_(sb_1__2__0_chany_bottom_out_133_[0]),
		.chany_bottom_out_135_(sb_1__2__0_chany_bottom_out_135_[0]),
		.chany_bottom_out_137_(sb_1__2__0_chany_bottom_out_137_[0]),
		.chany_bottom_out_139_(sb_1__2__0_chany_bottom_out_139_[0]),
		.chany_bottom_out_141_(sb_1__2__0_chany_bottom_out_141_[0]),
		.chany_bottom_out_143_(sb_1__2__0_chany_bottom_out_143_[0]),
		.chany_bottom_out_145_(sb_1__2__0_chany_bottom_out_145_[0]),
		.chany_bottom_out_147_(sb_1__2__0_chany_bottom_out_147_[0]),
		.chany_bottom_out_149_(sb_1__2__0_chany_bottom_out_149_[0]),
		.chany_bottom_out_151_(sb_1__2__0_chany_bottom_out_151_[0]),
		.chany_bottom_out_153_(sb_1__2__0_chany_bottom_out_153_[0]),
		.chany_bottom_out_155_(sb_1__2__0_chany_bottom_out_155_[0]),
		.chany_bottom_out_157_(sb_1__2__0_chany_bottom_out_157_[0]),
		.chany_bottom_out_159_(sb_1__2__0_chany_bottom_out_159_[0]),
		.chany_bottom_out_161_(sb_1__2__0_chany_bottom_out_161_[0]),
		.chany_bottom_out_163_(sb_1__2__0_chany_bottom_out_163_[0]),
		.chany_bottom_out_165_(sb_1__2__0_chany_bottom_out_165_[0]),
		.chany_bottom_out_167_(sb_1__2__0_chany_bottom_out_167_[0]),
		.chany_bottom_out_169_(sb_1__2__0_chany_bottom_out_169_[0]),
		.chany_bottom_out_171_(sb_1__2__0_chany_bottom_out_171_[0]),
		.chany_bottom_out_173_(sb_1__2__0_chany_bottom_out_173_[0]),
		.chany_bottom_out_175_(sb_1__2__0_chany_bottom_out_175_[0]),
		.chany_bottom_out_177_(sb_1__2__0_chany_bottom_out_177_[0]),
		.chany_bottom_out_179_(sb_1__2__0_chany_bottom_out_179_[0]),
		.chany_bottom_out_181_(sb_1__2__0_chany_bottom_out_181_[0]),
		.chany_bottom_out_183_(sb_1__2__0_chany_bottom_out_183_[0]),
		.chany_bottom_out_185_(sb_1__2__0_chany_bottom_out_185_[0]),
		.chany_bottom_out_187_(sb_1__2__0_chany_bottom_out_187_[0]),
		.chany_bottom_out_189_(sb_1__2__0_chany_bottom_out_189_[0]),
		.chany_bottom_out_191_(sb_1__2__0_chany_bottom_out_191_[0]),
		.chany_bottom_out_193_(sb_1__2__0_chany_bottom_out_193_[0]),
		.chany_bottom_out_195_(sb_1__2__0_chany_bottom_out_195_[0]),
		.chany_bottom_out_197_(sb_1__2__0_chany_bottom_out_197_[0]),
		.chany_bottom_out_199_(sb_1__2__0_chany_bottom_out_199_[0]),
		.chanx_left_out_1_(sb_1__2__0_chanx_left_out_1_[0]),
		.chanx_left_out_3_(sb_1__2__0_chanx_left_out_3_[0]),
		.chanx_left_out_5_(sb_1__2__0_chanx_left_out_5_[0]),
		.chanx_left_out_7_(sb_1__2__0_chanx_left_out_7_[0]),
		.chanx_left_out_9_(sb_1__2__0_chanx_left_out_9_[0]),
		.chanx_left_out_11_(sb_1__2__0_chanx_left_out_11_[0]),
		.chanx_left_out_13_(sb_1__2__0_chanx_left_out_13_[0]),
		.chanx_left_out_15_(sb_1__2__0_chanx_left_out_15_[0]),
		.chanx_left_out_17_(sb_1__2__0_chanx_left_out_17_[0]),
		.chanx_left_out_19_(sb_1__2__0_chanx_left_out_19_[0]),
		.chanx_left_out_21_(sb_1__2__0_chanx_left_out_21_[0]),
		.chanx_left_out_23_(sb_1__2__0_chanx_left_out_23_[0]),
		.chanx_left_out_25_(sb_1__2__0_chanx_left_out_25_[0]),
		.chanx_left_out_27_(sb_1__2__0_chanx_left_out_27_[0]),
		.chanx_left_out_29_(sb_1__2__0_chanx_left_out_29_[0]),
		.chanx_left_out_31_(sb_1__2__0_chanx_left_out_31_[0]),
		.chanx_left_out_33_(sb_1__2__0_chanx_left_out_33_[0]),
		.chanx_left_out_35_(sb_1__2__0_chanx_left_out_35_[0]),
		.chanx_left_out_37_(sb_1__2__0_chanx_left_out_37_[0]),
		.chanx_left_out_39_(sb_1__2__0_chanx_left_out_39_[0]),
		.chanx_left_out_41_(sb_1__2__0_chanx_left_out_41_[0]),
		.chanx_left_out_43_(sb_1__2__0_chanx_left_out_43_[0]),
		.chanx_left_out_45_(sb_1__2__0_chanx_left_out_45_[0]),
		.chanx_left_out_47_(sb_1__2__0_chanx_left_out_47_[0]),
		.chanx_left_out_49_(sb_1__2__0_chanx_left_out_49_[0]),
		.chanx_left_out_51_(sb_1__2__0_chanx_left_out_51_[0]),
		.chanx_left_out_53_(sb_1__2__0_chanx_left_out_53_[0]),
		.chanx_left_out_55_(sb_1__2__0_chanx_left_out_55_[0]),
		.chanx_left_out_57_(sb_1__2__0_chanx_left_out_57_[0]),
		.chanx_left_out_59_(sb_1__2__0_chanx_left_out_59_[0]),
		.chanx_left_out_61_(sb_1__2__0_chanx_left_out_61_[0]),
		.chanx_left_out_63_(sb_1__2__0_chanx_left_out_63_[0]),
		.chanx_left_out_65_(sb_1__2__0_chanx_left_out_65_[0]),
		.chanx_left_out_67_(sb_1__2__0_chanx_left_out_67_[0]),
		.chanx_left_out_69_(sb_1__2__0_chanx_left_out_69_[0]),
		.chanx_left_out_71_(sb_1__2__0_chanx_left_out_71_[0]),
		.chanx_left_out_73_(sb_1__2__0_chanx_left_out_73_[0]),
		.chanx_left_out_75_(sb_1__2__0_chanx_left_out_75_[0]),
		.chanx_left_out_77_(sb_1__2__0_chanx_left_out_77_[0]),
		.chanx_left_out_79_(sb_1__2__0_chanx_left_out_79_[0]),
		.chanx_left_out_81_(sb_1__2__0_chanx_left_out_81_[0]),
		.chanx_left_out_83_(sb_1__2__0_chanx_left_out_83_[0]),
		.chanx_left_out_85_(sb_1__2__0_chanx_left_out_85_[0]),
		.chanx_left_out_87_(sb_1__2__0_chanx_left_out_87_[0]),
		.chanx_left_out_89_(sb_1__2__0_chanx_left_out_89_[0]),
		.chanx_left_out_91_(sb_1__2__0_chanx_left_out_91_[0]),
		.chanx_left_out_93_(sb_1__2__0_chanx_left_out_93_[0]),
		.chanx_left_out_95_(sb_1__2__0_chanx_left_out_95_[0]),
		.chanx_left_out_97_(sb_1__2__0_chanx_left_out_97_[0]),
		.chanx_left_out_99_(sb_1__2__0_chanx_left_out_99_[0]),
		.chanx_left_out_101_(sb_1__2__0_chanx_left_out_101_[0]),
		.chanx_left_out_103_(sb_1__2__0_chanx_left_out_103_[0]),
		.chanx_left_out_105_(sb_1__2__0_chanx_left_out_105_[0]),
		.chanx_left_out_107_(sb_1__2__0_chanx_left_out_107_[0]),
		.chanx_left_out_109_(sb_1__2__0_chanx_left_out_109_[0]),
		.chanx_left_out_111_(sb_1__2__0_chanx_left_out_111_[0]),
		.chanx_left_out_113_(sb_1__2__0_chanx_left_out_113_[0]),
		.chanx_left_out_115_(sb_1__2__0_chanx_left_out_115_[0]),
		.chanx_left_out_117_(sb_1__2__0_chanx_left_out_117_[0]),
		.chanx_left_out_119_(sb_1__2__0_chanx_left_out_119_[0]),
		.chanx_left_out_121_(sb_1__2__0_chanx_left_out_121_[0]),
		.chanx_left_out_123_(sb_1__2__0_chanx_left_out_123_[0]),
		.chanx_left_out_125_(sb_1__2__0_chanx_left_out_125_[0]),
		.chanx_left_out_127_(sb_1__2__0_chanx_left_out_127_[0]),
		.chanx_left_out_129_(sb_1__2__0_chanx_left_out_129_[0]),
		.chanx_left_out_131_(sb_1__2__0_chanx_left_out_131_[0]),
		.chanx_left_out_133_(sb_1__2__0_chanx_left_out_133_[0]),
		.chanx_left_out_135_(sb_1__2__0_chanx_left_out_135_[0]),
		.chanx_left_out_137_(sb_1__2__0_chanx_left_out_137_[0]),
		.chanx_left_out_139_(sb_1__2__0_chanx_left_out_139_[0]),
		.chanx_left_out_141_(sb_1__2__0_chanx_left_out_141_[0]),
		.chanx_left_out_143_(sb_1__2__0_chanx_left_out_143_[0]),
		.chanx_left_out_145_(sb_1__2__0_chanx_left_out_145_[0]),
		.chanx_left_out_147_(sb_1__2__0_chanx_left_out_147_[0]),
		.chanx_left_out_149_(sb_1__2__0_chanx_left_out_149_[0]),
		.chanx_left_out_151_(sb_1__2__0_chanx_left_out_151_[0]),
		.chanx_left_out_153_(sb_1__2__0_chanx_left_out_153_[0]),
		.chanx_left_out_155_(sb_1__2__0_chanx_left_out_155_[0]),
		.chanx_left_out_157_(sb_1__2__0_chanx_left_out_157_[0]),
		.chanx_left_out_159_(sb_1__2__0_chanx_left_out_159_[0]),
		.chanx_left_out_161_(sb_1__2__0_chanx_left_out_161_[0]),
		.chanx_left_out_163_(sb_1__2__0_chanx_left_out_163_[0]),
		.chanx_left_out_165_(sb_1__2__0_chanx_left_out_165_[0]),
		.chanx_left_out_167_(sb_1__2__0_chanx_left_out_167_[0]),
		.chanx_left_out_169_(sb_1__2__0_chanx_left_out_169_[0]),
		.chanx_left_out_171_(sb_1__2__0_chanx_left_out_171_[0]),
		.chanx_left_out_173_(sb_1__2__0_chanx_left_out_173_[0]),
		.chanx_left_out_175_(sb_1__2__0_chanx_left_out_175_[0]),
		.chanx_left_out_177_(sb_1__2__0_chanx_left_out_177_[0]),
		.chanx_left_out_179_(sb_1__2__0_chanx_left_out_179_[0]),
		.chanx_left_out_181_(sb_1__2__0_chanx_left_out_181_[0]),
		.chanx_left_out_183_(sb_1__2__0_chanx_left_out_183_[0]),
		.chanx_left_out_185_(sb_1__2__0_chanx_left_out_185_[0]),
		.chanx_left_out_187_(sb_1__2__0_chanx_left_out_187_[0]),
		.chanx_left_out_189_(sb_1__2__0_chanx_left_out_189_[0]),
		.chanx_left_out_191_(sb_1__2__0_chanx_left_out_191_[0]),
		.chanx_left_out_193_(sb_1__2__0_chanx_left_out_193_[0]),
		.chanx_left_out_195_(sb_1__2__0_chanx_left_out_195_[0]),
		.chanx_left_out_197_(sb_1__2__0_chanx_left_out_197_[0]),
		.chanx_left_out_199_(sb_1__2__0_chanx_left_out_199_[0]),
		.ccff_tail(sb_1__2__0_ccff_tail[0]));

	sb_2__0_ sb_2__0_ (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.chany_top_in_1_(cby_2__1__0_chany_out_1_[0]),
		.chany_top_in_3_(cby_2__1__0_chany_out_3_[0]),
		.chany_top_in_5_(cby_2__1__0_chany_out_5_[0]),
		.chany_top_in_7_(cby_2__1__0_chany_out_7_[0]),
		.chany_top_in_9_(cby_2__1__0_chany_out_9_[0]),
		.chany_top_in_11_(cby_2__1__0_chany_out_11_[0]),
		.chany_top_in_13_(cby_2__1__0_chany_out_13_[0]),
		.chany_top_in_15_(cby_2__1__0_chany_out_15_[0]),
		.chany_top_in_17_(cby_2__1__0_chany_out_17_[0]),
		.chany_top_in_19_(cby_2__1__0_chany_out_19_[0]),
		.chany_top_in_21_(cby_2__1__0_chany_out_21_[0]),
		.chany_top_in_23_(cby_2__1__0_chany_out_23_[0]),
		.chany_top_in_25_(cby_2__1__0_chany_out_25_[0]),
		.chany_top_in_27_(cby_2__1__0_chany_out_27_[0]),
		.chany_top_in_29_(cby_2__1__0_chany_out_29_[0]),
		.chany_top_in_31_(cby_2__1__0_chany_out_31_[0]),
		.chany_top_in_33_(cby_2__1__0_chany_out_33_[0]),
		.chany_top_in_35_(cby_2__1__0_chany_out_35_[0]),
		.chany_top_in_37_(cby_2__1__0_chany_out_37_[0]),
		.chany_top_in_39_(cby_2__1__0_chany_out_39_[0]),
		.chany_top_in_41_(cby_2__1__0_chany_out_41_[0]),
		.chany_top_in_43_(cby_2__1__0_chany_out_43_[0]),
		.chany_top_in_45_(cby_2__1__0_chany_out_45_[0]),
		.chany_top_in_47_(cby_2__1__0_chany_out_47_[0]),
		.chany_top_in_49_(cby_2__1__0_chany_out_49_[0]),
		.chany_top_in_51_(cby_2__1__0_chany_out_51_[0]),
		.chany_top_in_53_(cby_2__1__0_chany_out_53_[0]),
		.chany_top_in_55_(cby_2__1__0_chany_out_55_[0]),
		.chany_top_in_57_(cby_2__1__0_chany_out_57_[0]),
		.chany_top_in_59_(cby_2__1__0_chany_out_59_[0]),
		.chany_top_in_61_(cby_2__1__0_chany_out_61_[0]),
		.chany_top_in_63_(cby_2__1__0_chany_out_63_[0]),
		.chany_top_in_65_(cby_2__1__0_chany_out_65_[0]),
		.chany_top_in_67_(cby_2__1__0_chany_out_67_[0]),
		.chany_top_in_69_(cby_2__1__0_chany_out_69_[0]),
		.chany_top_in_71_(cby_2__1__0_chany_out_71_[0]),
		.chany_top_in_73_(cby_2__1__0_chany_out_73_[0]),
		.chany_top_in_75_(cby_2__1__0_chany_out_75_[0]),
		.chany_top_in_77_(cby_2__1__0_chany_out_77_[0]),
		.chany_top_in_79_(cby_2__1__0_chany_out_79_[0]),
		.chany_top_in_81_(cby_2__1__0_chany_out_81_[0]),
		.chany_top_in_83_(cby_2__1__0_chany_out_83_[0]),
		.chany_top_in_85_(cby_2__1__0_chany_out_85_[0]),
		.chany_top_in_87_(cby_2__1__0_chany_out_87_[0]),
		.chany_top_in_89_(cby_2__1__0_chany_out_89_[0]),
		.chany_top_in_91_(cby_2__1__0_chany_out_91_[0]),
		.chany_top_in_93_(cby_2__1__0_chany_out_93_[0]),
		.chany_top_in_95_(cby_2__1__0_chany_out_95_[0]),
		.chany_top_in_97_(cby_2__1__0_chany_out_97_[0]),
		.chany_top_in_99_(cby_2__1__0_chany_out_99_[0]),
		.chany_top_in_101_(cby_2__1__0_chany_out_101_[0]),
		.chany_top_in_103_(cby_2__1__0_chany_out_103_[0]),
		.chany_top_in_105_(cby_2__1__0_chany_out_105_[0]),
		.chany_top_in_107_(cby_2__1__0_chany_out_107_[0]),
		.chany_top_in_109_(cby_2__1__0_chany_out_109_[0]),
		.chany_top_in_111_(cby_2__1__0_chany_out_111_[0]),
		.chany_top_in_113_(cby_2__1__0_chany_out_113_[0]),
		.chany_top_in_115_(cby_2__1__0_chany_out_115_[0]),
		.chany_top_in_117_(cby_2__1__0_chany_out_117_[0]),
		.chany_top_in_119_(cby_2__1__0_chany_out_119_[0]),
		.chany_top_in_121_(cby_2__1__0_chany_out_121_[0]),
		.chany_top_in_123_(cby_2__1__0_chany_out_123_[0]),
		.chany_top_in_125_(cby_2__1__0_chany_out_125_[0]),
		.chany_top_in_127_(cby_2__1__0_chany_out_127_[0]),
		.chany_top_in_129_(cby_2__1__0_chany_out_129_[0]),
		.chany_top_in_131_(cby_2__1__0_chany_out_131_[0]),
		.chany_top_in_133_(cby_2__1__0_chany_out_133_[0]),
		.chany_top_in_135_(cby_2__1__0_chany_out_135_[0]),
		.chany_top_in_137_(cby_2__1__0_chany_out_137_[0]),
		.chany_top_in_139_(cby_2__1__0_chany_out_139_[0]),
		.chany_top_in_141_(cby_2__1__0_chany_out_141_[0]),
		.chany_top_in_143_(cby_2__1__0_chany_out_143_[0]),
		.chany_top_in_145_(cby_2__1__0_chany_out_145_[0]),
		.chany_top_in_147_(cby_2__1__0_chany_out_147_[0]),
		.chany_top_in_149_(cby_2__1__0_chany_out_149_[0]),
		.chany_top_in_151_(cby_2__1__0_chany_out_151_[0]),
		.chany_top_in_153_(cby_2__1__0_chany_out_153_[0]),
		.chany_top_in_155_(cby_2__1__0_chany_out_155_[0]),
		.chany_top_in_157_(cby_2__1__0_chany_out_157_[0]),
		.chany_top_in_159_(cby_2__1__0_chany_out_159_[0]),
		.chany_top_in_161_(cby_2__1__0_chany_out_161_[0]),
		.chany_top_in_163_(cby_2__1__0_chany_out_163_[0]),
		.chany_top_in_165_(cby_2__1__0_chany_out_165_[0]),
		.chany_top_in_167_(cby_2__1__0_chany_out_167_[0]),
		.chany_top_in_169_(cby_2__1__0_chany_out_169_[0]),
		.chany_top_in_171_(cby_2__1__0_chany_out_171_[0]),
		.chany_top_in_173_(cby_2__1__0_chany_out_173_[0]),
		.chany_top_in_175_(cby_2__1__0_chany_out_175_[0]),
		.chany_top_in_177_(cby_2__1__0_chany_out_177_[0]),
		.chany_top_in_179_(cby_2__1__0_chany_out_179_[0]),
		.chany_top_in_181_(cby_2__1__0_chany_out_181_[0]),
		.chany_top_in_183_(cby_2__1__0_chany_out_183_[0]),
		.chany_top_in_185_(cby_2__1__0_chany_out_185_[0]),
		.chany_top_in_187_(cby_2__1__0_chany_out_187_[0]),
		.chany_top_in_189_(cby_2__1__0_chany_out_189_[0]),
		.chany_top_in_191_(cby_2__1__0_chany_out_191_[0]),
		.chany_top_in_193_(cby_2__1__0_chany_out_193_[0]),
		.chany_top_in_195_(cby_2__1__0_chany_out_195_[0]),
		.chany_top_in_197_(cby_2__1__0_chany_out_197_[0]),
		.chany_top_in_199_(cby_2__1__0_chany_out_199_[0]),
		.top_left_grid_pin_44_(grid_clb_1_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_1_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_1_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_1_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_1_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_1_right_width_0_height_0__pin_49_lower[0]),
		.top_left_grid_pin_50_(grid_clb_1_right_width_0_height_0__pin_50_lower[0]),
		.top_left_grid_pin_51_(grid_clb_1_right_width_0_height_0__pin_51_lower[0]),
		.top_left_grid_pin_52_(grid_clb_1_right_width_0_height_0__pin_52_lower[0]),
		.top_left_grid_pin_53_(grid_clb_1_right_width_0_height_0__pin_53_lower[0]),
		.top_right_grid_pin_1_(grid_io_right_0_left_width_0_height_0__pin_1_lower[0]),
		.chanx_left_in_0_(cbx_1__0__1_chanx_out_0_[0]),
		.chanx_left_in_2_(cbx_1__0__1_chanx_out_2_[0]),
		.chanx_left_in_4_(cbx_1__0__1_chanx_out_4_[0]),
		.chanx_left_in_6_(cbx_1__0__1_chanx_out_6_[0]),
		.chanx_left_in_8_(cbx_1__0__1_chanx_out_8_[0]),
		.chanx_left_in_10_(cbx_1__0__1_chanx_out_10_[0]),
		.chanx_left_in_12_(cbx_1__0__1_chanx_out_12_[0]),
		.chanx_left_in_14_(cbx_1__0__1_chanx_out_14_[0]),
		.chanx_left_in_16_(cbx_1__0__1_chanx_out_16_[0]),
		.chanx_left_in_18_(cbx_1__0__1_chanx_out_18_[0]),
		.chanx_left_in_20_(cbx_1__0__1_chanx_out_20_[0]),
		.chanx_left_in_22_(cbx_1__0__1_chanx_out_22_[0]),
		.chanx_left_in_24_(cbx_1__0__1_chanx_out_24_[0]),
		.chanx_left_in_26_(cbx_1__0__1_chanx_out_26_[0]),
		.chanx_left_in_28_(cbx_1__0__1_chanx_out_28_[0]),
		.chanx_left_in_30_(cbx_1__0__1_chanx_out_30_[0]),
		.chanx_left_in_32_(cbx_1__0__1_chanx_out_32_[0]),
		.chanx_left_in_34_(cbx_1__0__1_chanx_out_34_[0]),
		.chanx_left_in_36_(cbx_1__0__1_chanx_out_36_[0]),
		.chanx_left_in_38_(cbx_1__0__1_chanx_out_38_[0]),
		.chanx_left_in_40_(cbx_1__0__1_chanx_out_40_[0]),
		.chanx_left_in_42_(cbx_1__0__1_chanx_out_42_[0]),
		.chanx_left_in_44_(cbx_1__0__1_chanx_out_44_[0]),
		.chanx_left_in_46_(cbx_1__0__1_chanx_out_46_[0]),
		.chanx_left_in_48_(cbx_1__0__1_chanx_out_48_[0]),
		.chanx_left_in_50_(cbx_1__0__1_chanx_out_50_[0]),
		.chanx_left_in_52_(cbx_1__0__1_chanx_out_52_[0]),
		.chanx_left_in_54_(cbx_1__0__1_chanx_out_54_[0]),
		.chanx_left_in_56_(cbx_1__0__1_chanx_out_56_[0]),
		.chanx_left_in_58_(cbx_1__0__1_chanx_out_58_[0]),
		.chanx_left_in_60_(cbx_1__0__1_chanx_out_60_[0]),
		.chanx_left_in_62_(cbx_1__0__1_chanx_out_62_[0]),
		.chanx_left_in_64_(cbx_1__0__1_chanx_out_64_[0]),
		.chanx_left_in_66_(cbx_1__0__1_chanx_out_66_[0]),
		.chanx_left_in_68_(cbx_1__0__1_chanx_out_68_[0]),
		.chanx_left_in_70_(cbx_1__0__1_chanx_out_70_[0]),
		.chanx_left_in_72_(cbx_1__0__1_chanx_out_72_[0]),
		.chanx_left_in_74_(cbx_1__0__1_chanx_out_74_[0]),
		.chanx_left_in_76_(cbx_1__0__1_chanx_out_76_[0]),
		.chanx_left_in_78_(cbx_1__0__1_chanx_out_78_[0]),
		.chanx_left_in_80_(cbx_1__0__1_chanx_out_80_[0]),
		.chanx_left_in_82_(cbx_1__0__1_chanx_out_82_[0]),
		.chanx_left_in_84_(cbx_1__0__1_chanx_out_84_[0]),
		.chanx_left_in_86_(cbx_1__0__1_chanx_out_86_[0]),
		.chanx_left_in_88_(cbx_1__0__1_chanx_out_88_[0]),
		.chanx_left_in_90_(cbx_1__0__1_chanx_out_90_[0]),
		.chanx_left_in_92_(cbx_1__0__1_chanx_out_92_[0]),
		.chanx_left_in_94_(cbx_1__0__1_chanx_out_94_[0]),
		.chanx_left_in_96_(cbx_1__0__1_chanx_out_96_[0]),
		.chanx_left_in_98_(cbx_1__0__1_chanx_out_98_[0]),
		.chanx_left_in_100_(cbx_1__0__1_chanx_out_100_[0]),
		.chanx_left_in_102_(cbx_1__0__1_chanx_out_102_[0]),
		.chanx_left_in_104_(cbx_1__0__1_chanx_out_104_[0]),
		.chanx_left_in_106_(cbx_1__0__1_chanx_out_106_[0]),
		.chanx_left_in_108_(cbx_1__0__1_chanx_out_108_[0]),
		.chanx_left_in_110_(cbx_1__0__1_chanx_out_110_[0]),
		.chanx_left_in_112_(cbx_1__0__1_chanx_out_112_[0]),
		.chanx_left_in_114_(cbx_1__0__1_chanx_out_114_[0]),
		.chanx_left_in_116_(cbx_1__0__1_chanx_out_116_[0]),
		.chanx_left_in_118_(cbx_1__0__1_chanx_out_118_[0]),
		.chanx_left_in_120_(cbx_1__0__1_chanx_out_120_[0]),
		.chanx_left_in_122_(cbx_1__0__1_chanx_out_122_[0]),
		.chanx_left_in_124_(cbx_1__0__1_chanx_out_124_[0]),
		.chanx_left_in_126_(cbx_1__0__1_chanx_out_126_[0]),
		.chanx_left_in_128_(cbx_1__0__1_chanx_out_128_[0]),
		.chanx_left_in_130_(cbx_1__0__1_chanx_out_130_[0]),
		.chanx_left_in_132_(cbx_1__0__1_chanx_out_132_[0]),
		.chanx_left_in_134_(cbx_1__0__1_chanx_out_134_[0]),
		.chanx_left_in_136_(cbx_1__0__1_chanx_out_136_[0]),
		.chanx_left_in_138_(cbx_1__0__1_chanx_out_138_[0]),
		.chanx_left_in_140_(cbx_1__0__1_chanx_out_140_[0]),
		.chanx_left_in_142_(cbx_1__0__1_chanx_out_142_[0]),
		.chanx_left_in_144_(cbx_1__0__1_chanx_out_144_[0]),
		.chanx_left_in_146_(cbx_1__0__1_chanx_out_146_[0]),
		.chanx_left_in_148_(cbx_1__0__1_chanx_out_148_[0]),
		.chanx_left_in_150_(cbx_1__0__1_chanx_out_150_[0]),
		.chanx_left_in_152_(cbx_1__0__1_chanx_out_152_[0]),
		.chanx_left_in_154_(cbx_1__0__1_chanx_out_154_[0]),
		.chanx_left_in_156_(cbx_1__0__1_chanx_out_156_[0]),
		.chanx_left_in_158_(cbx_1__0__1_chanx_out_158_[0]),
		.chanx_left_in_160_(cbx_1__0__1_chanx_out_160_[0]),
		.chanx_left_in_162_(cbx_1__0__1_chanx_out_162_[0]),
		.chanx_left_in_164_(cbx_1__0__1_chanx_out_164_[0]),
		.chanx_left_in_166_(cbx_1__0__1_chanx_out_166_[0]),
		.chanx_left_in_168_(cbx_1__0__1_chanx_out_168_[0]),
		.chanx_left_in_170_(cbx_1__0__1_chanx_out_170_[0]),
		.chanx_left_in_172_(cbx_1__0__1_chanx_out_172_[0]),
		.chanx_left_in_174_(cbx_1__0__1_chanx_out_174_[0]),
		.chanx_left_in_176_(cbx_1__0__1_chanx_out_176_[0]),
		.chanx_left_in_178_(cbx_1__0__1_chanx_out_178_[0]),
		.chanx_left_in_180_(cbx_1__0__1_chanx_out_180_[0]),
		.chanx_left_in_182_(cbx_1__0__1_chanx_out_182_[0]),
		.chanx_left_in_184_(cbx_1__0__1_chanx_out_184_[0]),
		.chanx_left_in_186_(cbx_1__0__1_chanx_out_186_[0]),
		.chanx_left_in_188_(cbx_1__0__1_chanx_out_188_[0]),
		.chanx_left_in_190_(cbx_1__0__1_chanx_out_190_[0]),
		.chanx_left_in_192_(cbx_1__0__1_chanx_out_192_[0]),
		.chanx_left_in_194_(cbx_1__0__1_chanx_out_194_[0]),
		.chanx_left_in_196_(cbx_1__0__1_chanx_out_196_[0]),
		.chanx_left_in_198_(cbx_1__0__1_chanx_out_198_[0]),
		.left_top_grid_pin_54_(grid_clb_1_bottom_width_0_height_0__pin_54_lower[0]),
		.left_top_grid_pin_55_(grid_clb_1_bottom_width_0_height_0__pin_55_lower[0]),
		.left_top_grid_pin_56_(grid_clb_1_bottom_width_0_height_0__pin_56_lower[0]),
		.left_top_grid_pin_57_(grid_clb_1_bottom_width_0_height_0__pin_57_lower[0]),
		.left_top_grid_pin_58_(grid_clb_1_bottom_width_0_height_0__pin_58_lower[0]),
		.left_top_grid_pin_59_(grid_clb_1_bottom_width_0_height_0__pin_59_lower[0]),
		.left_top_grid_pin_60_(grid_clb_1_bottom_width_0_height_0__pin_60_lower[0]),
		.left_top_grid_pin_61_(grid_clb_1_bottom_width_0_height_0__pin_61_lower[0]),
		.left_top_grid_pin_62_(grid_clb_1_bottom_width_0_height_0__pin_62_lower[0]),
		.left_top_grid_pin_63_(grid_clb_1_bottom_width_0_height_0__pin_63_lower[0]),
		.left_top_grid_pin_66_(grid_clb_1_bottom_width_0_height_0__pin_66_lower[0]),
		.left_top_grid_pin_67_(grid_clb_1_bottom_width_0_height_0__pin_67_lower[0]),
		.left_bottom_grid_pin_1_(grid_io_bottom_1_top_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_clb_spypad_0_ccff_tail[0]),
		.chany_top_out_0_(sb_2__0__0_chany_top_out_0_[0]),
		.chany_top_out_2_(sb_2__0__0_chany_top_out_2_[0]),
		.chany_top_out_4_(sb_2__0__0_chany_top_out_4_[0]),
		.chany_top_out_6_(sb_2__0__0_chany_top_out_6_[0]),
		.chany_top_out_8_(sb_2__0__0_chany_top_out_8_[0]),
		.chany_top_out_10_(sb_2__0__0_chany_top_out_10_[0]),
		.chany_top_out_12_(sb_2__0__0_chany_top_out_12_[0]),
		.chany_top_out_14_(sb_2__0__0_chany_top_out_14_[0]),
		.chany_top_out_16_(sb_2__0__0_chany_top_out_16_[0]),
		.chany_top_out_18_(sb_2__0__0_chany_top_out_18_[0]),
		.chany_top_out_20_(sb_2__0__0_chany_top_out_20_[0]),
		.chany_top_out_22_(sb_2__0__0_chany_top_out_22_[0]),
		.chany_top_out_24_(sb_2__0__0_chany_top_out_24_[0]),
		.chany_top_out_26_(sb_2__0__0_chany_top_out_26_[0]),
		.chany_top_out_28_(sb_2__0__0_chany_top_out_28_[0]),
		.chany_top_out_30_(sb_2__0__0_chany_top_out_30_[0]),
		.chany_top_out_32_(sb_2__0__0_chany_top_out_32_[0]),
		.chany_top_out_34_(sb_2__0__0_chany_top_out_34_[0]),
		.chany_top_out_36_(sb_2__0__0_chany_top_out_36_[0]),
		.chany_top_out_38_(sb_2__0__0_chany_top_out_38_[0]),
		.chany_top_out_40_(sb_2__0__0_chany_top_out_40_[0]),
		.chany_top_out_42_(sb_2__0__0_chany_top_out_42_[0]),
		.chany_top_out_44_(sb_2__0__0_chany_top_out_44_[0]),
		.chany_top_out_46_(sb_2__0__0_chany_top_out_46_[0]),
		.chany_top_out_48_(sb_2__0__0_chany_top_out_48_[0]),
		.chany_top_out_50_(sb_2__0__0_chany_top_out_50_[0]),
		.chany_top_out_52_(sb_2__0__0_chany_top_out_52_[0]),
		.chany_top_out_54_(sb_2__0__0_chany_top_out_54_[0]),
		.chany_top_out_56_(sb_2__0__0_chany_top_out_56_[0]),
		.chany_top_out_58_(sb_2__0__0_chany_top_out_58_[0]),
		.chany_top_out_60_(sb_2__0__0_chany_top_out_60_[0]),
		.chany_top_out_62_(sb_2__0__0_chany_top_out_62_[0]),
		.chany_top_out_64_(sb_2__0__0_chany_top_out_64_[0]),
		.chany_top_out_66_(sb_2__0__0_chany_top_out_66_[0]),
		.chany_top_out_68_(sb_2__0__0_chany_top_out_68_[0]),
		.chany_top_out_70_(sb_2__0__0_chany_top_out_70_[0]),
		.chany_top_out_72_(sb_2__0__0_chany_top_out_72_[0]),
		.chany_top_out_74_(sb_2__0__0_chany_top_out_74_[0]),
		.chany_top_out_76_(sb_2__0__0_chany_top_out_76_[0]),
		.chany_top_out_78_(sb_2__0__0_chany_top_out_78_[0]),
		.chany_top_out_80_(sb_2__0__0_chany_top_out_80_[0]),
		.chany_top_out_82_(sb_2__0__0_chany_top_out_82_[0]),
		.chany_top_out_84_(sb_2__0__0_chany_top_out_84_[0]),
		.chany_top_out_86_(sb_2__0__0_chany_top_out_86_[0]),
		.chany_top_out_88_(sb_2__0__0_chany_top_out_88_[0]),
		.chany_top_out_90_(sb_2__0__0_chany_top_out_90_[0]),
		.chany_top_out_92_(sb_2__0__0_chany_top_out_92_[0]),
		.chany_top_out_94_(sb_2__0__0_chany_top_out_94_[0]),
		.chany_top_out_96_(sb_2__0__0_chany_top_out_96_[0]),
		.chany_top_out_98_(sb_2__0__0_chany_top_out_98_[0]),
		.chany_top_out_100_(sb_2__0__0_chany_top_out_100_[0]),
		.chany_top_out_102_(sb_2__0__0_chany_top_out_102_[0]),
		.chany_top_out_104_(sb_2__0__0_chany_top_out_104_[0]),
		.chany_top_out_106_(sb_2__0__0_chany_top_out_106_[0]),
		.chany_top_out_108_(sb_2__0__0_chany_top_out_108_[0]),
		.chany_top_out_110_(sb_2__0__0_chany_top_out_110_[0]),
		.chany_top_out_112_(sb_2__0__0_chany_top_out_112_[0]),
		.chany_top_out_114_(sb_2__0__0_chany_top_out_114_[0]),
		.chany_top_out_116_(sb_2__0__0_chany_top_out_116_[0]),
		.chany_top_out_118_(sb_2__0__0_chany_top_out_118_[0]),
		.chany_top_out_120_(sb_2__0__0_chany_top_out_120_[0]),
		.chany_top_out_122_(sb_2__0__0_chany_top_out_122_[0]),
		.chany_top_out_124_(sb_2__0__0_chany_top_out_124_[0]),
		.chany_top_out_126_(sb_2__0__0_chany_top_out_126_[0]),
		.chany_top_out_128_(sb_2__0__0_chany_top_out_128_[0]),
		.chany_top_out_130_(sb_2__0__0_chany_top_out_130_[0]),
		.chany_top_out_132_(sb_2__0__0_chany_top_out_132_[0]),
		.chany_top_out_134_(sb_2__0__0_chany_top_out_134_[0]),
		.chany_top_out_136_(sb_2__0__0_chany_top_out_136_[0]),
		.chany_top_out_138_(sb_2__0__0_chany_top_out_138_[0]),
		.chany_top_out_140_(sb_2__0__0_chany_top_out_140_[0]),
		.chany_top_out_142_(sb_2__0__0_chany_top_out_142_[0]),
		.chany_top_out_144_(sb_2__0__0_chany_top_out_144_[0]),
		.chany_top_out_146_(sb_2__0__0_chany_top_out_146_[0]),
		.chany_top_out_148_(sb_2__0__0_chany_top_out_148_[0]),
		.chany_top_out_150_(sb_2__0__0_chany_top_out_150_[0]),
		.chany_top_out_152_(sb_2__0__0_chany_top_out_152_[0]),
		.chany_top_out_154_(sb_2__0__0_chany_top_out_154_[0]),
		.chany_top_out_156_(sb_2__0__0_chany_top_out_156_[0]),
		.chany_top_out_158_(sb_2__0__0_chany_top_out_158_[0]),
		.chany_top_out_160_(sb_2__0__0_chany_top_out_160_[0]),
		.chany_top_out_162_(sb_2__0__0_chany_top_out_162_[0]),
		.chany_top_out_164_(sb_2__0__0_chany_top_out_164_[0]),
		.chany_top_out_166_(sb_2__0__0_chany_top_out_166_[0]),
		.chany_top_out_168_(sb_2__0__0_chany_top_out_168_[0]),
		.chany_top_out_170_(sb_2__0__0_chany_top_out_170_[0]),
		.chany_top_out_172_(sb_2__0__0_chany_top_out_172_[0]),
		.chany_top_out_174_(sb_2__0__0_chany_top_out_174_[0]),
		.chany_top_out_176_(sb_2__0__0_chany_top_out_176_[0]),
		.chany_top_out_178_(sb_2__0__0_chany_top_out_178_[0]),
		.chany_top_out_180_(sb_2__0__0_chany_top_out_180_[0]),
		.chany_top_out_182_(sb_2__0__0_chany_top_out_182_[0]),
		.chany_top_out_184_(sb_2__0__0_chany_top_out_184_[0]),
		.chany_top_out_186_(sb_2__0__0_chany_top_out_186_[0]),
		.chany_top_out_188_(sb_2__0__0_chany_top_out_188_[0]),
		.chany_top_out_190_(sb_2__0__0_chany_top_out_190_[0]),
		.chany_top_out_192_(sb_2__0__0_chany_top_out_192_[0]),
		.chany_top_out_194_(sb_2__0__0_chany_top_out_194_[0]),
		.chany_top_out_196_(sb_2__0__0_chany_top_out_196_[0]),
		.chany_top_out_198_(sb_2__0__0_chany_top_out_198_[0]),
		.chanx_left_out_1_(sb_2__0__0_chanx_left_out_1_[0]),
		.chanx_left_out_3_(sb_2__0__0_chanx_left_out_3_[0]),
		.chanx_left_out_5_(sb_2__0__0_chanx_left_out_5_[0]),
		.chanx_left_out_7_(sb_2__0__0_chanx_left_out_7_[0]),
		.chanx_left_out_9_(sb_2__0__0_chanx_left_out_9_[0]),
		.chanx_left_out_11_(sb_2__0__0_chanx_left_out_11_[0]),
		.chanx_left_out_13_(sb_2__0__0_chanx_left_out_13_[0]),
		.chanx_left_out_15_(sb_2__0__0_chanx_left_out_15_[0]),
		.chanx_left_out_17_(sb_2__0__0_chanx_left_out_17_[0]),
		.chanx_left_out_19_(sb_2__0__0_chanx_left_out_19_[0]),
		.chanx_left_out_21_(sb_2__0__0_chanx_left_out_21_[0]),
		.chanx_left_out_23_(sb_2__0__0_chanx_left_out_23_[0]),
		.chanx_left_out_25_(sb_2__0__0_chanx_left_out_25_[0]),
		.chanx_left_out_27_(sb_2__0__0_chanx_left_out_27_[0]),
		.chanx_left_out_29_(sb_2__0__0_chanx_left_out_29_[0]),
		.chanx_left_out_31_(sb_2__0__0_chanx_left_out_31_[0]),
		.chanx_left_out_33_(sb_2__0__0_chanx_left_out_33_[0]),
		.chanx_left_out_35_(sb_2__0__0_chanx_left_out_35_[0]),
		.chanx_left_out_37_(sb_2__0__0_chanx_left_out_37_[0]),
		.chanx_left_out_39_(sb_2__0__0_chanx_left_out_39_[0]),
		.chanx_left_out_41_(sb_2__0__0_chanx_left_out_41_[0]),
		.chanx_left_out_43_(sb_2__0__0_chanx_left_out_43_[0]),
		.chanx_left_out_45_(sb_2__0__0_chanx_left_out_45_[0]),
		.chanx_left_out_47_(sb_2__0__0_chanx_left_out_47_[0]),
		.chanx_left_out_49_(sb_2__0__0_chanx_left_out_49_[0]),
		.chanx_left_out_51_(sb_2__0__0_chanx_left_out_51_[0]),
		.chanx_left_out_53_(sb_2__0__0_chanx_left_out_53_[0]),
		.chanx_left_out_55_(sb_2__0__0_chanx_left_out_55_[0]),
		.chanx_left_out_57_(sb_2__0__0_chanx_left_out_57_[0]),
		.chanx_left_out_59_(sb_2__0__0_chanx_left_out_59_[0]),
		.chanx_left_out_61_(sb_2__0__0_chanx_left_out_61_[0]),
		.chanx_left_out_63_(sb_2__0__0_chanx_left_out_63_[0]),
		.chanx_left_out_65_(sb_2__0__0_chanx_left_out_65_[0]),
		.chanx_left_out_67_(sb_2__0__0_chanx_left_out_67_[0]),
		.chanx_left_out_69_(sb_2__0__0_chanx_left_out_69_[0]),
		.chanx_left_out_71_(sb_2__0__0_chanx_left_out_71_[0]),
		.chanx_left_out_73_(sb_2__0__0_chanx_left_out_73_[0]),
		.chanx_left_out_75_(sb_2__0__0_chanx_left_out_75_[0]),
		.chanx_left_out_77_(sb_2__0__0_chanx_left_out_77_[0]),
		.chanx_left_out_79_(sb_2__0__0_chanx_left_out_79_[0]),
		.chanx_left_out_81_(sb_2__0__0_chanx_left_out_81_[0]),
		.chanx_left_out_83_(sb_2__0__0_chanx_left_out_83_[0]),
		.chanx_left_out_85_(sb_2__0__0_chanx_left_out_85_[0]),
		.chanx_left_out_87_(sb_2__0__0_chanx_left_out_87_[0]),
		.chanx_left_out_89_(sb_2__0__0_chanx_left_out_89_[0]),
		.chanx_left_out_91_(sb_2__0__0_chanx_left_out_91_[0]),
		.chanx_left_out_93_(sb_2__0__0_chanx_left_out_93_[0]),
		.chanx_left_out_95_(sb_2__0__0_chanx_left_out_95_[0]),
		.chanx_left_out_97_(sb_2__0__0_chanx_left_out_97_[0]),
		.chanx_left_out_99_(sb_2__0__0_chanx_left_out_99_[0]),
		.chanx_left_out_101_(sb_2__0__0_chanx_left_out_101_[0]),
		.chanx_left_out_103_(sb_2__0__0_chanx_left_out_103_[0]),
		.chanx_left_out_105_(sb_2__0__0_chanx_left_out_105_[0]),
		.chanx_left_out_107_(sb_2__0__0_chanx_left_out_107_[0]),
		.chanx_left_out_109_(sb_2__0__0_chanx_left_out_109_[0]),
		.chanx_left_out_111_(sb_2__0__0_chanx_left_out_111_[0]),
		.chanx_left_out_113_(sb_2__0__0_chanx_left_out_113_[0]),
		.chanx_left_out_115_(sb_2__0__0_chanx_left_out_115_[0]),
		.chanx_left_out_117_(sb_2__0__0_chanx_left_out_117_[0]),
		.chanx_left_out_119_(sb_2__0__0_chanx_left_out_119_[0]),
		.chanx_left_out_121_(sb_2__0__0_chanx_left_out_121_[0]),
		.chanx_left_out_123_(sb_2__0__0_chanx_left_out_123_[0]),
		.chanx_left_out_125_(sb_2__0__0_chanx_left_out_125_[0]),
		.chanx_left_out_127_(sb_2__0__0_chanx_left_out_127_[0]),
		.chanx_left_out_129_(sb_2__0__0_chanx_left_out_129_[0]),
		.chanx_left_out_131_(sb_2__0__0_chanx_left_out_131_[0]),
		.chanx_left_out_133_(sb_2__0__0_chanx_left_out_133_[0]),
		.chanx_left_out_135_(sb_2__0__0_chanx_left_out_135_[0]),
		.chanx_left_out_137_(sb_2__0__0_chanx_left_out_137_[0]),
		.chanx_left_out_139_(sb_2__0__0_chanx_left_out_139_[0]),
		.chanx_left_out_141_(sb_2__0__0_chanx_left_out_141_[0]),
		.chanx_left_out_143_(sb_2__0__0_chanx_left_out_143_[0]),
		.chanx_left_out_145_(sb_2__0__0_chanx_left_out_145_[0]),
		.chanx_left_out_147_(sb_2__0__0_chanx_left_out_147_[0]),
		.chanx_left_out_149_(sb_2__0__0_chanx_left_out_149_[0]),
		.chanx_left_out_151_(sb_2__0__0_chanx_left_out_151_[0]),
		.chanx_left_out_153_(sb_2__0__0_chanx_left_out_153_[0]),
		.chanx_left_out_155_(sb_2__0__0_chanx_left_out_155_[0]),
		.chanx_left_out_157_(sb_2__0__0_chanx_left_out_157_[0]),
		.chanx_left_out_159_(sb_2__0__0_chanx_left_out_159_[0]),
		.chanx_left_out_161_(sb_2__0__0_chanx_left_out_161_[0]),
		.chanx_left_out_163_(sb_2__0__0_chanx_left_out_163_[0]),
		.chanx_left_out_165_(sb_2__0__0_chanx_left_out_165_[0]),
		.chanx_left_out_167_(sb_2__0__0_chanx_left_out_167_[0]),
		.chanx_left_out_169_(sb_2__0__0_chanx_left_out_169_[0]),
		.chanx_left_out_171_(sb_2__0__0_chanx_left_out_171_[0]),
		.chanx_left_out_173_(sb_2__0__0_chanx_left_out_173_[0]),
		.chanx_left_out_175_(sb_2__0__0_chanx_left_out_175_[0]),
		.chanx_left_out_177_(sb_2__0__0_chanx_left_out_177_[0]),
		.chanx_left_out_179_(sb_2__0__0_chanx_left_out_179_[0]),
		.chanx_left_out_181_(sb_2__0__0_chanx_left_out_181_[0]),
		.chanx_left_out_183_(sb_2__0__0_chanx_left_out_183_[0]),
		.chanx_left_out_185_(sb_2__0__0_chanx_left_out_185_[0]),
		.chanx_left_out_187_(sb_2__0__0_chanx_left_out_187_[0]),
		.chanx_left_out_189_(sb_2__0__0_chanx_left_out_189_[0]),
		.chanx_left_out_191_(sb_2__0__0_chanx_left_out_191_[0]),
		.chanx_left_out_193_(sb_2__0__0_chanx_left_out_193_[0]),
		.chanx_left_out_195_(sb_2__0__0_chanx_left_out_195_[0]),
		.chanx_left_out_197_(sb_2__0__0_chanx_left_out_197_[0]),
		.chanx_left_out_199_(sb_2__0__0_chanx_left_out_199_[0]),
		.ccff_tail(sb_2__0__0_ccff_tail[0]));

	sb_2__1_ sb_2__1_ (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.chany_top_in_1_(cby_2__1__1_chany_out_1_[0]),
		.chany_top_in_3_(cby_2__1__1_chany_out_3_[0]),
		.chany_top_in_5_(cby_2__1__1_chany_out_5_[0]),
		.chany_top_in_7_(cby_2__1__1_chany_out_7_[0]),
		.chany_top_in_9_(cby_2__1__1_chany_out_9_[0]),
		.chany_top_in_11_(cby_2__1__1_chany_out_11_[0]),
		.chany_top_in_13_(cby_2__1__1_chany_out_13_[0]),
		.chany_top_in_15_(cby_2__1__1_chany_out_15_[0]),
		.chany_top_in_17_(cby_2__1__1_chany_out_17_[0]),
		.chany_top_in_19_(cby_2__1__1_chany_out_19_[0]),
		.chany_top_in_21_(cby_2__1__1_chany_out_21_[0]),
		.chany_top_in_23_(cby_2__1__1_chany_out_23_[0]),
		.chany_top_in_25_(cby_2__1__1_chany_out_25_[0]),
		.chany_top_in_27_(cby_2__1__1_chany_out_27_[0]),
		.chany_top_in_29_(cby_2__1__1_chany_out_29_[0]),
		.chany_top_in_31_(cby_2__1__1_chany_out_31_[0]),
		.chany_top_in_33_(cby_2__1__1_chany_out_33_[0]),
		.chany_top_in_35_(cby_2__1__1_chany_out_35_[0]),
		.chany_top_in_37_(cby_2__1__1_chany_out_37_[0]),
		.chany_top_in_39_(cby_2__1__1_chany_out_39_[0]),
		.chany_top_in_41_(cby_2__1__1_chany_out_41_[0]),
		.chany_top_in_43_(cby_2__1__1_chany_out_43_[0]),
		.chany_top_in_45_(cby_2__1__1_chany_out_45_[0]),
		.chany_top_in_47_(cby_2__1__1_chany_out_47_[0]),
		.chany_top_in_49_(cby_2__1__1_chany_out_49_[0]),
		.chany_top_in_51_(cby_2__1__1_chany_out_51_[0]),
		.chany_top_in_53_(cby_2__1__1_chany_out_53_[0]),
		.chany_top_in_55_(cby_2__1__1_chany_out_55_[0]),
		.chany_top_in_57_(cby_2__1__1_chany_out_57_[0]),
		.chany_top_in_59_(cby_2__1__1_chany_out_59_[0]),
		.chany_top_in_61_(cby_2__1__1_chany_out_61_[0]),
		.chany_top_in_63_(cby_2__1__1_chany_out_63_[0]),
		.chany_top_in_65_(cby_2__1__1_chany_out_65_[0]),
		.chany_top_in_67_(cby_2__1__1_chany_out_67_[0]),
		.chany_top_in_69_(cby_2__1__1_chany_out_69_[0]),
		.chany_top_in_71_(cby_2__1__1_chany_out_71_[0]),
		.chany_top_in_73_(cby_2__1__1_chany_out_73_[0]),
		.chany_top_in_75_(cby_2__1__1_chany_out_75_[0]),
		.chany_top_in_77_(cby_2__1__1_chany_out_77_[0]),
		.chany_top_in_79_(cby_2__1__1_chany_out_79_[0]),
		.chany_top_in_81_(cby_2__1__1_chany_out_81_[0]),
		.chany_top_in_83_(cby_2__1__1_chany_out_83_[0]),
		.chany_top_in_85_(cby_2__1__1_chany_out_85_[0]),
		.chany_top_in_87_(cby_2__1__1_chany_out_87_[0]),
		.chany_top_in_89_(cby_2__1__1_chany_out_89_[0]),
		.chany_top_in_91_(cby_2__1__1_chany_out_91_[0]),
		.chany_top_in_93_(cby_2__1__1_chany_out_93_[0]),
		.chany_top_in_95_(cby_2__1__1_chany_out_95_[0]),
		.chany_top_in_97_(cby_2__1__1_chany_out_97_[0]),
		.chany_top_in_99_(cby_2__1__1_chany_out_99_[0]),
		.chany_top_in_101_(cby_2__1__1_chany_out_101_[0]),
		.chany_top_in_103_(cby_2__1__1_chany_out_103_[0]),
		.chany_top_in_105_(cby_2__1__1_chany_out_105_[0]),
		.chany_top_in_107_(cby_2__1__1_chany_out_107_[0]),
		.chany_top_in_109_(cby_2__1__1_chany_out_109_[0]),
		.chany_top_in_111_(cby_2__1__1_chany_out_111_[0]),
		.chany_top_in_113_(cby_2__1__1_chany_out_113_[0]),
		.chany_top_in_115_(cby_2__1__1_chany_out_115_[0]),
		.chany_top_in_117_(cby_2__1__1_chany_out_117_[0]),
		.chany_top_in_119_(cby_2__1__1_chany_out_119_[0]),
		.chany_top_in_121_(cby_2__1__1_chany_out_121_[0]),
		.chany_top_in_123_(cby_2__1__1_chany_out_123_[0]),
		.chany_top_in_125_(cby_2__1__1_chany_out_125_[0]),
		.chany_top_in_127_(cby_2__1__1_chany_out_127_[0]),
		.chany_top_in_129_(cby_2__1__1_chany_out_129_[0]),
		.chany_top_in_131_(cby_2__1__1_chany_out_131_[0]),
		.chany_top_in_133_(cby_2__1__1_chany_out_133_[0]),
		.chany_top_in_135_(cby_2__1__1_chany_out_135_[0]),
		.chany_top_in_137_(cby_2__1__1_chany_out_137_[0]),
		.chany_top_in_139_(cby_2__1__1_chany_out_139_[0]),
		.chany_top_in_141_(cby_2__1__1_chany_out_141_[0]),
		.chany_top_in_143_(cby_2__1__1_chany_out_143_[0]),
		.chany_top_in_145_(cby_2__1__1_chany_out_145_[0]),
		.chany_top_in_147_(cby_2__1__1_chany_out_147_[0]),
		.chany_top_in_149_(cby_2__1__1_chany_out_149_[0]),
		.chany_top_in_151_(cby_2__1__1_chany_out_151_[0]),
		.chany_top_in_153_(cby_2__1__1_chany_out_153_[0]),
		.chany_top_in_155_(cby_2__1__1_chany_out_155_[0]),
		.chany_top_in_157_(cby_2__1__1_chany_out_157_[0]),
		.chany_top_in_159_(cby_2__1__1_chany_out_159_[0]),
		.chany_top_in_161_(cby_2__1__1_chany_out_161_[0]),
		.chany_top_in_163_(cby_2__1__1_chany_out_163_[0]),
		.chany_top_in_165_(cby_2__1__1_chany_out_165_[0]),
		.chany_top_in_167_(cby_2__1__1_chany_out_167_[0]),
		.chany_top_in_169_(cby_2__1__1_chany_out_169_[0]),
		.chany_top_in_171_(cby_2__1__1_chany_out_171_[0]),
		.chany_top_in_173_(cby_2__1__1_chany_out_173_[0]),
		.chany_top_in_175_(cby_2__1__1_chany_out_175_[0]),
		.chany_top_in_177_(cby_2__1__1_chany_out_177_[0]),
		.chany_top_in_179_(cby_2__1__1_chany_out_179_[0]),
		.chany_top_in_181_(cby_2__1__1_chany_out_181_[0]),
		.chany_top_in_183_(cby_2__1__1_chany_out_183_[0]),
		.chany_top_in_185_(cby_2__1__1_chany_out_185_[0]),
		.chany_top_in_187_(cby_2__1__1_chany_out_187_[0]),
		.chany_top_in_189_(cby_2__1__1_chany_out_189_[0]),
		.chany_top_in_191_(cby_2__1__1_chany_out_191_[0]),
		.chany_top_in_193_(cby_2__1__1_chany_out_193_[0]),
		.chany_top_in_195_(cby_2__1__1_chany_out_195_[0]),
		.chany_top_in_197_(cby_2__1__1_chany_out_197_[0]),
		.chany_top_in_199_(cby_2__1__1_chany_out_199_[0]),
		.top_left_grid_pin_44_(grid_clb_2_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_2_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_2_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_2_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_2_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_2_right_width_0_height_0__pin_49_lower[0]),
		.top_left_grid_pin_50_(grid_clb_2_right_width_0_height_0__pin_50_lower[0]),
		.top_left_grid_pin_51_(grid_clb_2_right_width_0_height_0__pin_51_lower[0]),
		.top_left_grid_pin_52_(grid_clb_2_right_width_0_height_0__pin_52_lower[0]),
		.top_left_grid_pin_53_(grid_clb_2_right_width_0_height_0__pin_53_lower[0]),
		.top_right_grid_pin_1_(grid_io_right_1_left_width_0_height_0__pin_1_lower[0]),
		.chany_bottom_in_0_(cby_2__1__0_chany_out_0_[0]),
		.chany_bottom_in_2_(cby_2__1__0_chany_out_2_[0]),
		.chany_bottom_in_4_(cby_2__1__0_chany_out_4_[0]),
		.chany_bottom_in_6_(cby_2__1__0_chany_out_6_[0]),
		.chany_bottom_in_8_(cby_2__1__0_chany_out_8_[0]),
		.chany_bottom_in_10_(cby_2__1__0_chany_out_10_[0]),
		.chany_bottom_in_12_(cby_2__1__0_chany_out_12_[0]),
		.chany_bottom_in_14_(cby_2__1__0_chany_out_14_[0]),
		.chany_bottom_in_16_(cby_2__1__0_chany_out_16_[0]),
		.chany_bottom_in_18_(cby_2__1__0_chany_out_18_[0]),
		.chany_bottom_in_20_(cby_2__1__0_chany_out_20_[0]),
		.chany_bottom_in_22_(cby_2__1__0_chany_out_22_[0]),
		.chany_bottom_in_24_(cby_2__1__0_chany_out_24_[0]),
		.chany_bottom_in_26_(cby_2__1__0_chany_out_26_[0]),
		.chany_bottom_in_28_(cby_2__1__0_chany_out_28_[0]),
		.chany_bottom_in_30_(cby_2__1__0_chany_out_30_[0]),
		.chany_bottom_in_32_(cby_2__1__0_chany_out_32_[0]),
		.chany_bottom_in_34_(cby_2__1__0_chany_out_34_[0]),
		.chany_bottom_in_36_(cby_2__1__0_chany_out_36_[0]),
		.chany_bottom_in_38_(cby_2__1__0_chany_out_38_[0]),
		.chany_bottom_in_40_(cby_2__1__0_chany_out_40_[0]),
		.chany_bottom_in_42_(cby_2__1__0_chany_out_42_[0]),
		.chany_bottom_in_44_(cby_2__1__0_chany_out_44_[0]),
		.chany_bottom_in_46_(cby_2__1__0_chany_out_46_[0]),
		.chany_bottom_in_48_(cby_2__1__0_chany_out_48_[0]),
		.chany_bottom_in_50_(cby_2__1__0_chany_out_50_[0]),
		.chany_bottom_in_52_(cby_2__1__0_chany_out_52_[0]),
		.chany_bottom_in_54_(cby_2__1__0_chany_out_54_[0]),
		.chany_bottom_in_56_(cby_2__1__0_chany_out_56_[0]),
		.chany_bottom_in_58_(cby_2__1__0_chany_out_58_[0]),
		.chany_bottom_in_60_(cby_2__1__0_chany_out_60_[0]),
		.chany_bottom_in_62_(cby_2__1__0_chany_out_62_[0]),
		.chany_bottom_in_64_(cby_2__1__0_chany_out_64_[0]),
		.chany_bottom_in_66_(cby_2__1__0_chany_out_66_[0]),
		.chany_bottom_in_68_(cby_2__1__0_chany_out_68_[0]),
		.chany_bottom_in_70_(cby_2__1__0_chany_out_70_[0]),
		.chany_bottom_in_72_(cby_2__1__0_chany_out_72_[0]),
		.chany_bottom_in_74_(cby_2__1__0_chany_out_74_[0]),
		.chany_bottom_in_76_(cby_2__1__0_chany_out_76_[0]),
		.chany_bottom_in_78_(cby_2__1__0_chany_out_78_[0]),
		.chany_bottom_in_80_(cby_2__1__0_chany_out_80_[0]),
		.chany_bottom_in_82_(cby_2__1__0_chany_out_82_[0]),
		.chany_bottom_in_84_(cby_2__1__0_chany_out_84_[0]),
		.chany_bottom_in_86_(cby_2__1__0_chany_out_86_[0]),
		.chany_bottom_in_88_(cby_2__1__0_chany_out_88_[0]),
		.chany_bottom_in_90_(cby_2__1__0_chany_out_90_[0]),
		.chany_bottom_in_92_(cby_2__1__0_chany_out_92_[0]),
		.chany_bottom_in_94_(cby_2__1__0_chany_out_94_[0]),
		.chany_bottom_in_96_(cby_2__1__0_chany_out_96_[0]),
		.chany_bottom_in_98_(cby_2__1__0_chany_out_98_[0]),
		.chany_bottom_in_100_(cby_2__1__0_chany_out_100_[0]),
		.chany_bottom_in_102_(cby_2__1__0_chany_out_102_[0]),
		.chany_bottom_in_104_(cby_2__1__0_chany_out_104_[0]),
		.chany_bottom_in_106_(cby_2__1__0_chany_out_106_[0]),
		.chany_bottom_in_108_(cby_2__1__0_chany_out_108_[0]),
		.chany_bottom_in_110_(cby_2__1__0_chany_out_110_[0]),
		.chany_bottom_in_112_(cby_2__1__0_chany_out_112_[0]),
		.chany_bottom_in_114_(cby_2__1__0_chany_out_114_[0]),
		.chany_bottom_in_116_(cby_2__1__0_chany_out_116_[0]),
		.chany_bottom_in_118_(cby_2__1__0_chany_out_118_[0]),
		.chany_bottom_in_120_(cby_2__1__0_chany_out_120_[0]),
		.chany_bottom_in_122_(cby_2__1__0_chany_out_122_[0]),
		.chany_bottom_in_124_(cby_2__1__0_chany_out_124_[0]),
		.chany_bottom_in_126_(cby_2__1__0_chany_out_126_[0]),
		.chany_bottom_in_128_(cby_2__1__0_chany_out_128_[0]),
		.chany_bottom_in_130_(cby_2__1__0_chany_out_130_[0]),
		.chany_bottom_in_132_(cby_2__1__0_chany_out_132_[0]),
		.chany_bottom_in_134_(cby_2__1__0_chany_out_134_[0]),
		.chany_bottom_in_136_(cby_2__1__0_chany_out_136_[0]),
		.chany_bottom_in_138_(cby_2__1__0_chany_out_138_[0]),
		.chany_bottom_in_140_(cby_2__1__0_chany_out_140_[0]),
		.chany_bottom_in_142_(cby_2__1__0_chany_out_142_[0]),
		.chany_bottom_in_144_(cby_2__1__0_chany_out_144_[0]),
		.chany_bottom_in_146_(cby_2__1__0_chany_out_146_[0]),
		.chany_bottom_in_148_(cby_2__1__0_chany_out_148_[0]),
		.chany_bottom_in_150_(cby_2__1__0_chany_out_150_[0]),
		.chany_bottom_in_152_(cby_2__1__0_chany_out_152_[0]),
		.chany_bottom_in_154_(cby_2__1__0_chany_out_154_[0]),
		.chany_bottom_in_156_(cby_2__1__0_chany_out_156_[0]),
		.chany_bottom_in_158_(cby_2__1__0_chany_out_158_[0]),
		.chany_bottom_in_160_(cby_2__1__0_chany_out_160_[0]),
		.chany_bottom_in_162_(cby_2__1__0_chany_out_162_[0]),
		.chany_bottom_in_164_(cby_2__1__0_chany_out_164_[0]),
		.chany_bottom_in_166_(cby_2__1__0_chany_out_166_[0]),
		.chany_bottom_in_168_(cby_2__1__0_chany_out_168_[0]),
		.chany_bottom_in_170_(cby_2__1__0_chany_out_170_[0]),
		.chany_bottom_in_172_(cby_2__1__0_chany_out_172_[0]),
		.chany_bottom_in_174_(cby_2__1__0_chany_out_174_[0]),
		.chany_bottom_in_176_(cby_2__1__0_chany_out_176_[0]),
		.chany_bottom_in_178_(cby_2__1__0_chany_out_178_[0]),
		.chany_bottom_in_180_(cby_2__1__0_chany_out_180_[0]),
		.chany_bottom_in_182_(cby_2__1__0_chany_out_182_[0]),
		.chany_bottom_in_184_(cby_2__1__0_chany_out_184_[0]),
		.chany_bottom_in_186_(cby_2__1__0_chany_out_186_[0]),
		.chany_bottom_in_188_(cby_2__1__0_chany_out_188_[0]),
		.chany_bottom_in_190_(cby_2__1__0_chany_out_190_[0]),
		.chany_bottom_in_192_(cby_2__1__0_chany_out_192_[0]),
		.chany_bottom_in_194_(cby_2__1__0_chany_out_194_[0]),
		.chany_bottom_in_196_(cby_2__1__0_chany_out_196_[0]),
		.chany_bottom_in_198_(cby_2__1__0_chany_out_198_[0]),
		.bottom_right_grid_pin_1_(grid_io_right_0_left_width_0_height_0__pin_1_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_1_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_1_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_1_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_1_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_1_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_1_right_width_0_height_0__pin_49_upper[0]),
		.bottom_left_grid_pin_50_(grid_clb_1_right_width_0_height_0__pin_50_upper[0]),
		.bottom_left_grid_pin_51_(grid_clb_1_right_width_0_height_0__pin_51_upper[0]),
		.bottom_left_grid_pin_52_(grid_clb_1_right_width_0_height_0__pin_52_upper[0]),
		.bottom_left_grid_pin_53_(grid_clb_1_right_width_0_height_0__pin_53_upper[0]),
		.chanx_left_in_0_(cbx_1__1__1_chanx_out_0_[0]),
		.chanx_left_in_2_(cbx_1__1__1_chanx_out_2_[0]),
		.chanx_left_in_4_(cbx_1__1__1_chanx_out_4_[0]),
		.chanx_left_in_6_(cbx_1__1__1_chanx_out_6_[0]),
		.chanx_left_in_8_(cbx_1__1__1_chanx_out_8_[0]),
		.chanx_left_in_10_(cbx_1__1__1_chanx_out_10_[0]),
		.chanx_left_in_12_(cbx_1__1__1_chanx_out_12_[0]),
		.chanx_left_in_14_(cbx_1__1__1_chanx_out_14_[0]),
		.chanx_left_in_16_(cbx_1__1__1_chanx_out_16_[0]),
		.chanx_left_in_18_(cbx_1__1__1_chanx_out_18_[0]),
		.chanx_left_in_20_(cbx_1__1__1_chanx_out_20_[0]),
		.chanx_left_in_22_(cbx_1__1__1_chanx_out_22_[0]),
		.chanx_left_in_24_(cbx_1__1__1_chanx_out_24_[0]),
		.chanx_left_in_26_(cbx_1__1__1_chanx_out_26_[0]),
		.chanx_left_in_28_(cbx_1__1__1_chanx_out_28_[0]),
		.chanx_left_in_30_(cbx_1__1__1_chanx_out_30_[0]),
		.chanx_left_in_32_(cbx_1__1__1_chanx_out_32_[0]),
		.chanx_left_in_34_(cbx_1__1__1_chanx_out_34_[0]),
		.chanx_left_in_36_(cbx_1__1__1_chanx_out_36_[0]),
		.chanx_left_in_38_(cbx_1__1__1_chanx_out_38_[0]),
		.chanx_left_in_40_(cbx_1__1__1_chanx_out_40_[0]),
		.chanx_left_in_42_(cbx_1__1__1_chanx_out_42_[0]),
		.chanx_left_in_44_(cbx_1__1__1_chanx_out_44_[0]),
		.chanx_left_in_46_(cbx_1__1__1_chanx_out_46_[0]),
		.chanx_left_in_48_(cbx_1__1__1_chanx_out_48_[0]),
		.chanx_left_in_50_(cbx_1__1__1_chanx_out_50_[0]),
		.chanx_left_in_52_(cbx_1__1__1_chanx_out_52_[0]),
		.chanx_left_in_54_(cbx_1__1__1_chanx_out_54_[0]),
		.chanx_left_in_56_(cbx_1__1__1_chanx_out_56_[0]),
		.chanx_left_in_58_(cbx_1__1__1_chanx_out_58_[0]),
		.chanx_left_in_60_(cbx_1__1__1_chanx_out_60_[0]),
		.chanx_left_in_62_(cbx_1__1__1_chanx_out_62_[0]),
		.chanx_left_in_64_(cbx_1__1__1_chanx_out_64_[0]),
		.chanx_left_in_66_(cbx_1__1__1_chanx_out_66_[0]),
		.chanx_left_in_68_(cbx_1__1__1_chanx_out_68_[0]),
		.chanx_left_in_70_(cbx_1__1__1_chanx_out_70_[0]),
		.chanx_left_in_72_(cbx_1__1__1_chanx_out_72_[0]),
		.chanx_left_in_74_(cbx_1__1__1_chanx_out_74_[0]),
		.chanx_left_in_76_(cbx_1__1__1_chanx_out_76_[0]),
		.chanx_left_in_78_(cbx_1__1__1_chanx_out_78_[0]),
		.chanx_left_in_80_(cbx_1__1__1_chanx_out_80_[0]),
		.chanx_left_in_82_(cbx_1__1__1_chanx_out_82_[0]),
		.chanx_left_in_84_(cbx_1__1__1_chanx_out_84_[0]),
		.chanx_left_in_86_(cbx_1__1__1_chanx_out_86_[0]),
		.chanx_left_in_88_(cbx_1__1__1_chanx_out_88_[0]),
		.chanx_left_in_90_(cbx_1__1__1_chanx_out_90_[0]),
		.chanx_left_in_92_(cbx_1__1__1_chanx_out_92_[0]),
		.chanx_left_in_94_(cbx_1__1__1_chanx_out_94_[0]),
		.chanx_left_in_96_(cbx_1__1__1_chanx_out_96_[0]),
		.chanx_left_in_98_(cbx_1__1__1_chanx_out_98_[0]),
		.chanx_left_in_100_(cbx_1__1__1_chanx_out_100_[0]),
		.chanx_left_in_102_(cbx_1__1__1_chanx_out_102_[0]),
		.chanx_left_in_104_(cbx_1__1__1_chanx_out_104_[0]),
		.chanx_left_in_106_(cbx_1__1__1_chanx_out_106_[0]),
		.chanx_left_in_108_(cbx_1__1__1_chanx_out_108_[0]),
		.chanx_left_in_110_(cbx_1__1__1_chanx_out_110_[0]),
		.chanx_left_in_112_(cbx_1__1__1_chanx_out_112_[0]),
		.chanx_left_in_114_(cbx_1__1__1_chanx_out_114_[0]),
		.chanx_left_in_116_(cbx_1__1__1_chanx_out_116_[0]),
		.chanx_left_in_118_(cbx_1__1__1_chanx_out_118_[0]),
		.chanx_left_in_120_(cbx_1__1__1_chanx_out_120_[0]),
		.chanx_left_in_122_(cbx_1__1__1_chanx_out_122_[0]),
		.chanx_left_in_124_(cbx_1__1__1_chanx_out_124_[0]),
		.chanx_left_in_126_(cbx_1__1__1_chanx_out_126_[0]),
		.chanx_left_in_128_(cbx_1__1__1_chanx_out_128_[0]),
		.chanx_left_in_130_(cbx_1__1__1_chanx_out_130_[0]),
		.chanx_left_in_132_(cbx_1__1__1_chanx_out_132_[0]),
		.chanx_left_in_134_(cbx_1__1__1_chanx_out_134_[0]),
		.chanx_left_in_136_(cbx_1__1__1_chanx_out_136_[0]),
		.chanx_left_in_138_(cbx_1__1__1_chanx_out_138_[0]),
		.chanx_left_in_140_(cbx_1__1__1_chanx_out_140_[0]),
		.chanx_left_in_142_(cbx_1__1__1_chanx_out_142_[0]),
		.chanx_left_in_144_(cbx_1__1__1_chanx_out_144_[0]),
		.chanx_left_in_146_(cbx_1__1__1_chanx_out_146_[0]),
		.chanx_left_in_148_(cbx_1__1__1_chanx_out_148_[0]),
		.chanx_left_in_150_(cbx_1__1__1_chanx_out_150_[0]),
		.chanx_left_in_152_(cbx_1__1__1_chanx_out_152_[0]),
		.chanx_left_in_154_(cbx_1__1__1_chanx_out_154_[0]),
		.chanx_left_in_156_(cbx_1__1__1_chanx_out_156_[0]),
		.chanx_left_in_158_(cbx_1__1__1_chanx_out_158_[0]),
		.chanx_left_in_160_(cbx_1__1__1_chanx_out_160_[0]),
		.chanx_left_in_162_(cbx_1__1__1_chanx_out_162_[0]),
		.chanx_left_in_164_(cbx_1__1__1_chanx_out_164_[0]),
		.chanx_left_in_166_(cbx_1__1__1_chanx_out_166_[0]),
		.chanx_left_in_168_(cbx_1__1__1_chanx_out_168_[0]),
		.chanx_left_in_170_(cbx_1__1__1_chanx_out_170_[0]),
		.chanx_left_in_172_(cbx_1__1__1_chanx_out_172_[0]),
		.chanx_left_in_174_(cbx_1__1__1_chanx_out_174_[0]),
		.chanx_left_in_176_(cbx_1__1__1_chanx_out_176_[0]),
		.chanx_left_in_178_(cbx_1__1__1_chanx_out_178_[0]),
		.chanx_left_in_180_(cbx_1__1__1_chanx_out_180_[0]),
		.chanx_left_in_182_(cbx_1__1__1_chanx_out_182_[0]),
		.chanx_left_in_184_(cbx_1__1__1_chanx_out_184_[0]),
		.chanx_left_in_186_(cbx_1__1__1_chanx_out_186_[0]),
		.chanx_left_in_188_(cbx_1__1__1_chanx_out_188_[0]),
		.chanx_left_in_190_(cbx_1__1__1_chanx_out_190_[0]),
		.chanx_left_in_192_(cbx_1__1__1_chanx_out_192_[0]),
		.chanx_left_in_194_(cbx_1__1__1_chanx_out_194_[0]),
		.chanx_left_in_196_(cbx_1__1__1_chanx_out_196_[0]),
		.chanx_left_in_198_(cbx_1__1__1_chanx_out_198_[0]),
		.left_top_grid_pin_54_(grid_clb_2_bottom_width_0_height_0__pin_54_lower[0]),
		.left_top_grid_pin_55_(grid_clb_2_bottom_width_0_height_0__pin_55_lower[0]),
		.left_top_grid_pin_56_(grid_clb_2_bottom_width_0_height_0__pin_56_lower[0]),
		.left_top_grid_pin_57_(grid_clb_2_bottom_width_0_height_0__pin_57_lower[0]),
		.left_top_grid_pin_58_(grid_clb_2_bottom_width_0_height_0__pin_58_lower[0]),
		.left_top_grid_pin_59_(grid_clb_2_bottom_width_0_height_0__pin_59_lower[0]),
		.left_top_grid_pin_60_(grid_clb_2_bottom_width_0_height_0__pin_60_lower[0]),
		.left_top_grid_pin_61_(grid_clb_2_bottom_width_0_height_0__pin_61_lower[0]),
		.left_top_grid_pin_62_(grid_clb_2_bottom_width_0_height_0__pin_62_lower[0]),
		.left_top_grid_pin_63_(grid_clb_2_bottom_width_0_height_0__pin_63_lower[0]),
		.left_top_grid_pin_66_(grid_clb_2_bottom_width_0_height_0__pin_66_lower[0]),
		.left_top_grid_pin_67_(grid_clb_2_bottom_width_0_height_0__pin_67_lower[0]),
		.ccff_head(grid_clb_1_ccff_tail[0]),
		.chany_top_out_0_(sb_2__1__0_chany_top_out_0_[0]),
		.chany_top_out_2_(sb_2__1__0_chany_top_out_2_[0]),
		.chany_top_out_4_(sb_2__1__0_chany_top_out_4_[0]),
		.chany_top_out_6_(sb_2__1__0_chany_top_out_6_[0]),
		.chany_top_out_8_(sb_2__1__0_chany_top_out_8_[0]),
		.chany_top_out_10_(sb_2__1__0_chany_top_out_10_[0]),
		.chany_top_out_12_(sb_2__1__0_chany_top_out_12_[0]),
		.chany_top_out_14_(sb_2__1__0_chany_top_out_14_[0]),
		.chany_top_out_16_(sb_2__1__0_chany_top_out_16_[0]),
		.chany_top_out_18_(sb_2__1__0_chany_top_out_18_[0]),
		.chany_top_out_20_(sb_2__1__0_chany_top_out_20_[0]),
		.chany_top_out_22_(sb_2__1__0_chany_top_out_22_[0]),
		.chany_top_out_24_(sb_2__1__0_chany_top_out_24_[0]),
		.chany_top_out_26_(sb_2__1__0_chany_top_out_26_[0]),
		.chany_top_out_28_(sb_2__1__0_chany_top_out_28_[0]),
		.chany_top_out_30_(sb_2__1__0_chany_top_out_30_[0]),
		.chany_top_out_32_(sb_2__1__0_chany_top_out_32_[0]),
		.chany_top_out_34_(sb_2__1__0_chany_top_out_34_[0]),
		.chany_top_out_36_(sb_2__1__0_chany_top_out_36_[0]),
		.chany_top_out_38_(sb_2__1__0_chany_top_out_38_[0]),
		.chany_top_out_40_(sb_2__1__0_chany_top_out_40_[0]),
		.chany_top_out_42_(sb_2__1__0_chany_top_out_42_[0]),
		.chany_top_out_44_(sb_2__1__0_chany_top_out_44_[0]),
		.chany_top_out_46_(sb_2__1__0_chany_top_out_46_[0]),
		.chany_top_out_48_(sb_2__1__0_chany_top_out_48_[0]),
		.chany_top_out_50_(sb_2__1__0_chany_top_out_50_[0]),
		.chany_top_out_52_(sb_2__1__0_chany_top_out_52_[0]),
		.chany_top_out_54_(sb_2__1__0_chany_top_out_54_[0]),
		.chany_top_out_56_(sb_2__1__0_chany_top_out_56_[0]),
		.chany_top_out_58_(sb_2__1__0_chany_top_out_58_[0]),
		.chany_top_out_60_(sb_2__1__0_chany_top_out_60_[0]),
		.chany_top_out_62_(sb_2__1__0_chany_top_out_62_[0]),
		.chany_top_out_64_(sb_2__1__0_chany_top_out_64_[0]),
		.chany_top_out_66_(sb_2__1__0_chany_top_out_66_[0]),
		.chany_top_out_68_(sb_2__1__0_chany_top_out_68_[0]),
		.chany_top_out_70_(sb_2__1__0_chany_top_out_70_[0]),
		.chany_top_out_72_(sb_2__1__0_chany_top_out_72_[0]),
		.chany_top_out_74_(sb_2__1__0_chany_top_out_74_[0]),
		.chany_top_out_76_(sb_2__1__0_chany_top_out_76_[0]),
		.chany_top_out_78_(sb_2__1__0_chany_top_out_78_[0]),
		.chany_top_out_80_(sb_2__1__0_chany_top_out_80_[0]),
		.chany_top_out_82_(sb_2__1__0_chany_top_out_82_[0]),
		.chany_top_out_84_(sb_2__1__0_chany_top_out_84_[0]),
		.chany_top_out_86_(sb_2__1__0_chany_top_out_86_[0]),
		.chany_top_out_88_(sb_2__1__0_chany_top_out_88_[0]),
		.chany_top_out_90_(sb_2__1__0_chany_top_out_90_[0]),
		.chany_top_out_92_(sb_2__1__0_chany_top_out_92_[0]),
		.chany_top_out_94_(sb_2__1__0_chany_top_out_94_[0]),
		.chany_top_out_96_(sb_2__1__0_chany_top_out_96_[0]),
		.chany_top_out_98_(sb_2__1__0_chany_top_out_98_[0]),
		.chany_top_out_100_(sb_2__1__0_chany_top_out_100_[0]),
		.chany_top_out_102_(sb_2__1__0_chany_top_out_102_[0]),
		.chany_top_out_104_(sb_2__1__0_chany_top_out_104_[0]),
		.chany_top_out_106_(sb_2__1__0_chany_top_out_106_[0]),
		.chany_top_out_108_(sb_2__1__0_chany_top_out_108_[0]),
		.chany_top_out_110_(sb_2__1__0_chany_top_out_110_[0]),
		.chany_top_out_112_(sb_2__1__0_chany_top_out_112_[0]),
		.chany_top_out_114_(sb_2__1__0_chany_top_out_114_[0]),
		.chany_top_out_116_(sb_2__1__0_chany_top_out_116_[0]),
		.chany_top_out_118_(sb_2__1__0_chany_top_out_118_[0]),
		.chany_top_out_120_(sb_2__1__0_chany_top_out_120_[0]),
		.chany_top_out_122_(sb_2__1__0_chany_top_out_122_[0]),
		.chany_top_out_124_(sb_2__1__0_chany_top_out_124_[0]),
		.chany_top_out_126_(sb_2__1__0_chany_top_out_126_[0]),
		.chany_top_out_128_(sb_2__1__0_chany_top_out_128_[0]),
		.chany_top_out_130_(sb_2__1__0_chany_top_out_130_[0]),
		.chany_top_out_132_(sb_2__1__0_chany_top_out_132_[0]),
		.chany_top_out_134_(sb_2__1__0_chany_top_out_134_[0]),
		.chany_top_out_136_(sb_2__1__0_chany_top_out_136_[0]),
		.chany_top_out_138_(sb_2__1__0_chany_top_out_138_[0]),
		.chany_top_out_140_(sb_2__1__0_chany_top_out_140_[0]),
		.chany_top_out_142_(sb_2__1__0_chany_top_out_142_[0]),
		.chany_top_out_144_(sb_2__1__0_chany_top_out_144_[0]),
		.chany_top_out_146_(sb_2__1__0_chany_top_out_146_[0]),
		.chany_top_out_148_(sb_2__1__0_chany_top_out_148_[0]),
		.chany_top_out_150_(sb_2__1__0_chany_top_out_150_[0]),
		.chany_top_out_152_(sb_2__1__0_chany_top_out_152_[0]),
		.chany_top_out_154_(sb_2__1__0_chany_top_out_154_[0]),
		.chany_top_out_156_(sb_2__1__0_chany_top_out_156_[0]),
		.chany_top_out_158_(sb_2__1__0_chany_top_out_158_[0]),
		.chany_top_out_160_(sb_2__1__0_chany_top_out_160_[0]),
		.chany_top_out_162_(sb_2__1__0_chany_top_out_162_[0]),
		.chany_top_out_164_(sb_2__1__0_chany_top_out_164_[0]),
		.chany_top_out_166_(sb_2__1__0_chany_top_out_166_[0]),
		.chany_top_out_168_(sb_2__1__0_chany_top_out_168_[0]),
		.chany_top_out_170_(sb_2__1__0_chany_top_out_170_[0]),
		.chany_top_out_172_(sb_2__1__0_chany_top_out_172_[0]),
		.chany_top_out_174_(sb_2__1__0_chany_top_out_174_[0]),
		.chany_top_out_176_(sb_2__1__0_chany_top_out_176_[0]),
		.chany_top_out_178_(sb_2__1__0_chany_top_out_178_[0]),
		.chany_top_out_180_(sb_2__1__0_chany_top_out_180_[0]),
		.chany_top_out_182_(sb_2__1__0_chany_top_out_182_[0]),
		.chany_top_out_184_(sb_2__1__0_chany_top_out_184_[0]),
		.chany_top_out_186_(sb_2__1__0_chany_top_out_186_[0]),
		.chany_top_out_188_(sb_2__1__0_chany_top_out_188_[0]),
		.chany_top_out_190_(sb_2__1__0_chany_top_out_190_[0]),
		.chany_top_out_192_(sb_2__1__0_chany_top_out_192_[0]),
		.chany_top_out_194_(sb_2__1__0_chany_top_out_194_[0]),
		.chany_top_out_196_(sb_2__1__0_chany_top_out_196_[0]),
		.chany_top_out_198_(sb_2__1__0_chany_top_out_198_[0]),
		.chany_bottom_out_1_(sb_2__1__0_chany_bottom_out_1_[0]),
		.chany_bottom_out_3_(sb_2__1__0_chany_bottom_out_3_[0]),
		.chany_bottom_out_5_(sb_2__1__0_chany_bottom_out_5_[0]),
		.chany_bottom_out_7_(sb_2__1__0_chany_bottom_out_7_[0]),
		.chany_bottom_out_9_(sb_2__1__0_chany_bottom_out_9_[0]),
		.chany_bottom_out_11_(sb_2__1__0_chany_bottom_out_11_[0]),
		.chany_bottom_out_13_(sb_2__1__0_chany_bottom_out_13_[0]),
		.chany_bottom_out_15_(sb_2__1__0_chany_bottom_out_15_[0]),
		.chany_bottom_out_17_(sb_2__1__0_chany_bottom_out_17_[0]),
		.chany_bottom_out_19_(sb_2__1__0_chany_bottom_out_19_[0]),
		.chany_bottom_out_21_(sb_2__1__0_chany_bottom_out_21_[0]),
		.chany_bottom_out_23_(sb_2__1__0_chany_bottom_out_23_[0]),
		.chany_bottom_out_25_(sb_2__1__0_chany_bottom_out_25_[0]),
		.chany_bottom_out_27_(sb_2__1__0_chany_bottom_out_27_[0]),
		.chany_bottom_out_29_(sb_2__1__0_chany_bottom_out_29_[0]),
		.chany_bottom_out_31_(sb_2__1__0_chany_bottom_out_31_[0]),
		.chany_bottom_out_33_(sb_2__1__0_chany_bottom_out_33_[0]),
		.chany_bottom_out_35_(sb_2__1__0_chany_bottom_out_35_[0]),
		.chany_bottom_out_37_(sb_2__1__0_chany_bottom_out_37_[0]),
		.chany_bottom_out_39_(sb_2__1__0_chany_bottom_out_39_[0]),
		.chany_bottom_out_41_(sb_2__1__0_chany_bottom_out_41_[0]),
		.chany_bottom_out_43_(sb_2__1__0_chany_bottom_out_43_[0]),
		.chany_bottom_out_45_(sb_2__1__0_chany_bottom_out_45_[0]),
		.chany_bottom_out_47_(sb_2__1__0_chany_bottom_out_47_[0]),
		.chany_bottom_out_49_(sb_2__1__0_chany_bottom_out_49_[0]),
		.chany_bottom_out_51_(sb_2__1__0_chany_bottom_out_51_[0]),
		.chany_bottom_out_53_(sb_2__1__0_chany_bottom_out_53_[0]),
		.chany_bottom_out_55_(sb_2__1__0_chany_bottom_out_55_[0]),
		.chany_bottom_out_57_(sb_2__1__0_chany_bottom_out_57_[0]),
		.chany_bottom_out_59_(sb_2__1__0_chany_bottom_out_59_[0]),
		.chany_bottom_out_61_(sb_2__1__0_chany_bottom_out_61_[0]),
		.chany_bottom_out_63_(sb_2__1__0_chany_bottom_out_63_[0]),
		.chany_bottom_out_65_(sb_2__1__0_chany_bottom_out_65_[0]),
		.chany_bottom_out_67_(sb_2__1__0_chany_bottom_out_67_[0]),
		.chany_bottom_out_69_(sb_2__1__0_chany_bottom_out_69_[0]),
		.chany_bottom_out_71_(sb_2__1__0_chany_bottom_out_71_[0]),
		.chany_bottom_out_73_(sb_2__1__0_chany_bottom_out_73_[0]),
		.chany_bottom_out_75_(sb_2__1__0_chany_bottom_out_75_[0]),
		.chany_bottom_out_77_(sb_2__1__0_chany_bottom_out_77_[0]),
		.chany_bottom_out_79_(sb_2__1__0_chany_bottom_out_79_[0]),
		.chany_bottom_out_81_(sb_2__1__0_chany_bottom_out_81_[0]),
		.chany_bottom_out_83_(sb_2__1__0_chany_bottom_out_83_[0]),
		.chany_bottom_out_85_(sb_2__1__0_chany_bottom_out_85_[0]),
		.chany_bottom_out_87_(sb_2__1__0_chany_bottom_out_87_[0]),
		.chany_bottom_out_89_(sb_2__1__0_chany_bottom_out_89_[0]),
		.chany_bottom_out_91_(sb_2__1__0_chany_bottom_out_91_[0]),
		.chany_bottom_out_93_(sb_2__1__0_chany_bottom_out_93_[0]),
		.chany_bottom_out_95_(sb_2__1__0_chany_bottom_out_95_[0]),
		.chany_bottom_out_97_(sb_2__1__0_chany_bottom_out_97_[0]),
		.chany_bottom_out_99_(sb_2__1__0_chany_bottom_out_99_[0]),
		.chany_bottom_out_101_(sb_2__1__0_chany_bottom_out_101_[0]),
		.chany_bottom_out_103_(sb_2__1__0_chany_bottom_out_103_[0]),
		.chany_bottom_out_105_(sb_2__1__0_chany_bottom_out_105_[0]),
		.chany_bottom_out_107_(sb_2__1__0_chany_bottom_out_107_[0]),
		.chany_bottom_out_109_(sb_2__1__0_chany_bottom_out_109_[0]),
		.chany_bottom_out_111_(sb_2__1__0_chany_bottom_out_111_[0]),
		.chany_bottom_out_113_(sb_2__1__0_chany_bottom_out_113_[0]),
		.chany_bottom_out_115_(sb_2__1__0_chany_bottom_out_115_[0]),
		.chany_bottom_out_117_(sb_2__1__0_chany_bottom_out_117_[0]),
		.chany_bottom_out_119_(sb_2__1__0_chany_bottom_out_119_[0]),
		.chany_bottom_out_121_(sb_2__1__0_chany_bottom_out_121_[0]),
		.chany_bottom_out_123_(sb_2__1__0_chany_bottom_out_123_[0]),
		.chany_bottom_out_125_(sb_2__1__0_chany_bottom_out_125_[0]),
		.chany_bottom_out_127_(sb_2__1__0_chany_bottom_out_127_[0]),
		.chany_bottom_out_129_(sb_2__1__0_chany_bottom_out_129_[0]),
		.chany_bottom_out_131_(sb_2__1__0_chany_bottom_out_131_[0]),
		.chany_bottom_out_133_(sb_2__1__0_chany_bottom_out_133_[0]),
		.chany_bottom_out_135_(sb_2__1__0_chany_bottom_out_135_[0]),
		.chany_bottom_out_137_(sb_2__1__0_chany_bottom_out_137_[0]),
		.chany_bottom_out_139_(sb_2__1__0_chany_bottom_out_139_[0]),
		.chany_bottom_out_141_(sb_2__1__0_chany_bottom_out_141_[0]),
		.chany_bottom_out_143_(sb_2__1__0_chany_bottom_out_143_[0]),
		.chany_bottom_out_145_(sb_2__1__0_chany_bottom_out_145_[0]),
		.chany_bottom_out_147_(sb_2__1__0_chany_bottom_out_147_[0]),
		.chany_bottom_out_149_(sb_2__1__0_chany_bottom_out_149_[0]),
		.chany_bottom_out_151_(sb_2__1__0_chany_bottom_out_151_[0]),
		.chany_bottom_out_153_(sb_2__1__0_chany_bottom_out_153_[0]),
		.chany_bottom_out_155_(sb_2__1__0_chany_bottom_out_155_[0]),
		.chany_bottom_out_157_(sb_2__1__0_chany_bottom_out_157_[0]),
		.chany_bottom_out_159_(sb_2__1__0_chany_bottom_out_159_[0]),
		.chany_bottom_out_161_(sb_2__1__0_chany_bottom_out_161_[0]),
		.chany_bottom_out_163_(sb_2__1__0_chany_bottom_out_163_[0]),
		.chany_bottom_out_165_(sb_2__1__0_chany_bottom_out_165_[0]),
		.chany_bottom_out_167_(sb_2__1__0_chany_bottom_out_167_[0]),
		.chany_bottom_out_169_(sb_2__1__0_chany_bottom_out_169_[0]),
		.chany_bottom_out_171_(sb_2__1__0_chany_bottom_out_171_[0]),
		.chany_bottom_out_173_(sb_2__1__0_chany_bottom_out_173_[0]),
		.chany_bottom_out_175_(sb_2__1__0_chany_bottom_out_175_[0]),
		.chany_bottom_out_177_(sb_2__1__0_chany_bottom_out_177_[0]),
		.chany_bottom_out_179_(sb_2__1__0_chany_bottom_out_179_[0]),
		.chany_bottom_out_181_(sb_2__1__0_chany_bottom_out_181_[0]),
		.chany_bottom_out_183_(sb_2__1__0_chany_bottom_out_183_[0]),
		.chany_bottom_out_185_(sb_2__1__0_chany_bottom_out_185_[0]),
		.chany_bottom_out_187_(sb_2__1__0_chany_bottom_out_187_[0]),
		.chany_bottom_out_189_(sb_2__1__0_chany_bottom_out_189_[0]),
		.chany_bottom_out_191_(sb_2__1__0_chany_bottom_out_191_[0]),
		.chany_bottom_out_193_(sb_2__1__0_chany_bottom_out_193_[0]),
		.chany_bottom_out_195_(sb_2__1__0_chany_bottom_out_195_[0]),
		.chany_bottom_out_197_(sb_2__1__0_chany_bottom_out_197_[0]),
		.chany_bottom_out_199_(sb_2__1__0_chany_bottom_out_199_[0]),
		.chanx_left_out_1_(sb_2__1__0_chanx_left_out_1_[0]),
		.chanx_left_out_3_(sb_2__1__0_chanx_left_out_3_[0]),
		.chanx_left_out_5_(sb_2__1__0_chanx_left_out_5_[0]),
		.chanx_left_out_7_(sb_2__1__0_chanx_left_out_7_[0]),
		.chanx_left_out_9_(sb_2__1__0_chanx_left_out_9_[0]),
		.chanx_left_out_11_(sb_2__1__0_chanx_left_out_11_[0]),
		.chanx_left_out_13_(sb_2__1__0_chanx_left_out_13_[0]),
		.chanx_left_out_15_(sb_2__1__0_chanx_left_out_15_[0]),
		.chanx_left_out_17_(sb_2__1__0_chanx_left_out_17_[0]),
		.chanx_left_out_19_(sb_2__1__0_chanx_left_out_19_[0]),
		.chanx_left_out_21_(sb_2__1__0_chanx_left_out_21_[0]),
		.chanx_left_out_23_(sb_2__1__0_chanx_left_out_23_[0]),
		.chanx_left_out_25_(sb_2__1__0_chanx_left_out_25_[0]),
		.chanx_left_out_27_(sb_2__1__0_chanx_left_out_27_[0]),
		.chanx_left_out_29_(sb_2__1__0_chanx_left_out_29_[0]),
		.chanx_left_out_31_(sb_2__1__0_chanx_left_out_31_[0]),
		.chanx_left_out_33_(sb_2__1__0_chanx_left_out_33_[0]),
		.chanx_left_out_35_(sb_2__1__0_chanx_left_out_35_[0]),
		.chanx_left_out_37_(sb_2__1__0_chanx_left_out_37_[0]),
		.chanx_left_out_39_(sb_2__1__0_chanx_left_out_39_[0]),
		.chanx_left_out_41_(sb_2__1__0_chanx_left_out_41_[0]),
		.chanx_left_out_43_(sb_2__1__0_chanx_left_out_43_[0]),
		.chanx_left_out_45_(sb_2__1__0_chanx_left_out_45_[0]),
		.chanx_left_out_47_(sb_2__1__0_chanx_left_out_47_[0]),
		.chanx_left_out_49_(sb_2__1__0_chanx_left_out_49_[0]),
		.chanx_left_out_51_(sb_2__1__0_chanx_left_out_51_[0]),
		.chanx_left_out_53_(sb_2__1__0_chanx_left_out_53_[0]),
		.chanx_left_out_55_(sb_2__1__0_chanx_left_out_55_[0]),
		.chanx_left_out_57_(sb_2__1__0_chanx_left_out_57_[0]),
		.chanx_left_out_59_(sb_2__1__0_chanx_left_out_59_[0]),
		.chanx_left_out_61_(sb_2__1__0_chanx_left_out_61_[0]),
		.chanx_left_out_63_(sb_2__1__0_chanx_left_out_63_[0]),
		.chanx_left_out_65_(sb_2__1__0_chanx_left_out_65_[0]),
		.chanx_left_out_67_(sb_2__1__0_chanx_left_out_67_[0]),
		.chanx_left_out_69_(sb_2__1__0_chanx_left_out_69_[0]),
		.chanx_left_out_71_(sb_2__1__0_chanx_left_out_71_[0]),
		.chanx_left_out_73_(sb_2__1__0_chanx_left_out_73_[0]),
		.chanx_left_out_75_(sb_2__1__0_chanx_left_out_75_[0]),
		.chanx_left_out_77_(sb_2__1__0_chanx_left_out_77_[0]),
		.chanx_left_out_79_(sb_2__1__0_chanx_left_out_79_[0]),
		.chanx_left_out_81_(sb_2__1__0_chanx_left_out_81_[0]),
		.chanx_left_out_83_(sb_2__1__0_chanx_left_out_83_[0]),
		.chanx_left_out_85_(sb_2__1__0_chanx_left_out_85_[0]),
		.chanx_left_out_87_(sb_2__1__0_chanx_left_out_87_[0]),
		.chanx_left_out_89_(sb_2__1__0_chanx_left_out_89_[0]),
		.chanx_left_out_91_(sb_2__1__0_chanx_left_out_91_[0]),
		.chanx_left_out_93_(sb_2__1__0_chanx_left_out_93_[0]),
		.chanx_left_out_95_(sb_2__1__0_chanx_left_out_95_[0]),
		.chanx_left_out_97_(sb_2__1__0_chanx_left_out_97_[0]),
		.chanx_left_out_99_(sb_2__1__0_chanx_left_out_99_[0]),
		.chanx_left_out_101_(sb_2__1__0_chanx_left_out_101_[0]),
		.chanx_left_out_103_(sb_2__1__0_chanx_left_out_103_[0]),
		.chanx_left_out_105_(sb_2__1__0_chanx_left_out_105_[0]),
		.chanx_left_out_107_(sb_2__1__0_chanx_left_out_107_[0]),
		.chanx_left_out_109_(sb_2__1__0_chanx_left_out_109_[0]),
		.chanx_left_out_111_(sb_2__1__0_chanx_left_out_111_[0]),
		.chanx_left_out_113_(sb_2__1__0_chanx_left_out_113_[0]),
		.chanx_left_out_115_(sb_2__1__0_chanx_left_out_115_[0]),
		.chanx_left_out_117_(sb_2__1__0_chanx_left_out_117_[0]),
		.chanx_left_out_119_(sb_2__1__0_chanx_left_out_119_[0]),
		.chanx_left_out_121_(sb_2__1__0_chanx_left_out_121_[0]),
		.chanx_left_out_123_(sb_2__1__0_chanx_left_out_123_[0]),
		.chanx_left_out_125_(sb_2__1__0_chanx_left_out_125_[0]),
		.chanx_left_out_127_(sb_2__1__0_chanx_left_out_127_[0]),
		.chanx_left_out_129_(sb_2__1__0_chanx_left_out_129_[0]),
		.chanx_left_out_131_(sb_2__1__0_chanx_left_out_131_[0]),
		.chanx_left_out_133_(sb_2__1__0_chanx_left_out_133_[0]),
		.chanx_left_out_135_(sb_2__1__0_chanx_left_out_135_[0]),
		.chanx_left_out_137_(sb_2__1__0_chanx_left_out_137_[0]),
		.chanx_left_out_139_(sb_2__1__0_chanx_left_out_139_[0]),
		.chanx_left_out_141_(sb_2__1__0_chanx_left_out_141_[0]),
		.chanx_left_out_143_(sb_2__1__0_chanx_left_out_143_[0]),
		.chanx_left_out_145_(sb_2__1__0_chanx_left_out_145_[0]),
		.chanx_left_out_147_(sb_2__1__0_chanx_left_out_147_[0]),
		.chanx_left_out_149_(sb_2__1__0_chanx_left_out_149_[0]),
		.chanx_left_out_151_(sb_2__1__0_chanx_left_out_151_[0]),
		.chanx_left_out_153_(sb_2__1__0_chanx_left_out_153_[0]),
		.chanx_left_out_155_(sb_2__1__0_chanx_left_out_155_[0]),
		.chanx_left_out_157_(sb_2__1__0_chanx_left_out_157_[0]),
		.chanx_left_out_159_(sb_2__1__0_chanx_left_out_159_[0]),
		.chanx_left_out_161_(sb_2__1__0_chanx_left_out_161_[0]),
		.chanx_left_out_163_(sb_2__1__0_chanx_left_out_163_[0]),
		.chanx_left_out_165_(sb_2__1__0_chanx_left_out_165_[0]),
		.chanx_left_out_167_(sb_2__1__0_chanx_left_out_167_[0]),
		.chanx_left_out_169_(sb_2__1__0_chanx_left_out_169_[0]),
		.chanx_left_out_171_(sb_2__1__0_chanx_left_out_171_[0]),
		.chanx_left_out_173_(sb_2__1__0_chanx_left_out_173_[0]),
		.chanx_left_out_175_(sb_2__1__0_chanx_left_out_175_[0]),
		.chanx_left_out_177_(sb_2__1__0_chanx_left_out_177_[0]),
		.chanx_left_out_179_(sb_2__1__0_chanx_left_out_179_[0]),
		.chanx_left_out_181_(sb_2__1__0_chanx_left_out_181_[0]),
		.chanx_left_out_183_(sb_2__1__0_chanx_left_out_183_[0]),
		.chanx_left_out_185_(sb_2__1__0_chanx_left_out_185_[0]),
		.chanx_left_out_187_(sb_2__1__0_chanx_left_out_187_[0]),
		.chanx_left_out_189_(sb_2__1__0_chanx_left_out_189_[0]),
		.chanx_left_out_191_(sb_2__1__0_chanx_left_out_191_[0]),
		.chanx_left_out_193_(sb_2__1__0_chanx_left_out_193_[0]),
		.chanx_left_out_195_(sb_2__1__0_chanx_left_out_195_[0]),
		.chanx_left_out_197_(sb_2__1__0_chanx_left_out_197_[0]),
		.chanx_left_out_199_(sb_2__1__0_chanx_left_out_199_[0]),
		.ccff_tail(sb_2__1__0_ccff_tail[0]));

	sb_2__2_ sb_2__2_ (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.chany_bottom_in_0_(cby_2__1__1_chany_out_0_[0]),
		.chany_bottom_in_2_(cby_2__1__1_chany_out_2_[0]),
		.chany_bottom_in_4_(cby_2__1__1_chany_out_4_[0]),
		.chany_bottom_in_6_(cby_2__1__1_chany_out_6_[0]),
		.chany_bottom_in_8_(cby_2__1__1_chany_out_8_[0]),
		.chany_bottom_in_10_(cby_2__1__1_chany_out_10_[0]),
		.chany_bottom_in_12_(cby_2__1__1_chany_out_12_[0]),
		.chany_bottom_in_14_(cby_2__1__1_chany_out_14_[0]),
		.chany_bottom_in_16_(cby_2__1__1_chany_out_16_[0]),
		.chany_bottom_in_18_(cby_2__1__1_chany_out_18_[0]),
		.chany_bottom_in_20_(cby_2__1__1_chany_out_20_[0]),
		.chany_bottom_in_22_(cby_2__1__1_chany_out_22_[0]),
		.chany_bottom_in_24_(cby_2__1__1_chany_out_24_[0]),
		.chany_bottom_in_26_(cby_2__1__1_chany_out_26_[0]),
		.chany_bottom_in_28_(cby_2__1__1_chany_out_28_[0]),
		.chany_bottom_in_30_(cby_2__1__1_chany_out_30_[0]),
		.chany_bottom_in_32_(cby_2__1__1_chany_out_32_[0]),
		.chany_bottom_in_34_(cby_2__1__1_chany_out_34_[0]),
		.chany_bottom_in_36_(cby_2__1__1_chany_out_36_[0]),
		.chany_bottom_in_38_(cby_2__1__1_chany_out_38_[0]),
		.chany_bottom_in_40_(cby_2__1__1_chany_out_40_[0]),
		.chany_bottom_in_42_(cby_2__1__1_chany_out_42_[0]),
		.chany_bottom_in_44_(cby_2__1__1_chany_out_44_[0]),
		.chany_bottom_in_46_(cby_2__1__1_chany_out_46_[0]),
		.chany_bottom_in_48_(cby_2__1__1_chany_out_48_[0]),
		.chany_bottom_in_50_(cby_2__1__1_chany_out_50_[0]),
		.chany_bottom_in_52_(cby_2__1__1_chany_out_52_[0]),
		.chany_bottom_in_54_(cby_2__1__1_chany_out_54_[0]),
		.chany_bottom_in_56_(cby_2__1__1_chany_out_56_[0]),
		.chany_bottom_in_58_(cby_2__1__1_chany_out_58_[0]),
		.chany_bottom_in_60_(cby_2__1__1_chany_out_60_[0]),
		.chany_bottom_in_62_(cby_2__1__1_chany_out_62_[0]),
		.chany_bottom_in_64_(cby_2__1__1_chany_out_64_[0]),
		.chany_bottom_in_66_(cby_2__1__1_chany_out_66_[0]),
		.chany_bottom_in_68_(cby_2__1__1_chany_out_68_[0]),
		.chany_bottom_in_70_(cby_2__1__1_chany_out_70_[0]),
		.chany_bottom_in_72_(cby_2__1__1_chany_out_72_[0]),
		.chany_bottom_in_74_(cby_2__1__1_chany_out_74_[0]),
		.chany_bottom_in_76_(cby_2__1__1_chany_out_76_[0]),
		.chany_bottom_in_78_(cby_2__1__1_chany_out_78_[0]),
		.chany_bottom_in_80_(cby_2__1__1_chany_out_80_[0]),
		.chany_bottom_in_82_(cby_2__1__1_chany_out_82_[0]),
		.chany_bottom_in_84_(cby_2__1__1_chany_out_84_[0]),
		.chany_bottom_in_86_(cby_2__1__1_chany_out_86_[0]),
		.chany_bottom_in_88_(cby_2__1__1_chany_out_88_[0]),
		.chany_bottom_in_90_(cby_2__1__1_chany_out_90_[0]),
		.chany_bottom_in_92_(cby_2__1__1_chany_out_92_[0]),
		.chany_bottom_in_94_(cby_2__1__1_chany_out_94_[0]),
		.chany_bottom_in_96_(cby_2__1__1_chany_out_96_[0]),
		.chany_bottom_in_98_(cby_2__1__1_chany_out_98_[0]),
		.chany_bottom_in_100_(cby_2__1__1_chany_out_100_[0]),
		.chany_bottom_in_102_(cby_2__1__1_chany_out_102_[0]),
		.chany_bottom_in_104_(cby_2__1__1_chany_out_104_[0]),
		.chany_bottom_in_106_(cby_2__1__1_chany_out_106_[0]),
		.chany_bottom_in_108_(cby_2__1__1_chany_out_108_[0]),
		.chany_bottom_in_110_(cby_2__1__1_chany_out_110_[0]),
		.chany_bottom_in_112_(cby_2__1__1_chany_out_112_[0]),
		.chany_bottom_in_114_(cby_2__1__1_chany_out_114_[0]),
		.chany_bottom_in_116_(cby_2__1__1_chany_out_116_[0]),
		.chany_bottom_in_118_(cby_2__1__1_chany_out_118_[0]),
		.chany_bottom_in_120_(cby_2__1__1_chany_out_120_[0]),
		.chany_bottom_in_122_(cby_2__1__1_chany_out_122_[0]),
		.chany_bottom_in_124_(cby_2__1__1_chany_out_124_[0]),
		.chany_bottom_in_126_(cby_2__1__1_chany_out_126_[0]),
		.chany_bottom_in_128_(cby_2__1__1_chany_out_128_[0]),
		.chany_bottom_in_130_(cby_2__1__1_chany_out_130_[0]),
		.chany_bottom_in_132_(cby_2__1__1_chany_out_132_[0]),
		.chany_bottom_in_134_(cby_2__1__1_chany_out_134_[0]),
		.chany_bottom_in_136_(cby_2__1__1_chany_out_136_[0]),
		.chany_bottom_in_138_(cby_2__1__1_chany_out_138_[0]),
		.chany_bottom_in_140_(cby_2__1__1_chany_out_140_[0]),
		.chany_bottom_in_142_(cby_2__1__1_chany_out_142_[0]),
		.chany_bottom_in_144_(cby_2__1__1_chany_out_144_[0]),
		.chany_bottom_in_146_(cby_2__1__1_chany_out_146_[0]),
		.chany_bottom_in_148_(cby_2__1__1_chany_out_148_[0]),
		.chany_bottom_in_150_(cby_2__1__1_chany_out_150_[0]),
		.chany_bottom_in_152_(cby_2__1__1_chany_out_152_[0]),
		.chany_bottom_in_154_(cby_2__1__1_chany_out_154_[0]),
		.chany_bottom_in_156_(cby_2__1__1_chany_out_156_[0]),
		.chany_bottom_in_158_(cby_2__1__1_chany_out_158_[0]),
		.chany_bottom_in_160_(cby_2__1__1_chany_out_160_[0]),
		.chany_bottom_in_162_(cby_2__1__1_chany_out_162_[0]),
		.chany_bottom_in_164_(cby_2__1__1_chany_out_164_[0]),
		.chany_bottom_in_166_(cby_2__1__1_chany_out_166_[0]),
		.chany_bottom_in_168_(cby_2__1__1_chany_out_168_[0]),
		.chany_bottom_in_170_(cby_2__1__1_chany_out_170_[0]),
		.chany_bottom_in_172_(cby_2__1__1_chany_out_172_[0]),
		.chany_bottom_in_174_(cby_2__1__1_chany_out_174_[0]),
		.chany_bottom_in_176_(cby_2__1__1_chany_out_176_[0]),
		.chany_bottom_in_178_(cby_2__1__1_chany_out_178_[0]),
		.chany_bottom_in_180_(cby_2__1__1_chany_out_180_[0]),
		.chany_bottom_in_182_(cby_2__1__1_chany_out_182_[0]),
		.chany_bottom_in_184_(cby_2__1__1_chany_out_184_[0]),
		.chany_bottom_in_186_(cby_2__1__1_chany_out_186_[0]),
		.chany_bottom_in_188_(cby_2__1__1_chany_out_188_[0]),
		.chany_bottom_in_190_(cby_2__1__1_chany_out_190_[0]),
		.chany_bottom_in_192_(cby_2__1__1_chany_out_192_[0]),
		.chany_bottom_in_194_(cby_2__1__1_chany_out_194_[0]),
		.chany_bottom_in_196_(cby_2__1__1_chany_out_196_[0]),
		.chany_bottom_in_198_(cby_2__1__1_chany_out_198_[0]),
		.bottom_right_grid_pin_1_(grid_io_right_1_left_width_0_height_0__pin_1_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_2_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_2_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_2_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_2_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_2_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_2_right_width_0_height_0__pin_49_upper[0]),
		.bottom_left_grid_pin_50_(grid_clb_2_right_width_0_height_0__pin_50_upper[0]),
		.bottom_left_grid_pin_51_(grid_clb_2_right_width_0_height_0__pin_51_upper[0]),
		.bottom_left_grid_pin_52_(grid_clb_2_right_width_0_height_0__pin_52_upper[0]),
		.bottom_left_grid_pin_53_(grid_clb_2_right_width_0_height_0__pin_53_upper[0]),
		.chanx_left_in_0_(cbx_1__2__1_chanx_out_0_[0]),
		.chanx_left_in_2_(cbx_1__2__1_chanx_out_2_[0]),
		.chanx_left_in_4_(cbx_1__2__1_chanx_out_4_[0]),
		.chanx_left_in_6_(cbx_1__2__1_chanx_out_6_[0]),
		.chanx_left_in_8_(cbx_1__2__1_chanx_out_8_[0]),
		.chanx_left_in_10_(cbx_1__2__1_chanx_out_10_[0]),
		.chanx_left_in_12_(cbx_1__2__1_chanx_out_12_[0]),
		.chanx_left_in_14_(cbx_1__2__1_chanx_out_14_[0]),
		.chanx_left_in_16_(cbx_1__2__1_chanx_out_16_[0]),
		.chanx_left_in_18_(cbx_1__2__1_chanx_out_18_[0]),
		.chanx_left_in_20_(cbx_1__2__1_chanx_out_20_[0]),
		.chanx_left_in_22_(cbx_1__2__1_chanx_out_22_[0]),
		.chanx_left_in_24_(cbx_1__2__1_chanx_out_24_[0]),
		.chanx_left_in_26_(cbx_1__2__1_chanx_out_26_[0]),
		.chanx_left_in_28_(cbx_1__2__1_chanx_out_28_[0]),
		.chanx_left_in_30_(cbx_1__2__1_chanx_out_30_[0]),
		.chanx_left_in_32_(cbx_1__2__1_chanx_out_32_[0]),
		.chanx_left_in_34_(cbx_1__2__1_chanx_out_34_[0]),
		.chanx_left_in_36_(cbx_1__2__1_chanx_out_36_[0]),
		.chanx_left_in_38_(cbx_1__2__1_chanx_out_38_[0]),
		.chanx_left_in_40_(cbx_1__2__1_chanx_out_40_[0]),
		.chanx_left_in_42_(cbx_1__2__1_chanx_out_42_[0]),
		.chanx_left_in_44_(cbx_1__2__1_chanx_out_44_[0]),
		.chanx_left_in_46_(cbx_1__2__1_chanx_out_46_[0]),
		.chanx_left_in_48_(cbx_1__2__1_chanx_out_48_[0]),
		.chanx_left_in_50_(cbx_1__2__1_chanx_out_50_[0]),
		.chanx_left_in_52_(cbx_1__2__1_chanx_out_52_[0]),
		.chanx_left_in_54_(cbx_1__2__1_chanx_out_54_[0]),
		.chanx_left_in_56_(cbx_1__2__1_chanx_out_56_[0]),
		.chanx_left_in_58_(cbx_1__2__1_chanx_out_58_[0]),
		.chanx_left_in_60_(cbx_1__2__1_chanx_out_60_[0]),
		.chanx_left_in_62_(cbx_1__2__1_chanx_out_62_[0]),
		.chanx_left_in_64_(cbx_1__2__1_chanx_out_64_[0]),
		.chanx_left_in_66_(cbx_1__2__1_chanx_out_66_[0]),
		.chanx_left_in_68_(cbx_1__2__1_chanx_out_68_[0]),
		.chanx_left_in_70_(cbx_1__2__1_chanx_out_70_[0]),
		.chanx_left_in_72_(cbx_1__2__1_chanx_out_72_[0]),
		.chanx_left_in_74_(cbx_1__2__1_chanx_out_74_[0]),
		.chanx_left_in_76_(cbx_1__2__1_chanx_out_76_[0]),
		.chanx_left_in_78_(cbx_1__2__1_chanx_out_78_[0]),
		.chanx_left_in_80_(cbx_1__2__1_chanx_out_80_[0]),
		.chanx_left_in_82_(cbx_1__2__1_chanx_out_82_[0]),
		.chanx_left_in_84_(cbx_1__2__1_chanx_out_84_[0]),
		.chanx_left_in_86_(cbx_1__2__1_chanx_out_86_[0]),
		.chanx_left_in_88_(cbx_1__2__1_chanx_out_88_[0]),
		.chanx_left_in_90_(cbx_1__2__1_chanx_out_90_[0]),
		.chanx_left_in_92_(cbx_1__2__1_chanx_out_92_[0]),
		.chanx_left_in_94_(cbx_1__2__1_chanx_out_94_[0]),
		.chanx_left_in_96_(cbx_1__2__1_chanx_out_96_[0]),
		.chanx_left_in_98_(cbx_1__2__1_chanx_out_98_[0]),
		.chanx_left_in_100_(cbx_1__2__1_chanx_out_100_[0]),
		.chanx_left_in_102_(cbx_1__2__1_chanx_out_102_[0]),
		.chanx_left_in_104_(cbx_1__2__1_chanx_out_104_[0]),
		.chanx_left_in_106_(cbx_1__2__1_chanx_out_106_[0]),
		.chanx_left_in_108_(cbx_1__2__1_chanx_out_108_[0]),
		.chanx_left_in_110_(cbx_1__2__1_chanx_out_110_[0]),
		.chanx_left_in_112_(cbx_1__2__1_chanx_out_112_[0]),
		.chanx_left_in_114_(cbx_1__2__1_chanx_out_114_[0]),
		.chanx_left_in_116_(cbx_1__2__1_chanx_out_116_[0]),
		.chanx_left_in_118_(cbx_1__2__1_chanx_out_118_[0]),
		.chanx_left_in_120_(cbx_1__2__1_chanx_out_120_[0]),
		.chanx_left_in_122_(cbx_1__2__1_chanx_out_122_[0]),
		.chanx_left_in_124_(cbx_1__2__1_chanx_out_124_[0]),
		.chanx_left_in_126_(cbx_1__2__1_chanx_out_126_[0]),
		.chanx_left_in_128_(cbx_1__2__1_chanx_out_128_[0]),
		.chanx_left_in_130_(cbx_1__2__1_chanx_out_130_[0]),
		.chanx_left_in_132_(cbx_1__2__1_chanx_out_132_[0]),
		.chanx_left_in_134_(cbx_1__2__1_chanx_out_134_[0]),
		.chanx_left_in_136_(cbx_1__2__1_chanx_out_136_[0]),
		.chanx_left_in_138_(cbx_1__2__1_chanx_out_138_[0]),
		.chanx_left_in_140_(cbx_1__2__1_chanx_out_140_[0]),
		.chanx_left_in_142_(cbx_1__2__1_chanx_out_142_[0]),
		.chanx_left_in_144_(cbx_1__2__1_chanx_out_144_[0]),
		.chanx_left_in_146_(cbx_1__2__1_chanx_out_146_[0]),
		.chanx_left_in_148_(cbx_1__2__1_chanx_out_148_[0]),
		.chanx_left_in_150_(cbx_1__2__1_chanx_out_150_[0]),
		.chanx_left_in_152_(cbx_1__2__1_chanx_out_152_[0]),
		.chanx_left_in_154_(cbx_1__2__1_chanx_out_154_[0]),
		.chanx_left_in_156_(cbx_1__2__1_chanx_out_156_[0]),
		.chanx_left_in_158_(cbx_1__2__1_chanx_out_158_[0]),
		.chanx_left_in_160_(cbx_1__2__1_chanx_out_160_[0]),
		.chanx_left_in_162_(cbx_1__2__1_chanx_out_162_[0]),
		.chanx_left_in_164_(cbx_1__2__1_chanx_out_164_[0]),
		.chanx_left_in_166_(cbx_1__2__1_chanx_out_166_[0]),
		.chanx_left_in_168_(cbx_1__2__1_chanx_out_168_[0]),
		.chanx_left_in_170_(cbx_1__2__1_chanx_out_170_[0]),
		.chanx_left_in_172_(cbx_1__2__1_chanx_out_172_[0]),
		.chanx_left_in_174_(cbx_1__2__1_chanx_out_174_[0]),
		.chanx_left_in_176_(cbx_1__2__1_chanx_out_176_[0]),
		.chanx_left_in_178_(cbx_1__2__1_chanx_out_178_[0]),
		.chanx_left_in_180_(cbx_1__2__1_chanx_out_180_[0]),
		.chanx_left_in_182_(cbx_1__2__1_chanx_out_182_[0]),
		.chanx_left_in_184_(cbx_1__2__1_chanx_out_184_[0]),
		.chanx_left_in_186_(cbx_1__2__1_chanx_out_186_[0]),
		.chanx_left_in_188_(cbx_1__2__1_chanx_out_188_[0]),
		.chanx_left_in_190_(cbx_1__2__1_chanx_out_190_[0]),
		.chanx_left_in_192_(cbx_1__2__1_chanx_out_192_[0]),
		.chanx_left_in_194_(cbx_1__2__1_chanx_out_194_[0]),
		.chanx_left_in_196_(cbx_1__2__1_chanx_out_196_[0]),
		.chanx_left_in_198_(cbx_1__2__1_chanx_out_198_[0]),
		.left_top_grid_pin_1_(grid_io_top_1_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_io_right_1_ccff_tail[0]),
		.chany_bottom_out_1_(sb_2__2__0_chany_bottom_out_1_[0]),
		.chany_bottom_out_3_(sb_2__2__0_chany_bottom_out_3_[0]),
		.chany_bottom_out_5_(sb_2__2__0_chany_bottom_out_5_[0]),
		.chany_bottom_out_7_(sb_2__2__0_chany_bottom_out_7_[0]),
		.chany_bottom_out_9_(sb_2__2__0_chany_bottom_out_9_[0]),
		.chany_bottom_out_11_(sb_2__2__0_chany_bottom_out_11_[0]),
		.chany_bottom_out_13_(sb_2__2__0_chany_bottom_out_13_[0]),
		.chany_bottom_out_15_(sb_2__2__0_chany_bottom_out_15_[0]),
		.chany_bottom_out_17_(sb_2__2__0_chany_bottom_out_17_[0]),
		.chany_bottom_out_19_(sb_2__2__0_chany_bottom_out_19_[0]),
		.chany_bottom_out_21_(sb_2__2__0_chany_bottom_out_21_[0]),
		.chany_bottom_out_23_(sb_2__2__0_chany_bottom_out_23_[0]),
		.chany_bottom_out_25_(sb_2__2__0_chany_bottom_out_25_[0]),
		.chany_bottom_out_27_(sb_2__2__0_chany_bottom_out_27_[0]),
		.chany_bottom_out_29_(sb_2__2__0_chany_bottom_out_29_[0]),
		.chany_bottom_out_31_(sb_2__2__0_chany_bottom_out_31_[0]),
		.chany_bottom_out_33_(sb_2__2__0_chany_bottom_out_33_[0]),
		.chany_bottom_out_35_(sb_2__2__0_chany_bottom_out_35_[0]),
		.chany_bottom_out_37_(sb_2__2__0_chany_bottom_out_37_[0]),
		.chany_bottom_out_39_(sb_2__2__0_chany_bottom_out_39_[0]),
		.chany_bottom_out_41_(sb_2__2__0_chany_bottom_out_41_[0]),
		.chany_bottom_out_43_(sb_2__2__0_chany_bottom_out_43_[0]),
		.chany_bottom_out_45_(sb_2__2__0_chany_bottom_out_45_[0]),
		.chany_bottom_out_47_(sb_2__2__0_chany_bottom_out_47_[0]),
		.chany_bottom_out_49_(sb_2__2__0_chany_bottom_out_49_[0]),
		.chany_bottom_out_51_(sb_2__2__0_chany_bottom_out_51_[0]),
		.chany_bottom_out_53_(sb_2__2__0_chany_bottom_out_53_[0]),
		.chany_bottom_out_55_(sb_2__2__0_chany_bottom_out_55_[0]),
		.chany_bottom_out_57_(sb_2__2__0_chany_bottom_out_57_[0]),
		.chany_bottom_out_59_(sb_2__2__0_chany_bottom_out_59_[0]),
		.chany_bottom_out_61_(sb_2__2__0_chany_bottom_out_61_[0]),
		.chany_bottom_out_63_(sb_2__2__0_chany_bottom_out_63_[0]),
		.chany_bottom_out_65_(sb_2__2__0_chany_bottom_out_65_[0]),
		.chany_bottom_out_67_(sb_2__2__0_chany_bottom_out_67_[0]),
		.chany_bottom_out_69_(sb_2__2__0_chany_bottom_out_69_[0]),
		.chany_bottom_out_71_(sb_2__2__0_chany_bottom_out_71_[0]),
		.chany_bottom_out_73_(sb_2__2__0_chany_bottom_out_73_[0]),
		.chany_bottom_out_75_(sb_2__2__0_chany_bottom_out_75_[0]),
		.chany_bottom_out_77_(sb_2__2__0_chany_bottom_out_77_[0]),
		.chany_bottom_out_79_(sb_2__2__0_chany_bottom_out_79_[0]),
		.chany_bottom_out_81_(sb_2__2__0_chany_bottom_out_81_[0]),
		.chany_bottom_out_83_(sb_2__2__0_chany_bottom_out_83_[0]),
		.chany_bottom_out_85_(sb_2__2__0_chany_bottom_out_85_[0]),
		.chany_bottom_out_87_(sb_2__2__0_chany_bottom_out_87_[0]),
		.chany_bottom_out_89_(sb_2__2__0_chany_bottom_out_89_[0]),
		.chany_bottom_out_91_(sb_2__2__0_chany_bottom_out_91_[0]),
		.chany_bottom_out_93_(sb_2__2__0_chany_bottom_out_93_[0]),
		.chany_bottom_out_95_(sb_2__2__0_chany_bottom_out_95_[0]),
		.chany_bottom_out_97_(sb_2__2__0_chany_bottom_out_97_[0]),
		.chany_bottom_out_99_(sb_2__2__0_chany_bottom_out_99_[0]),
		.chany_bottom_out_101_(sb_2__2__0_chany_bottom_out_101_[0]),
		.chany_bottom_out_103_(sb_2__2__0_chany_bottom_out_103_[0]),
		.chany_bottom_out_105_(sb_2__2__0_chany_bottom_out_105_[0]),
		.chany_bottom_out_107_(sb_2__2__0_chany_bottom_out_107_[0]),
		.chany_bottom_out_109_(sb_2__2__0_chany_bottom_out_109_[0]),
		.chany_bottom_out_111_(sb_2__2__0_chany_bottom_out_111_[0]),
		.chany_bottom_out_113_(sb_2__2__0_chany_bottom_out_113_[0]),
		.chany_bottom_out_115_(sb_2__2__0_chany_bottom_out_115_[0]),
		.chany_bottom_out_117_(sb_2__2__0_chany_bottom_out_117_[0]),
		.chany_bottom_out_119_(sb_2__2__0_chany_bottom_out_119_[0]),
		.chany_bottom_out_121_(sb_2__2__0_chany_bottom_out_121_[0]),
		.chany_bottom_out_123_(sb_2__2__0_chany_bottom_out_123_[0]),
		.chany_bottom_out_125_(sb_2__2__0_chany_bottom_out_125_[0]),
		.chany_bottom_out_127_(sb_2__2__0_chany_bottom_out_127_[0]),
		.chany_bottom_out_129_(sb_2__2__0_chany_bottom_out_129_[0]),
		.chany_bottom_out_131_(sb_2__2__0_chany_bottom_out_131_[0]),
		.chany_bottom_out_133_(sb_2__2__0_chany_bottom_out_133_[0]),
		.chany_bottom_out_135_(sb_2__2__0_chany_bottom_out_135_[0]),
		.chany_bottom_out_137_(sb_2__2__0_chany_bottom_out_137_[0]),
		.chany_bottom_out_139_(sb_2__2__0_chany_bottom_out_139_[0]),
		.chany_bottom_out_141_(sb_2__2__0_chany_bottom_out_141_[0]),
		.chany_bottom_out_143_(sb_2__2__0_chany_bottom_out_143_[0]),
		.chany_bottom_out_145_(sb_2__2__0_chany_bottom_out_145_[0]),
		.chany_bottom_out_147_(sb_2__2__0_chany_bottom_out_147_[0]),
		.chany_bottom_out_149_(sb_2__2__0_chany_bottom_out_149_[0]),
		.chany_bottom_out_151_(sb_2__2__0_chany_bottom_out_151_[0]),
		.chany_bottom_out_153_(sb_2__2__0_chany_bottom_out_153_[0]),
		.chany_bottom_out_155_(sb_2__2__0_chany_bottom_out_155_[0]),
		.chany_bottom_out_157_(sb_2__2__0_chany_bottom_out_157_[0]),
		.chany_bottom_out_159_(sb_2__2__0_chany_bottom_out_159_[0]),
		.chany_bottom_out_161_(sb_2__2__0_chany_bottom_out_161_[0]),
		.chany_bottom_out_163_(sb_2__2__0_chany_bottom_out_163_[0]),
		.chany_bottom_out_165_(sb_2__2__0_chany_bottom_out_165_[0]),
		.chany_bottom_out_167_(sb_2__2__0_chany_bottom_out_167_[0]),
		.chany_bottom_out_169_(sb_2__2__0_chany_bottom_out_169_[0]),
		.chany_bottom_out_171_(sb_2__2__0_chany_bottom_out_171_[0]),
		.chany_bottom_out_173_(sb_2__2__0_chany_bottom_out_173_[0]),
		.chany_bottom_out_175_(sb_2__2__0_chany_bottom_out_175_[0]),
		.chany_bottom_out_177_(sb_2__2__0_chany_bottom_out_177_[0]),
		.chany_bottom_out_179_(sb_2__2__0_chany_bottom_out_179_[0]),
		.chany_bottom_out_181_(sb_2__2__0_chany_bottom_out_181_[0]),
		.chany_bottom_out_183_(sb_2__2__0_chany_bottom_out_183_[0]),
		.chany_bottom_out_185_(sb_2__2__0_chany_bottom_out_185_[0]),
		.chany_bottom_out_187_(sb_2__2__0_chany_bottom_out_187_[0]),
		.chany_bottom_out_189_(sb_2__2__0_chany_bottom_out_189_[0]),
		.chany_bottom_out_191_(sb_2__2__0_chany_bottom_out_191_[0]),
		.chany_bottom_out_193_(sb_2__2__0_chany_bottom_out_193_[0]),
		.chany_bottom_out_195_(sb_2__2__0_chany_bottom_out_195_[0]),
		.chany_bottom_out_197_(sb_2__2__0_chany_bottom_out_197_[0]),
		.chany_bottom_out_199_(sb_2__2__0_chany_bottom_out_199_[0]),
		.chanx_left_out_1_(sb_2__2__0_chanx_left_out_1_[0]),
		.chanx_left_out_3_(sb_2__2__0_chanx_left_out_3_[0]),
		.chanx_left_out_5_(sb_2__2__0_chanx_left_out_5_[0]),
		.chanx_left_out_7_(sb_2__2__0_chanx_left_out_7_[0]),
		.chanx_left_out_9_(sb_2__2__0_chanx_left_out_9_[0]),
		.chanx_left_out_11_(sb_2__2__0_chanx_left_out_11_[0]),
		.chanx_left_out_13_(sb_2__2__0_chanx_left_out_13_[0]),
		.chanx_left_out_15_(sb_2__2__0_chanx_left_out_15_[0]),
		.chanx_left_out_17_(sb_2__2__0_chanx_left_out_17_[0]),
		.chanx_left_out_19_(sb_2__2__0_chanx_left_out_19_[0]),
		.chanx_left_out_21_(sb_2__2__0_chanx_left_out_21_[0]),
		.chanx_left_out_23_(sb_2__2__0_chanx_left_out_23_[0]),
		.chanx_left_out_25_(sb_2__2__0_chanx_left_out_25_[0]),
		.chanx_left_out_27_(sb_2__2__0_chanx_left_out_27_[0]),
		.chanx_left_out_29_(sb_2__2__0_chanx_left_out_29_[0]),
		.chanx_left_out_31_(sb_2__2__0_chanx_left_out_31_[0]),
		.chanx_left_out_33_(sb_2__2__0_chanx_left_out_33_[0]),
		.chanx_left_out_35_(sb_2__2__0_chanx_left_out_35_[0]),
		.chanx_left_out_37_(sb_2__2__0_chanx_left_out_37_[0]),
		.chanx_left_out_39_(sb_2__2__0_chanx_left_out_39_[0]),
		.chanx_left_out_41_(sb_2__2__0_chanx_left_out_41_[0]),
		.chanx_left_out_43_(sb_2__2__0_chanx_left_out_43_[0]),
		.chanx_left_out_45_(sb_2__2__0_chanx_left_out_45_[0]),
		.chanx_left_out_47_(sb_2__2__0_chanx_left_out_47_[0]),
		.chanx_left_out_49_(sb_2__2__0_chanx_left_out_49_[0]),
		.chanx_left_out_51_(sb_2__2__0_chanx_left_out_51_[0]),
		.chanx_left_out_53_(sb_2__2__0_chanx_left_out_53_[0]),
		.chanx_left_out_55_(sb_2__2__0_chanx_left_out_55_[0]),
		.chanx_left_out_57_(sb_2__2__0_chanx_left_out_57_[0]),
		.chanx_left_out_59_(sb_2__2__0_chanx_left_out_59_[0]),
		.chanx_left_out_61_(sb_2__2__0_chanx_left_out_61_[0]),
		.chanx_left_out_63_(sb_2__2__0_chanx_left_out_63_[0]),
		.chanx_left_out_65_(sb_2__2__0_chanx_left_out_65_[0]),
		.chanx_left_out_67_(sb_2__2__0_chanx_left_out_67_[0]),
		.chanx_left_out_69_(sb_2__2__0_chanx_left_out_69_[0]),
		.chanx_left_out_71_(sb_2__2__0_chanx_left_out_71_[0]),
		.chanx_left_out_73_(sb_2__2__0_chanx_left_out_73_[0]),
		.chanx_left_out_75_(sb_2__2__0_chanx_left_out_75_[0]),
		.chanx_left_out_77_(sb_2__2__0_chanx_left_out_77_[0]),
		.chanx_left_out_79_(sb_2__2__0_chanx_left_out_79_[0]),
		.chanx_left_out_81_(sb_2__2__0_chanx_left_out_81_[0]),
		.chanx_left_out_83_(sb_2__2__0_chanx_left_out_83_[0]),
		.chanx_left_out_85_(sb_2__2__0_chanx_left_out_85_[0]),
		.chanx_left_out_87_(sb_2__2__0_chanx_left_out_87_[0]),
		.chanx_left_out_89_(sb_2__2__0_chanx_left_out_89_[0]),
		.chanx_left_out_91_(sb_2__2__0_chanx_left_out_91_[0]),
		.chanx_left_out_93_(sb_2__2__0_chanx_left_out_93_[0]),
		.chanx_left_out_95_(sb_2__2__0_chanx_left_out_95_[0]),
		.chanx_left_out_97_(sb_2__2__0_chanx_left_out_97_[0]),
		.chanx_left_out_99_(sb_2__2__0_chanx_left_out_99_[0]),
		.chanx_left_out_101_(sb_2__2__0_chanx_left_out_101_[0]),
		.chanx_left_out_103_(sb_2__2__0_chanx_left_out_103_[0]),
		.chanx_left_out_105_(sb_2__2__0_chanx_left_out_105_[0]),
		.chanx_left_out_107_(sb_2__2__0_chanx_left_out_107_[0]),
		.chanx_left_out_109_(sb_2__2__0_chanx_left_out_109_[0]),
		.chanx_left_out_111_(sb_2__2__0_chanx_left_out_111_[0]),
		.chanx_left_out_113_(sb_2__2__0_chanx_left_out_113_[0]),
		.chanx_left_out_115_(sb_2__2__0_chanx_left_out_115_[0]),
		.chanx_left_out_117_(sb_2__2__0_chanx_left_out_117_[0]),
		.chanx_left_out_119_(sb_2__2__0_chanx_left_out_119_[0]),
		.chanx_left_out_121_(sb_2__2__0_chanx_left_out_121_[0]),
		.chanx_left_out_123_(sb_2__2__0_chanx_left_out_123_[0]),
		.chanx_left_out_125_(sb_2__2__0_chanx_left_out_125_[0]),
		.chanx_left_out_127_(sb_2__2__0_chanx_left_out_127_[0]),
		.chanx_left_out_129_(sb_2__2__0_chanx_left_out_129_[0]),
		.chanx_left_out_131_(sb_2__2__0_chanx_left_out_131_[0]),
		.chanx_left_out_133_(sb_2__2__0_chanx_left_out_133_[0]),
		.chanx_left_out_135_(sb_2__2__0_chanx_left_out_135_[0]),
		.chanx_left_out_137_(sb_2__2__0_chanx_left_out_137_[0]),
		.chanx_left_out_139_(sb_2__2__0_chanx_left_out_139_[0]),
		.chanx_left_out_141_(sb_2__2__0_chanx_left_out_141_[0]),
		.chanx_left_out_143_(sb_2__2__0_chanx_left_out_143_[0]),
		.chanx_left_out_145_(sb_2__2__0_chanx_left_out_145_[0]),
		.chanx_left_out_147_(sb_2__2__0_chanx_left_out_147_[0]),
		.chanx_left_out_149_(sb_2__2__0_chanx_left_out_149_[0]),
		.chanx_left_out_151_(sb_2__2__0_chanx_left_out_151_[0]),
		.chanx_left_out_153_(sb_2__2__0_chanx_left_out_153_[0]),
		.chanx_left_out_155_(sb_2__2__0_chanx_left_out_155_[0]),
		.chanx_left_out_157_(sb_2__2__0_chanx_left_out_157_[0]),
		.chanx_left_out_159_(sb_2__2__0_chanx_left_out_159_[0]),
		.chanx_left_out_161_(sb_2__2__0_chanx_left_out_161_[0]),
		.chanx_left_out_163_(sb_2__2__0_chanx_left_out_163_[0]),
		.chanx_left_out_165_(sb_2__2__0_chanx_left_out_165_[0]),
		.chanx_left_out_167_(sb_2__2__0_chanx_left_out_167_[0]),
		.chanx_left_out_169_(sb_2__2__0_chanx_left_out_169_[0]),
		.chanx_left_out_171_(sb_2__2__0_chanx_left_out_171_[0]),
		.chanx_left_out_173_(sb_2__2__0_chanx_left_out_173_[0]),
		.chanx_left_out_175_(sb_2__2__0_chanx_left_out_175_[0]),
		.chanx_left_out_177_(sb_2__2__0_chanx_left_out_177_[0]),
		.chanx_left_out_179_(sb_2__2__0_chanx_left_out_179_[0]),
		.chanx_left_out_181_(sb_2__2__0_chanx_left_out_181_[0]),
		.chanx_left_out_183_(sb_2__2__0_chanx_left_out_183_[0]),
		.chanx_left_out_185_(sb_2__2__0_chanx_left_out_185_[0]),
		.chanx_left_out_187_(sb_2__2__0_chanx_left_out_187_[0]),
		.chanx_left_out_189_(sb_2__2__0_chanx_left_out_189_[0]),
		.chanx_left_out_191_(sb_2__2__0_chanx_left_out_191_[0]),
		.chanx_left_out_193_(sb_2__2__0_chanx_left_out_193_[0]),
		.chanx_left_out_195_(sb_2__2__0_chanx_left_out_195_[0]),
		.chanx_left_out_197_(sb_2__2__0_chanx_left_out_197_[0]),
		.chanx_left_out_199_(sb_2__2__0_chanx_left_out_199_[0]),
		.ccff_tail(sb_2__2__0_ccff_tail[0]));

	cbx_1__0_ cbx_1__0_ (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.chanx_in_0_(sb_0__0__0_chanx_right_out_0_[0]),
		.chanx_in_1_(sb_1__0__0_chanx_left_out_1_[0]),
		.chanx_in_2_(sb_0__0__0_chanx_right_out_2_[0]),
		.chanx_in_3_(sb_1__0__0_chanx_left_out_3_[0]),
		.chanx_in_4_(sb_0__0__0_chanx_right_out_4_[0]),
		.chanx_in_5_(sb_1__0__0_chanx_left_out_5_[0]),
		.chanx_in_6_(sb_0__0__0_chanx_right_out_6_[0]),
		.chanx_in_7_(sb_1__0__0_chanx_left_out_7_[0]),
		.chanx_in_8_(sb_0__0__0_chanx_right_out_8_[0]),
		.chanx_in_9_(sb_1__0__0_chanx_left_out_9_[0]),
		.chanx_in_10_(sb_0__0__0_chanx_right_out_10_[0]),
		.chanx_in_11_(sb_1__0__0_chanx_left_out_11_[0]),
		.chanx_in_12_(sb_0__0__0_chanx_right_out_12_[0]),
		.chanx_in_13_(sb_1__0__0_chanx_left_out_13_[0]),
		.chanx_in_14_(sb_0__0__0_chanx_right_out_14_[0]),
		.chanx_in_15_(sb_1__0__0_chanx_left_out_15_[0]),
		.chanx_in_16_(sb_0__0__0_chanx_right_out_16_[0]),
		.chanx_in_17_(sb_1__0__0_chanx_left_out_17_[0]),
		.chanx_in_18_(sb_0__0__0_chanx_right_out_18_[0]),
		.chanx_in_19_(sb_1__0__0_chanx_left_out_19_[0]),
		.chanx_in_20_(sb_0__0__0_chanx_right_out_20_[0]),
		.chanx_in_21_(sb_1__0__0_chanx_left_out_21_[0]),
		.chanx_in_22_(sb_0__0__0_chanx_right_out_22_[0]),
		.chanx_in_23_(sb_1__0__0_chanx_left_out_23_[0]),
		.chanx_in_24_(sb_0__0__0_chanx_right_out_24_[0]),
		.chanx_in_25_(sb_1__0__0_chanx_left_out_25_[0]),
		.chanx_in_26_(sb_0__0__0_chanx_right_out_26_[0]),
		.chanx_in_27_(sb_1__0__0_chanx_left_out_27_[0]),
		.chanx_in_28_(sb_0__0__0_chanx_right_out_28_[0]),
		.chanx_in_29_(sb_1__0__0_chanx_left_out_29_[0]),
		.chanx_in_30_(sb_0__0__0_chanx_right_out_30_[0]),
		.chanx_in_31_(sb_1__0__0_chanx_left_out_31_[0]),
		.chanx_in_32_(sb_0__0__0_chanx_right_out_32_[0]),
		.chanx_in_33_(sb_1__0__0_chanx_left_out_33_[0]),
		.chanx_in_34_(sb_0__0__0_chanx_right_out_34_[0]),
		.chanx_in_35_(sb_1__0__0_chanx_left_out_35_[0]),
		.chanx_in_36_(sb_0__0__0_chanx_right_out_36_[0]),
		.chanx_in_37_(sb_1__0__0_chanx_left_out_37_[0]),
		.chanx_in_38_(sb_0__0__0_chanx_right_out_38_[0]),
		.chanx_in_39_(sb_1__0__0_chanx_left_out_39_[0]),
		.chanx_in_40_(sb_0__0__0_chanx_right_out_40_[0]),
		.chanx_in_41_(sb_1__0__0_chanx_left_out_41_[0]),
		.chanx_in_42_(sb_0__0__0_chanx_right_out_42_[0]),
		.chanx_in_43_(sb_1__0__0_chanx_left_out_43_[0]),
		.chanx_in_44_(sb_0__0__0_chanx_right_out_44_[0]),
		.chanx_in_45_(sb_1__0__0_chanx_left_out_45_[0]),
		.chanx_in_46_(sb_0__0__0_chanx_right_out_46_[0]),
		.chanx_in_47_(sb_1__0__0_chanx_left_out_47_[0]),
		.chanx_in_48_(sb_0__0__0_chanx_right_out_48_[0]),
		.chanx_in_49_(sb_1__0__0_chanx_left_out_49_[0]),
		.chanx_in_50_(sb_0__0__0_chanx_right_out_50_[0]),
		.chanx_in_51_(sb_1__0__0_chanx_left_out_51_[0]),
		.chanx_in_52_(sb_0__0__0_chanx_right_out_52_[0]),
		.chanx_in_53_(sb_1__0__0_chanx_left_out_53_[0]),
		.chanx_in_54_(sb_0__0__0_chanx_right_out_54_[0]),
		.chanx_in_55_(sb_1__0__0_chanx_left_out_55_[0]),
		.chanx_in_56_(sb_0__0__0_chanx_right_out_56_[0]),
		.chanx_in_57_(sb_1__0__0_chanx_left_out_57_[0]),
		.chanx_in_58_(sb_0__0__0_chanx_right_out_58_[0]),
		.chanx_in_59_(sb_1__0__0_chanx_left_out_59_[0]),
		.chanx_in_60_(sb_0__0__0_chanx_right_out_60_[0]),
		.chanx_in_61_(sb_1__0__0_chanx_left_out_61_[0]),
		.chanx_in_62_(sb_0__0__0_chanx_right_out_62_[0]),
		.chanx_in_63_(sb_1__0__0_chanx_left_out_63_[0]),
		.chanx_in_64_(sb_0__0__0_chanx_right_out_64_[0]),
		.chanx_in_65_(sb_1__0__0_chanx_left_out_65_[0]),
		.chanx_in_66_(sb_0__0__0_chanx_right_out_66_[0]),
		.chanx_in_67_(sb_1__0__0_chanx_left_out_67_[0]),
		.chanx_in_68_(sb_0__0__0_chanx_right_out_68_[0]),
		.chanx_in_69_(sb_1__0__0_chanx_left_out_69_[0]),
		.chanx_in_70_(sb_0__0__0_chanx_right_out_70_[0]),
		.chanx_in_71_(sb_1__0__0_chanx_left_out_71_[0]),
		.chanx_in_72_(sb_0__0__0_chanx_right_out_72_[0]),
		.chanx_in_73_(sb_1__0__0_chanx_left_out_73_[0]),
		.chanx_in_74_(sb_0__0__0_chanx_right_out_74_[0]),
		.chanx_in_75_(sb_1__0__0_chanx_left_out_75_[0]),
		.chanx_in_76_(sb_0__0__0_chanx_right_out_76_[0]),
		.chanx_in_77_(sb_1__0__0_chanx_left_out_77_[0]),
		.chanx_in_78_(sb_0__0__0_chanx_right_out_78_[0]),
		.chanx_in_79_(sb_1__0__0_chanx_left_out_79_[0]),
		.chanx_in_80_(sb_0__0__0_chanx_right_out_80_[0]),
		.chanx_in_81_(sb_1__0__0_chanx_left_out_81_[0]),
		.chanx_in_82_(sb_0__0__0_chanx_right_out_82_[0]),
		.chanx_in_83_(sb_1__0__0_chanx_left_out_83_[0]),
		.chanx_in_84_(sb_0__0__0_chanx_right_out_84_[0]),
		.chanx_in_85_(sb_1__0__0_chanx_left_out_85_[0]),
		.chanx_in_86_(sb_0__0__0_chanx_right_out_86_[0]),
		.chanx_in_87_(sb_1__0__0_chanx_left_out_87_[0]),
		.chanx_in_88_(sb_0__0__0_chanx_right_out_88_[0]),
		.chanx_in_89_(sb_1__0__0_chanx_left_out_89_[0]),
		.chanx_in_90_(sb_0__0__0_chanx_right_out_90_[0]),
		.chanx_in_91_(sb_1__0__0_chanx_left_out_91_[0]),
		.chanx_in_92_(sb_0__0__0_chanx_right_out_92_[0]),
		.chanx_in_93_(sb_1__0__0_chanx_left_out_93_[0]),
		.chanx_in_94_(sb_0__0__0_chanx_right_out_94_[0]),
		.chanx_in_95_(sb_1__0__0_chanx_left_out_95_[0]),
		.chanx_in_96_(sb_0__0__0_chanx_right_out_96_[0]),
		.chanx_in_97_(sb_1__0__0_chanx_left_out_97_[0]),
		.chanx_in_98_(sb_0__0__0_chanx_right_out_98_[0]),
		.chanx_in_99_(sb_1__0__0_chanx_left_out_99_[0]),
		.chanx_in_100_(sb_0__0__0_chanx_right_out_100_[0]),
		.chanx_in_101_(sb_1__0__0_chanx_left_out_101_[0]),
		.chanx_in_102_(sb_0__0__0_chanx_right_out_102_[0]),
		.chanx_in_103_(sb_1__0__0_chanx_left_out_103_[0]),
		.chanx_in_104_(sb_0__0__0_chanx_right_out_104_[0]),
		.chanx_in_105_(sb_1__0__0_chanx_left_out_105_[0]),
		.chanx_in_106_(sb_0__0__0_chanx_right_out_106_[0]),
		.chanx_in_107_(sb_1__0__0_chanx_left_out_107_[0]),
		.chanx_in_108_(sb_0__0__0_chanx_right_out_108_[0]),
		.chanx_in_109_(sb_1__0__0_chanx_left_out_109_[0]),
		.chanx_in_110_(sb_0__0__0_chanx_right_out_110_[0]),
		.chanx_in_111_(sb_1__0__0_chanx_left_out_111_[0]),
		.chanx_in_112_(sb_0__0__0_chanx_right_out_112_[0]),
		.chanx_in_113_(sb_1__0__0_chanx_left_out_113_[0]),
		.chanx_in_114_(sb_0__0__0_chanx_right_out_114_[0]),
		.chanx_in_115_(sb_1__0__0_chanx_left_out_115_[0]),
		.chanx_in_116_(sb_0__0__0_chanx_right_out_116_[0]),
		.chanx_in_117_(sb_1__0__0_chanx_left_out_117_[0]),
		.chanx_in_118_(sb_0__0__0_chanx_right_out_118_[0]),
		.chanx_in_119_(sb_1__0__0_chanx_left_out_119_[0]),
		.chanx_in_120_(sb_0__0__0_chanx_right_out_120_[0]),
		.chanx_in_121_(sb_1__0__0_chanx_left_out_121_[0]),
		.chanx_in_122_(sb_0__0__0_chanx_right_out_122_[0]),
		.chanx_in_123_(sb_1__0__0_chanx_left_out_123_[0]),
		.chanx_in_124_(sb_0__0__0_chanx_right_out_124_[0]),
		.chanx_in_125_(sb_1__0__0_chanx_left_out_125_[0]),
		.chanx_in_126_(sb_0__0__0_chanx_right_out_126_[0]),
		.chanx_in_127_(sb_1__0__0_chanx_left_out_127_[0]),
		.chanx_in_128_(sb_0__0__0_chanx_right_out_128_[0]),
		.chanx_in_129_(sb_1__0__0_chanx_left_out_129_[0]),
		.chanx_in_130_(sb_0__0__0_chanx_right_out_130_[0]),
		.chanx_in_131_(sb_1__0__0_chanx_left_out_131_[0]),
		.chanx_in_132_(sb_0__0__0_chanx_right_out_132_[0]),
		.chanx_in_133_(sb_1__0__0_chanx_left_out_133_[0]),
		.chanx_in_134_(sb_0__0__0_chanx_right_out_134_[0]),
		.chanx_in_135_(sb_1__0__0_chanx_left_out_135_[0]),
		.chanx_in_136_(sb_0__0__0_chanx_right_out_136_[0]),
		.chanx_in_137_(sb_1__0__0_chanx_left_out_137_[0]),
		.chanx_in_138_(sb_0__0__0_chanx_right_out_138_[0]),
		.chanx_in_139_(sb_1__0__0_chanx_left_out_139_[0]),
		.chanx_in_140_(sb_0__0__0_chanx_right_out_140_[0]),
		.chanx_in_141_(sb_1__0__0_chanx_left_out_141_[0]),
		.chanx_in_142_(sb_0__0__0_chanx_right_out_142_[0]),
		.chanx_in_143_(sb_1__0__0_chanx_left_out_143_[0]),
		.chanx_in_144_(sb_0__0__0_chanx_right_out_144_[0]),
		.chanx_in_145_(sb_1__0__0_chanx_left_out_145_[0]),
		.chanx_in_146_(sb_0__0__0_chanx_right_out_146_[0]),
		.chanx_in_147_(sb_1__0__0_chanx_left_out_147_[0]),
		.chanx_in_148_(sb_0__0__0_chanx_right_out_148_[0]),
		.chanx_in_149_(sb_1__0__0_chanx_left_out_149_[0]),
		.chanx_in_150_(sb_0__0__0_chanx_right_out_150_[0]),
		.chanx_in_151_(sb_1__0__0_chanx_left_out_151_[0]),
		.chanx_in_152_(sb_0__0__0_chanx_right_out_152_[0]),
		.chanx_in_153_(sb_1__0__0_chanx_left_out_153_[0]),
		.chanx_in_154_(sb_0__0__0_chanx_right_out_154_[0]),
		.chanx_in_155_(sb_1__0__0_chanx_left_out_155_[0]),
		.chanx_in_156_(sb_0__0__0_chanx_right_out_156_[0]),
		.chanx_in_157_(sb_1__0__0_chanx_left_out_157_[0]),
		.chanx_in_158_(sb_0__0__0_chanx_right_out_158_[0]),
		.chanx_in_159_(sb_1__0__0_chanx_left_out_159_[0]),
		.chanx_in_160_(sb_0__0__0_chanx_right_out_160_[0]),
		.chanx_in_161_(sb_1__0__0_chanx_left_out_161_[0]),
		.chanx_in_162_(sb_0__0__0_chanx_right_out_162_[0]),
		.chanx_in_163_(sb_1__0__0_chanx_left_out_163_[0]),
		.chanx_in_164_(sb_0__0__0_chanx_right_out_164_[0]),
		.chanx_in_165_(sb_1__0__0_chanx_left_out_165_[0]),
		.chanx_in_166_(sb_0__0__0_chanx_right_out_166_[0]),
		.chanx_in_167_(sb_1__0__0_chanx_left_out_167_[0]),
		.chanx_in_168_(sb_0__0__0_chanx_right_out_168_[0]),
		.chanx_in_169_(sb_1__0__0_chanx_left_out_169_[0]),
		.chanx_in_170_(sb_0__0__0_chanx_right_out_170_[0]),
		.chanx_in_171_(sb_1__0__0_chanx_left_out_171_[0]),
		.chanx_in_172_(sb_0__0__0_chanx_right_out_172_[0]),
		.chanx_in_173_(sb_1__0__0_chanx_left_out_173_[0]),
		.chanx_in_174_(sb_0__0__0_chanx_right_out_174_[0]),
		.chanx_in_175_(sb_1__0__0_chanx_left_out_175_[0]),
		.chanx_in_176_(sb_0__0__0_chanx_right_out_176_[0]),
		.chanx_in_177_(sb_1__0__0_chanx_left_out_177_[0]),
		.chanx_in_178_(sb_0__0__0_chanx_right_out_178_[0]),
		.chanx_in_179_(sb_1__0__0_chanx_left_out_179_[0]),
		.chanx_in_180_(sb_0__0__0_chanx_right_out_180_[0]),
		.chanx_in_181_(sb_1__0__0_chanx_left_out_181_[0]),
		.chanx_in_182_(sb_0__0__0_chanx_right_out_182_[0]),
		.chanx_in_183_(sb_1__0__0_chanx_left_out_183_[0]),
		.chanx_in_184_(sb_0__0__0_chanx_right_out_184_[0]),
		.chanx_in_185_(sb_1__0__0_chanx_left_out_185_[0]),
		.chanx_in_186_(sb_0__0__0_chanx_right_out_186_[0]),
		.chanx_in_187_(sb_1__0__0_chanx_left_out_187_[0]),
		.chanx_in_188_(sb_0__0__0_chanx_right_out_188_[0]),
		.chanx_in_189_(sb_1__0__0_chanx_left_out_189_[0]),
		.chanx_in_190_(sb_0__0__0_chanx_right_out_190_[0]),
		.chanx_in_191_(sb_1__0__0_chanx_left_out_191_[0]),
		.chanx_in_192_(sb_0__0__0_chanx_right_out_192_[0]),
		.chanx_in_193_(sb_1__0__0_chanx_left_out_193_[0]),
		.chanx_in_194_(sb_0__0__0_chanx_right_out_194_[0]),
		.chanx_in_195_(sb_1__0__0_chanx_left_out_195_[0]),
		.chanx_in_196_(sb_0__0__0_chanx_right_out_196_[0]),
		.chanx_in_197_(sb_1__0__0_chanx_left_out_197_[0]),
		.chanx_in_198_(sb_0__0__0_chanx_right_out_198_[0]),
		.chanx_in_199_(sb_1__0__0_chanx_left_out_199_[0]),
		.ccff_head(sb_1__0__0_ccff_tail[0]),
		.chanx_out_0_(cbx_1__0__0_chanx_out_0_[0]),
		.chanx_out_1_(cbx_1__0__0_chanx_out_1_[0]),
		.chanx_out_2_(cbx_1__0__0_chanx_out_2_[0]),
		.chanx_out_3_(cbx_1__0__0_chanx_out_3_[0]),
		.chanx_out_4_(cbx_1__0__0_chanx_out_4_[0]),
		.chanx_out_5_(cbx_1__0__0_chanx_out_5_[0]),
		.chanx_out_6_(cbx_1__0__0_chanx_out_6_[0]),
		.chanx_out_7_(cbx_1__0__0_chanx_out_7_[0]),
		.chanx_out_8_(cbx_1__0__0_chanx_out_8_[0]),
		.chanx_out_9_(cbx_1__0__0_chanx_out_9_[0]),
		.chanx_out_10_(cbx_1__0__0_chanx_out_10_[0]),
		.chanx_out_11_(cbx_1__0__0_chanx_out_11_[0]),
		.chanx_out_12_(cbx_1__0__0_chanx_out_12_[0]),
		.chanx_out_13_(cbx_1__0__0_chanx_out_13_[0]),
		.chanx_out_14_(cbx_1__0__0_chanx_out_14_[0]),
		.chanx_out_15_(cbx_1__0__0_chanx_out_15_[0]),
		.chanx_out_16_(cbx_1__0__0_chanx_out_16_[0]),
		.chanx_out_17_(cbx_1__0__0_chanx_out_17_[0]),
		.chanx_out_18_(cbx_1__0__0_chanx_out_18_[0]),
		.chanx_out_19_(cbx_1__0__0_chanx_out_19_[0]),
		.chanx_out_20_(cbx_1__0__0_chanx_out_20_[0]),
		.chanx_out_21_(cbx_1__0__0_chanx_out_21_[0]),
		.chanx_out_22_(cbx_1__0__0_chanx_out_22_[0]),
		.chanx_out_23_(cbx_1__0__0_chanx_out_23_[0]),
		.chanx_out_24_(cbx_1__0__0_chanx_out_24_[0]),
		.chanx_out_25_(cbx_1__0__0_chanx_out_25_[0]),
		.chanx_out_26_(cbx_1__0__0_chanx_out_26_[0]),
		.chanx_out_27_(cbx_1__0__0_chanx_out_27_[0]),
		.chanx_out_28_(cbx_1__0__0_chanx_out_28_[0]),
		.chanx_out_29_(cbx_1__0__0_chanx_out_29_[0]),
		.chanx_out_30_(cbx_1__0__0_chanx_out_30_[0]),
		.chanx_out_31_(cbx_1__0__0_chanx_out_31_[0]),
		.chanx_out_32_(cbx_1__0__0_chanx_out_32_[0]),
		.chanx_out_33_(cbx_1__0__0_chanx_out_33_[0]),
		.chanx_out_34_(cbx_1__0__0_chanx_out_34_[0]),
		.chanx_out_35_(cbx_1__0__0_chanx_out_35_[0]),
		.chanx_out_36_(cbx_1__0__0_chanx_out_36_[0]),
		.chanx_out_37_(cbx_1__0__0_chanx_out_37_[0]),
		.chanx_out_38_(cbx_1__0__0_chanx_out_38_[0]),
		.chanx_out_39_(cbx_1__0__0_chanx_out_39_[0]),
		.chanx_out_40_(cbx_1__0__0_chanx_out_40_[0]),
		.chanx_out_41_(cbx_1__0__0_chanx_out_41_[0]),
		.chanx_out_42_(cbx_1__0__0_chanx_out_42_[0]),
		.chanx_out_43_(cbx_1__0__0_chanx_out_43_[0]),
		.chanx_out_44_(cbx_1__0__0_chanx_out_44_[0]),
		.chanx_out_45_(cbx_1__0__0_chanx_out_45_[0]),
		.chanx_out_46_(cbx_1__0__0_chanx_out_46_[0]),
		.chanx_out_47_(cbx_1__0__0_chanx_out_47_[0]),
		.chanx_out_48_(cbx_1__0__0_chanx_out_48_[0]),
		.chanx_out_49_(cbx_1__0__0_chanx_out_49_[0]),
		.chanx_out_50_(cbx_1__0__0_chanx_out_50_[0]),
		.chanx_out_51_(cbx_1__0__0_chanx_out_51_[0]),
		.chanx_out_52_(cbx_1__0__0_chanx_out_52_[0]),
		.chanx_out_53_(cbx_1__0__0_chanx_out_53_[0]),
		.chanx_out_54_(cbx_1__0__0_chanx_out_54_[0]),
		.chanx_out_55_(cbx_1__0__0_chanx_out_55_[0]),
		.chanx_out_56_(cbx_1__0__0_chanx_out_56_[0]),
		.chanx_out_57_(cbx_1__0__0_chanx_out_57_[0]),
		.chanx_out_58_(cbx_1__0__0_chanx_out_58_[0]),
		.chanx_out_59_(cbx_1__0__0_chanx_out_59_[0]),
		.chanx_out_60_(cbx_1__0__0_chanx_out_60_[0]),
		.chanx_out_61_(cbx_1__0__0_chanx_out_61_[0]),
		.chanx_out_62_(cbx_1__0__0_chanx_out_62_[0]),
		.chanx_out_63_(cbx_1__0__0_chanx_out_63_[0]),
		.chanx_out_64_(cbx_1__0__0_chanx_out_64_[0]),
		.chanx_out_65_(cbx_1__0__0_chanx_out_65_[0]),
		.chanx_out_66_(cbx_1__0__0_chanx_out_66_[0]),
		.chanx_out_67_(cbx_1__0__0_chanx_out_67_[0]),
		.chanx_out_68_(cbx_1__0__0_chanx_out_68_[0]),
		.chanx_out_69_(cbx_1__0__0_chanx_out_69_[0]),
		.chanx_out_70_(cbx_1__0__0_chanx_out_70_[0]),
		.chanx_out_71_(cbx_1__0__0_chanx_out_71_[0]),
		.chanx_out_72_(cbx_1__0__0_chanx_out_72_[0]),
		.chanx_out_73_(cbx_1__0__0_chanx_out_73_[0]),
		.chanx_out_74_(cbx_1__0__0_chanx_out_74_[0]),
		.chanx_out_75_(cbx_1__0__0_chanx_out_75_[0]),
		.chanx_out_76_(cbx_1__0__0_chanx_out_76_[0]),
		.chanx_out_77_(cbx_1__0__0_chanx_out_77_[0]),
		.chanx_out_78_(cbx_1__0__0_chanx_out_78_[0]),
		.chanx_out_79_(cbx_1__0__0_chanx_out_79_[0]),
		.chanx_out_80_(cbx_1__0__0_chanx_out_80_[0]),
		.chanx_out_81_(cbx_1__0__0_chanx_out_81_[0]),
		.chanx_out_82_(cbx_1__0__0_chanx_out_82_[0]),
		.chanx_out_83_(cbx_1__0__0_chanx_out_83_[0]),
		.chanx_out_84_(cbx_1__0__0_chanx_out_84_[0]),
		.chanx_out_85_(cbx_1__0__0_chanx_out_85_[0]),
		.chanx_out_86_(cbx_1__0__0_chanx_out_86_[0]),
		.chanx_out_87_(cbx_1__0__0_chanx_out_87_[0]),
		.chanx_out_88_(cbx_1__0__0_chanx_out_88_[0]),
		.chanx_out_89_(cbx_1__0__0_chanx_out_89_[0]),
		.chanx_out_90_(cbx_1__0__0_chanx_out_90_[0]),
		.chanx_out_91_(cbx_1__0__0_chanx_out_91_[0]),
		.chanx_out_92_(cbx_1__0__0_chanx_out_92_[0]),
		.chanx_out_93_(cbx_1__0__0_chanx_out_93_[0]),
		.chanx_out_94_(cbx_1__0__0_chanx_out_94_[0]),
		.chanx_out_95_(cbx_1__0__0_chanx_out_95_[0]),
		.chanx_out_96_(cbx_1__0__0_chanx_out_96_[0]),
		.chanx_out_97_(cbx_1__0__0_chanx_out_97_[0]),
		.chanx_out_98_(cbx_1__0__0_chanx_out_98_[0]),
		.chanx_out_99_(cbx_1__0__0_chanx_out_99_[0]),
		.chanx_out_100_(cbx_1__0__0_chanx_out_100_[0]),
		.chanx_out_101_(cbx_1__0__0_chanx_out_101_[0]),
		.chanx_out_102_(cbx_1__0__0_chanx_out_102_[0]),
		.chanx_out_103_(cbx_1__0__0_chanx_out_103_[0]),
		.chanx_out_104_(cbx_1__0__0_chanx_out_104_[0]),
		.chanx_out_105_(cbx_1__0__0_chanx_out_105_[0]),
		.chanx_out_106_(cbx_1__0__0_chanx_out_106_[0]),
		.chanx_out_107_(cbx_1__0__0_chanx_out_107_[0]),
		.chanx_out_108_(cbx_1__0__0_chanx_out_108_[0]),
		.chanx_out_109_(cbx_1__0__0_chanx_out_109_[0]),
		.chanx_out_110_(cbx_1__0__0_chanx_out_110_[0]),
		.chanx_out_111_(cbx_1__0__0_chanx_out_111_[0]),
		.chanx_out_112_(cbx_1__0__0_chanx_out_112_[0]),
		.chanx_out_113_(cbx_1__0__0_chanx_out_113_[0]),
		.chanx_out_114_(cbx_1__0__0_chanx_out_114_[0]),
		.chanx_out_115_(cbx_1__0__0_chanx_out_115_[0]),
		.chanx_out_116_(cbx_1__0__0_chanx_out_116_[0]),
		.chanx_out_117_(cbx_1__0__0_chanx_out_117_[0]),
		.chanx_out_118_(cbx_1__0__0_chanx_out_118_[0]),
		.chanx_out_119_(cbx_1__0__0_chanx_out_119_[0]),
		.chanx_out_120_(cbx_1__0__0_chanx_out_120_[0]),
		.chanx_out_121_(cbx_1__0__0_chanx_out_121_[0]),
		.chanx_out_122_(cbx_1__0__0_chanx_out_122_[0]),
		.chanx_out_123_(cbx_1__0__0_chanx_out_123_[0]),
		.chanx_out_124_(cbx_1__0__0_chanx_out_124_[0]),
		.chanx_out_125_(cbx_1__0__0_chanx_out_125_[0]),
		.chanx_out_126_(cbx_1__0__0_chanx_out_126_[0]),
		.chanx_out_127_(cbx_1__0__0_chanx_out_127_[0]),
		.chanx_out_128_(cbx_1__0__0_chanx_out_128_[0]),
		.chanx_out_129_(cbx_1__0__0_chanx_out_129_[0]),
		.chanx_out_130_(cbx_1__0__0_chanx_out_130_[0]),
		.chanx_out_131_(cbx_1__0__0_chanx_out_131_[0]),
		.chanx_out_132_(cbx_1__0__0_chanx_out_132_[0]),
		.chanx_out_133_(cbx_1__0__0_chanx_out_133_[0]),
		.chanx_out_134_(cbx_1__0__0_chanx_out_134_[0]),
		.chanx_out_135_(cbx_1__0__0_chanx_out_135_[0]),
		.chanx_out_136_(cbx_1__0__0_chanx_out_136_[0]),
		.chanx_out_137_(cbx_1__0__0_chanx_out_137_[0]),
		.chanx_out_138_(cbx_1__0__0_chanx_out_138_[0]),
		.chanx_out_139_(cbx_1__0__0_chanx_out_139_[0]),
		.chanx_out_140_(cbx_1__0__0_chanx_out_140_[0]),
		.chanx_out_141_(cbx_1__0__0_chanx_out_141_[0]),
		.chanx_out_142_(cbx_1__0__0_chanx_out_142_[0]),
		.chanx_out_143_(cbx_1__0__0_chanx_out_143_[0]),
		.chanx_out_144_(cbx_1__0__0_chanx_out_144_[0]),
		.chanx_out_145_(cbx_1__0__0_chanx_out_145_[0]),
		.chanx_out_146_(cbx_1__0__0_chanx_out_146_[0]),
		.chanx_out_147_(cbx_1__0__0_chanx_out_147_[0]),
		.chanx_out_148_(cbx_1__0__0_chanx_out_148_[0]),
		.chanx_out_149_(cbx_1__0__0_chanx_out_149_[0]),
		.chanx_out_150_(cbx_1__0__0_chanx_out_150_[0]),
		.chanx_out_151_(cbx_1__0__0_chanx_out_151_[0]),
		.chanx_out_152_(cbx_1__0__0_chanx_out_152_[0]),
		.chanx_out_153_(cbx_1__0__0_chanx_out_153_[0]),
		.chanx_out_154_(cbx_1__0__0_chanx_out_154_[0]),
		.chanx_out_155_(cbx_1__0__0_chanx_out_155_[0]),
		.chanx_out_156_(cbx_1__0__0_chanx_out_156_[0]),
		.chanx_out_157_(cbx_1__0__0_chanx_out_157_[0]),
		.chanx_out_158_(cbx_1__0__0_chanx_out_158_[0]),
		.chanx_out_159_(cbx_1__0__0_chanx_out_159_[0]),
		.chanx_out_160_(cbx_1__0__0_chanx_out_160_[0]),
		.chanx_out_161_(cbx_1__0__0_chanx_out_161_[0]),
		.chanx_out_162_(cbx_1__0__0_chanx_out_162_[0]),
		.chanx_out_163_(cbx_1__0__0_chanx_out_163_[0]),
		.chanx_out_164_(cbx_1__0__0_chanx_out_164_[0]),
		.chanx_out_165_(cbx_1__0__0_chanx_out_165_[0]),
		.chanx_out_166_(cbx_1__0__0_chanx_out_166_[0]),
		.chanx_out_167_(cbx_1__0__0_chanx_out_167_[0]),
		.chanx_out_168_(cbx_1__0__0_chanx_out_168_[0]),
		.chanx_out_169_(cbx_1__0__0_chanx_out_169_[0]),
		.chanx_out_170_(cbx_1__0__0_chanx_out_170_[0]),
		.chanx_out_171_(cbx_1__0__0_chanx_out_171_[0]),
		.chanx_out_172_(cbx_1__0__0_chanx_out_172_[0]),
		.chanx_out_173_(cbx_1__0__0_chanx_out_173_[0]),
		.chanx_out_174_(cbx_1__0__0_chanx_out_174_[0]),
		.chanx_out_175_(cbx_1__0__0_chanx_out_175_[0]),
		.chanx_out_176_(cbx_1__0__0_chanx_out_176_[0]),
		.chanx_out_177_(cbx_1__0__0_chanx_out_177_[0]),
		.chanx_out_178_(cbx_1__0__0_chanx_out_178_[0]),
		.chanx_out_179_(cbx_1__0__0_chanx_out_179_[0]),
		.chanx_out_180_(cbx_1__0__0_chanx_out_180_[0]),
		.chanx_out_181_(cbx_1__0__0_chanx_out_181_[0]),
		.chanx_out_182_(cbx_1__0__0_chanx_out_182_[0]),
		.chanx_out_183_(cbx_1__0__0_chanx_out_183_[0]),
		.chanx_out_184_(cbx_1__0__0_chanx_out_184_[0]),
		.chanx_out_185_(cbx_1__0__0_chanx_out_185_[0]),
		.chanx_out_186_(cbx_1__0__0_chanx_out_186_[0]),
		.chanx_out_187_(cbx_1__0__0_chanx_out_187_[0]),
		.chanx_out_188_(cbx_1__0__0_chanx_out_188_[0]),
		.chanx_out_189_(cbx_1__0__0_chanx_out_189_[0]),
		.chanx_out_190_(cbx_1__0__0_chanx_out_190_[0]),
		.chanx_out_191_(cbx_1__0__0_chanx_out_191_[0]),
		.chanx_out_192_(cbx_1__0__0_chanx_out_192_[0]),
		.chanx_out_193_(cbx_1__0__0_chanx_out_193_[0]),
		.chanx_out_194_(cbx_1__0__0_chanx_out_194_[0]),
		.chanx_out_195_(cbx_1__0__0_chanx_out_195_[0]),
		.chanx_out_196_(cbx_1__0__0_chanx_out_196_[0]),
		.chanx_out_197_(cbx_1__0__0_chanx_out_197_[0]),
		.chanx_out_198_(cbx_1__0__0_chanx_out_198_[0]),
		.chanx_out_199_(cbx_1__0__0_chanx_out_199_[0]),
		.top_grid_pin_20_(cbx_1__0__0_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__0__0_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__0__0_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__0__0_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__0__0_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__0__0_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__0__0_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__0__0_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__0__0_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__0__0_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__0__0_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__0__0_top_grid_pin_31_[0]),
		.top_grid_pin_32_(cbx_1__0__0_top_grid_pin_32_[0]),
		.top_grid_pin_33_(cbx_1__0__0_top_grid_pin_33_[0]),
		.top_grid_pin_34_(cbx_1__0__0_top_grid_pin_34_[0]),
		.top_grid_pin_35_(cbx_1__0__0_top_grid_pin_35_[0]),
		.top_grid_pin_36_(cbx_1__0__0_top_grid_pin_36_[0]),
		.top_grid_pin_37_(cbx_1__0__0_top_grid_pin_37_[0]),
		.top_grid_pin_38_(cbx_1__0__0_top_grid_pin_38_[0]),
		.top_grid_pin_39_(cbx_1__0__0_top_grid_pin_39_[0]),
		.bottom_grid_pin_0_(cbx_1__0__0_bottom_grid_pin_0_[0]),
		.ccff_tail(cbx_1__0__0_ccff_tail[0]));

	cbx_1__0_ cbx_2__0_ (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.chanx_in_0_(sb_1__0__0_chanx_right_out_0_[0]),
		.chanx_in_1_(sb_2__0__0_chanx_left_out_1_[0]),
		.chanx_in_2_(sb_1__0__0_chanx_right_out_2_[0]),
		.chanx_in_3_(sb_2__0__0_chanx_left_out_3_[0]),
		.chanx_in_4_(sb_1__0__0_chanx_right_out_4_[0]),
		.chanx_in_5_(sb_2__0__0_chanx_left_out_5_[0]),
		.chanx_in_6_(sb_1__0__0_chanx_right_out_6_[0]),
		.chanx_in_7_(sb_2__0__0_chanx_left_out_7_[0]),
		.chanx_in_8_(sb_1__0__0_chanx_right_out_8_[0]),
		.chanx_in_9_(sb_2__0__0_chanx_left_out_9_[0]),
		.chanx_in_10_(sb_1__0__0_chanx_right_out_10_[0]),
		.chanx_in_11_(sb_2__0__0_chanx_left_out_11_[0]),
		.chanx_in_12_(sb_1__0__0_chanx_right_out_12_[0]),
		.chanx_in_13_(sb_2__0__0_chanx_left_out_13_[0]),
		.chanx_in_14_(sb_1__0__0_chanx_right_out_14_[0]),
		.chanx_in_15_(sb_2__0__0_chanx_left_out_15_[0]),
		.chanx_in_16_(sb_1__0__0_chanx_right_out_16_[0]),
		.chanx_in_17_(sb_2__0__0_chanx_left_out_17_[0]),
		.chanx_in_18_(sb_1__0__0_chanx_right_out_18_[0]),
		.chanx_in_19_(sb_2__0__0_chanx_left_out_19_[0]),
		.chanx_in_20_(sb_1__0__0_chanx_right_out_20_[0]),
		.chanx_in_21_(sb_2__0__0_chanx_left_out_21_[0]),
		.chanx_in_22_(sb_1__0__0_chanx_right_out_22_[0]),
		.chanx_in_23_(sb_2__0__0_chanx_left_out_23_[0]),
		.chanx_in_24_(sb_1__0__0_chanx_right_out_24_[0]),
		.chanx_in_25_(sb_2__0__0_chanx_left_out_25_[0]),
		.chanx_in_26_(sb_1__0__0_chanx_right_out_26_[0]),
		.chanx_in_27_(sb_2__0__0_chanx_left_out_27_[0]),
		.chanx_in_28_(sb_1__0__0_chanx_right_out_28_[0]),
		.chanx_in_29_(sb_2__0__0_chanx_left_out_29_[0]),
		.chanx_in_30_(sb_1__0__0_chanx_right_out_30_[0]),
		.chanx_in_31_(sb_2__0__0_chanx_left_out_31_[0]),
		.chanx_in_32_(sb_1__0__0_chanx_right_out_32_[0]),
		.chanx_in_33_(sb_2__0__0_chanx_left_out_33_[0]),
		.chanx_in_34_(sb_1__0__0_chanx_right_out_34_[0]),
		.chanx_in_35_(sb_2__0__0_chanx_left_out_35_[0]),
		.chanx_in_36_(sb_1__0__0_chanx_right_out_36_[0]),
		.chanx_in_37_(sb_2__0__0_chanx_left_out_37_[0]),
		.chanx_in_38_(sb_1__0__0_chanx_right_out_38_[0]),
		.chanx_in_39_(sb_2__0__0_chanx_left_out_39_[0]),
		.chanx_in_40_(sb_1__0__0_chanx_right_out_40_[0]),
		.chanx_in_41_(sb_2__0__0_chanx_left_out_41_[0]),
		.chanx_in_42_(sb_1__0__0_chanx_right_out_42_[0]),
		.chanx_in_43_(sb_2__0__0_chanx_left_out_43_[0]),
		.chanx_in_44_(sb_1__0__0_chanx_right_out_44_[0]),
		.chanx_in_45_(sb_2__0__0_chanx_left_out_45_[0]),
		.chanx_in_46_(sb_1__0__0_chanx_right_out_46_[0]),
		.chanx_in_47_(sb_2__0__0_chanx_left_out_47_[0]),
		.chanx_in_48_(sb_1__0__0_chanx_right_out_48_[0]),
		.chanx_in_49_(sb_2__0__0_chanx_left_out_49_[0]),
		.chanx_in_50_(sb_1__0__0_chanx_right_out_50_[0]),
		.chanx_in_51_(sb_2__0__0_chanx_left_out_51_[0]),
		.chanx_in_52_(sb_1__0__0_chanx_right_out_52_[0]),
		.chanx_in_53_(sb_2__0__0_chanx_left_out_53_[0]),
		.chanx_in_54_(sb_1__0__0_chanx_right_out_54_[0]),
		.chanx_in_55_(sb_2__0__0_chanx_left_out_55_[0]),
		.chanx_in_56_(sb_1__0__0_chanx_right_out_56_[0]),
		.chanx_in_57_(sb_2__0__0_chanx_left_out_57_[0]),
		.chanx_in_58_(sb_1__0__0_chanx_right_out_58_[0]),
		.chanx_in_59_(sb_2__0__0_chanx_left_out_59_[0]),
		.chanx_in_60_(sb_1__0__0_chanx_right_out_60_[0]),
		.chanx_in_61_(sb_2__0__0_chanx_left_out_61_[0]),
		.chanx_in_62_(sb_1__0__0_chanx_right_out_62_[0]),
		.chanx_in_63_(sb_2__0__0_chanx_left_out_63_[0]),
		.chanx_in_64_(sb_1__0__0_chanx_right_out_64_[0]),
		.chanx_in_65_(sb_2__0__0_chanx_left_out_65_[0]),
		.chanx_in_66_(sb_1__0__0_chanx_right_out_66_[0]),
		.chanx_in_67_(sb_2__0__0_chanx_left_out_67_[0]),
		.chanx_in_68_(sb_1__0__0_chanx_right_out_68_[0]),
		.chanx_in_69_(sb_2__0__0_chanx_left_out_69_[0]),
		.chanx_in_70_(sb_1__0__0_chanx_right_out_70_[0]),
		.chanx_in_71_(sb_2__0__0_chanx_left_out_71_[0]),
		.chanx_in_72_(sb_1__0__0_chanx_right_out_72_[0]),
		.chanx_in_73_(sb_2__0__0_chanx_left_out_73_[0]),
		.chanx_in_74_(sb_1__0__0_chanx_right_out_74_[0]),
		.chanx_in_75_(sb_2__0__0_chanx_left_out_75_[0]),
		.chanx_in_76_(sb_1__0__0_chanx_right_out_76_[0]),
		.chanx_in_77_(sb_2__0__0_chanx_left_out_77_[0]),
		.chanx_in_78_(sb_1__0__0_chanx_right_out_78_[0]),
		.chanx_in_79_(sb_2__0__0_chanx_left_out_79_[0]),
		.chanx_in_80_(sb_1__0__0_chanx_right_out_80_[0]),
		.chanx_in_81_(sb_2__0__0_chanx_left_out_81_[0]),
		.chanx_in_82_(sb_1__0__0_chanx_right_out_82_[0]),
		.chanx_in_83_(sb_2__0__0_chanx_left_out_83_[0]),
		.chanx_in_84_(sb_1__0__0_chanx_right_out_84_[0]),
		.chanx_in_85_(sb_2__0__0_chanx_left_out_85_[0]),
		.chanx_in_86_(sb_1__0__0_chanx_right_out_86_[0]),
		.chanx_in_87_(sb_2__0__0_chanx_left_out_87_[0]),
		.chanx_in_88_(sb_1__0__0_chanx_right_out_88_[0]),
		.chanx_in_89_(sb_2__0__0_chanx_left_out_89_[0]),
		.chanx_in_90_(sb_1__0__0_chanx_right_out_90_[0]),
		.chanx_in_91_(sb_2__0__0_chanx_left_out_91_[0]),
		.chanx_in_92_(sb_1__0__0_chanx_right_out_92_[0]),
		.chanx_in_93_(sb_2__0__0_chanx_left_out_93_[0]),
		.chanx_in_94_(sb_1__0__0_chanx_right_out_94_[0]),
		.chanx_in_95_(sb_2__0__0_chanx_left_out_95_[0]),
		.chanx_in_96_(sb_1__0__0_chanx_right_out_96_[0]),
		.chanx_in_97_(sb_2__0__0_chanx_left_out_97_[0]),
		.chanx_in_98_(sb_1__0__0_chanx_right_out_98_[0]),
		.chanx_in_99_(sb_2__0__0_chanx_left_out_99_[0]),
		.chanx_in_100_(sb_1__0__0_chanx_right_out_100_[0]),
		.chanx_in_101_(sb_2__0__0_chanx_left_out_101_[0]),
		.chanx_in_102_(sb_1__0__0_chanx_right_out_102_[0]),
		.chanx_in_103_(sb_2__0__0_chanx_left_out_103_[0]),
		.chanx_in_104_(sb_1__0__0_chanx_right_out_104_[0]),
		.chanx_in_105_(sb_2__0__0_chanx_left_out_105_[0]),
		.chanx_in_106_(sb_1__0__0_chanx_right_out_106_[0]),
		.chanx_in_107_(sb_2__0__0_chanx_left_out_107_[0]),
		.chanx_in_108_(sb_1__0__0_chanx_right_out_108_[0]),
		.chanx_in_109_(sb_2__0__0_chanx_left_out_109_[0]),
		.chanx_in_110_(sb_1__0__0_chanx_right_out_110_[0]),
		.chanx_in_111_(sb_2__0__0_chanx_left_out_111_[0]),
		.chanx_in_112_(sb_1__0__0_chanx_right_out_112_[0]),
		.chanx_in_113_(sb_2__0__0_chanx_left_out_113_[0]),
		.chanx_in_114_(sb_1__0__0_chanx_right_out_114_[0]),
		.chanx_in_115_(sb_2__0__0_chanx_left_out_115_[0]),
		.chanx_in_116_(sb_1__0__0_chanx_right_out_116_[0]),
		.chanx_in_117_(sb_2__0__0_chanx_left_out_117_[0]),
		.chanx_in_118_(sb_1__0__0_chanx_right_out_118_[0]),
		.chanx_in_119_(sb_2__0__0_chanx_left_out_119_[0]),
		.chanx_in_120_(sb_1__0__0_chanx_right_out_120_[0]),
		.chanx_in_121_(sb_2__0__0_chanx_left_out_121_[0]),
		.chanx_in_122_(sb_1__0__0_chanx_right_out_122_[0]),
		.chanx_in_123_(sb_2__0__0_chanx_left_out_123_[0]),
		.chanx_in_124_(sb_1__0__0_chanx_right_out_124_[0]),
		.chanx_in_125_(sb_2__0__0_chanx_left_out_125_[0]),
		.chanx_in_126_(sb_1__0__0_chanx_right_out_126_[0]),
		.chanx_in_127_(sb_2__0__0_chanx_left_out_127_[0]),
		.chanx_in_128_(sb_1__0__0_chanx_right_out_128_[0]),
		.chanx_in_129_(sb_2__0__0_chanx_left_out_129_[0]),
		.chanx_in_130_(sb_1__0__0_chanx_right_out_130_[0]),
		.chanx_in_131_(sb_2__0__0_chanx_left_out_131_[0]),
		.chanx_in_132_(sb_1__0__0_chanx_right_out_132_[0]),
		.chanx_in_133_(sb_2__0__0_chanx_left_out_133_[0]),
		.chanx_in_134_(sb_1__0__0_chanx_right_out_134_[0]),
		.chanx_in_135_(sb_2__0__0_chanx_left_out_135_[0]),
		.chanx_in_136_(sb_1__0__0_chanx_right_out_136_[0]),
		.chanx_in_137_(sb_2__0__0_chanx_left_out_137_[0]),
		.chanx_in_138_(sb_1__0__0_chanx_right_out_138_[0]),
		.chanx_in_139_(sb_2__0__0_chanx_left_out_139_[0]),
		.chanx_in_140_(sb_1__0__0_chanx_right_out_140_[0]),
		.chanx_in_141_(sb_2__0__0_chanx_left_out_141_[0]),
		.chanx_in_142_(sb_1__0__0_chanx_right_out_142_[0]),
		.chanx_in_143_(sb_2__0__0_chanx_left_out_143_[0]),
		.chanx_in_144_(sb_1__0__0_chanx_right_out_144_[0]),
		.chanx_in_145_(sb_2__0__0_chanx_left_out_145_[0]),
		.chanx_in_146_(sb_1__0__0_chanx_right_out_146_[0]),
		.chanx_in_147_(sb_2__0__0_chanx_left_out_147_[0]),
		.chanx_in_148_(sb_1__0__0_chanx_right_out_148_[0]),
		.chanx_in_149_(sb_2__0__0_chanx_left_out_149_[0]),
		.chanx_in_150_(sb_1__0__0_chanx_right_out_150_[0]),
		.chanx_in_151_(sb_2__0__0_chanx_left_out_151_[0]),
		.chanx_in_152_(sb_1__0__0_chanx_right_out_152_[0]),
		.chanx_in_153_(sb_2__0__0_chanx_left_out_153_[0]),
		.chanx_in_154_(sb_1__0__0_chanx_right_out_154_[0]),
		.chanx_in_155_(sb_2__0__0_chanx_left_out_155_[0]),
		.chanx_in_156_(sb_1__0__0_chanx_right_out_156_[0]),
		.chanx_in_157_(sb_2__0__0_chanx_left_out_157_[0]),
		.chanx_in_158_(sb_1__0__0_chanx_right_out_158_[0]),
		.chanx_in_159_(sb_2__0__0_chanx_left_out_159_[0]),
		.chanx_in_160_(sb_1__0__0_chanx_right_out_160_[0]),
		.chanx_in_161_(sb_2__0__0_chanx_left_out_161_[0]),
		.chanx_in_162_(sb_1__0__0_chanx_right_out_162_[0]),
		.chanx_in_163_(sb_2__0__0_chanx_left_out_163_[0]),
		.chanx_in_164_(sb_1__0__0_chanx_right_out_164_[0]),
		.chanx_in_165_(sb_2__0__0_chanx_left_out_165_[0]),
		.chanx_in_166_(sb_1__0__0_chanx_right_out_166_[0]),
		.chanx_in_167_(sb_2__0__0_chanx_left_out_167_[0]),
		.chanx_in_168_(sb_1__0__0_chanx_right_out_168_[0]),
		.chanx_in_169_(sb_2__0__0_chanx_left_out_169_[0]),
		.chanx_in_170_(sb_1__0__0_chanx_right_out_170_[0]),
		.chanx_in_171_(sb_2__0__0_chanx_left_out_171_[0]),
		.chanx_in_172_(sb_1__0__0_chanx_right_out_172_[0]),
		.chanx_in_173_(sb_2__0__0_chanx_left_out_173_[0]),
		.chanx_in_174_(sb_1__0__0_chanx_right_out_174_[0]),
		.chanx_in_175_(sb_2__0__0_chanx_left_out_175_[0]),
		.chanx_in_176_(sb_1__0__0_chanx_right_out_176_[0]),
		.chanx_in_177_(sb_2__0__0_chanx_left_out_177_[0]),
		.chanx_in_178_(sb_1__0__0_chanx_right_out_178_[0]),
		.chanx_in_179_(sb_2__0__0_chanx_left_out_179_[0]),
		.chanx_in_180_(sb_1__0__0_chanx_right_out_180_[0]),
		.chanx_in_181_(sb_2__0__0_chanx_left_out_181_[0]),
		.chanx_in_182_(sb_1__0__0_chanx_right_out_182_[0]),
		.chanx_in_183_(sb_2__0__0_chanx_left_out_183_[0]),
		.chanx_in_184_(sb_1__0__0_chanx_right_out_184_[0]),
		.chanx_in_185_(sb_2__0__0_chanx_left_out_185_[0]),
		.chanx_in_186_(sb_1__0__0_chanx_right_out_186_[0]),
		.chanx_in_187_(sb_2__0__0_chanx_left_out_187_[0]),
		.chanx_in_188_(sb_1__0__0_chanx_right_out_188_[0]),
		.chanx_in_189_(sb_2__0__0_chanx_left_out_189_[0]),
		.chanx_in_190_(sb_1__0__0_chanx_right_out_190_[0]),
		.chanx_in_191_(sb_2__0__0_chanx_left_out_191_[0]),
		.chanx_in_192_(sb_1__0__0_chanx_right_out_192_[0]),
		.chanx_in_193_(sb_2__0__0_chanx_left_out_193_[0]),
		.chanx_in_194_(sb_1__0__0_chanx_right_out_194_[0]),
		.chanx_in_195_(sb_2__0__0_chanx_left_out_195_[0]),
		.chanx_in_196_(sb_1__0__0_chanx_right_out_196_[0]),
		.chanx_in_197_(sb_2__0__0_chanx_left_out_197_[0]),
		.chanx_in_198_(sb_1__0__0_chanx_right_out_198_[0]),
		.chanx_in_199_(sb_2__0__0_chanx_left_out_199_[0]),
		.ccff_head(sb_2__0__0_ccff_tail[0]),
		.chanx_out_0_(cbx_1__0__1_chanx_out_0_[0]),
		.chanx_out_1_(cbx_1__0__1_chanx_out_1_[0]),
		.chanx_out_2_(cbx_1__0__1_chanx_out_2_[0]),
		.chanx_out_3_(cbx_1__0__1_chanx_out_3_[0]),
		.chanx_out_4_(cbx_1__0__1_chanx_out_4_[0]),
		.chanx_out_5_(cbx_1__0__1_chanx_out_5_[0]),
		.chanx_out_6_(cbx_1__0__1_chanx_out_6_[0]),
		.chanx_out_7_(cbx_1__0__1_chanx_out_7_[0]),
		.chanx_out_8_(cbx_1__0__1_chanx_out_8_[0]),
		.chanx_out_9_(cbx_1__0__1_chanx_out_9_[0]),
		.chanx_out_10_(cbx_1__0__1_chanx_out_10_[0]),
		.chanx_out_11_(cbx_1__0__1_chanx_out_11_[0]),
		.chanx_out_12_(cbx_1__0__1_chanx_out_12_[0]),
		.chanx_out_13_(cbx_1__0__1_chanx_out_13_[0]),
		.chanx_out_14_(cbx_1__0__1_chanx_out_14_[0]),
		.chanx_out_15_(cbx_1__0__1_chanx_out_15_[0]),
		.chanx_out_16_(cbx_1__0__1_chanx_out_16_[0]),
		.chanx_out_17_(cbx_1__0__1_chanx_out_17_[0]),
		.chanx_out_18_(cbx_1__0__1_chanx_out_18_[0]),
		.chanx_out_19_(cbx_1__0__1_chanx_out_19_[0]),
		.chanx_out_20_(cbx_1__0__1_chanx_out_20_[0]),
		.chanx_out_21_(cbx_1__0__1_chanx_out_21_[0]),
		.chanx_out_22_(cbx_1__0__1_chanx_out_22_[0]),
		.chanx_out_23_(cbx_1__0__1_chanx_out_23_[0]),
		.chanx_out_24_(cbx_1__0__1_chanx_out_24_[0]),
		.chanx_out_25_(cbx_1__0__1_chanx_out_25_[0]),
		.chanx_out_26_(cbx_1__0__1_chanx_out_26_[0]),
		.chanx_out_27_(cbx_1__0__1_chanx_out_27_[0]),
		.chanx_out_28_(cbx_1__0__1_chanx_out_28_[0]),
		.chanx_out_29_(cbx_1__0__1_chanx_out_29_[0]),
		.chanx_out_30_(cbx_1__0__1_chanx_out_30_[0]),
		.chanx_out_31_(cbx_1__0__1_chanx_out_31_[0]),
		.chanx_out_32_(cbx_1__0__1_chanx_out_32_[0]),
		.chanx_out_33_(cbx_1__0__1_chanx_out_33_[0]),
		.chanx_out_34_(cbx_1__0__1_chanx_out_34_[0]),
		.chanx_out_35_(cbx_1__0__1_chanx_out_35_[0]),
		.chanx_out_36_(cbx_1__0__1_chanx_out_36_[0]),
		.chanx_out_37_(cbx_1__0__1_chanx_out_37_[0]),
		.chanx_out_38_(cbx_1__0__1_chanx_out_38_[0]),
		.chanx_out_39_(cbx_1__0__1_chanx_out_39_[0]),
		.chanx_out_40_(cbx_1__0__1_chanx_out_40_[0]),
		.chanx_out_41_(cbx_1__0__1_chanx_out_41_[0]),
		.chanx_out_42_(cbx_1__0__1_chanx_out_42_[0]),
		.chanx_out_43_(cbx_1__0__1_chanx_out_43_[0]),
		.chanx_out_44_(cbx_1__0__1_chanx_out_44_[0]),
		.chanx_out_45_(cbx_1__0__1_chanx_out_45_[0]),
		.chanx_out_46_(cbx_1__0__1_chanx_out_46_[0]),
		.chanx_out_47_(cbx_1__0__1_chanx_out_47_[0]),
		.chanx_out_48_(cbx_1__0__1_chanx_out_48_[0]),
		.chanx_out_49_(cbx_1__0__1_chanx_out_49_[0]),
		.chanx_out_50_(cbx_1__0__1_chanx_out_50_[0]),
		.chanx_out_51_(cbx_1__0__1_chanx_out_51_[0]),
		.chanx_out_52_(cbx_1__0__1_chanx_out_52_[0]),
		.chanx_out_53_(cbx_1__0__1_chanx_out_53_[0]),
		.chanx_out_54_(cbx_1__0__1_chanx_out_54_[0]),
		.chanx_out_55_(cbx_1__0__1_chanx_out_55_[0]),
		.chanx_out_56_(cbx_1__0__1_chanx_out_56_[0]),
		.chanx_out_57_(cbx_1__0__1_chanx_out_57_[0]),
		.chanx_out_58_(cbx_1__0__1_chanx_out_58_[0]),
		.chanx_out_59_(cbx_1__0__1_chanx_out_59_[0]),
		.chanx_out_60_(cbx_1__0__1_chanx_out_60_[0]),
		.chanx_out_61_(cbx_1__0__1_chanx_out_61_[0]),
		.chanx_out_62_(cbx_1__0__1_chanx_out_62_[0]),
		.chanx_out_63_(cbx_1__0__1_chanx_out_63_[0]),
		.chanx_out_64_(cbx_1__0__1_chanx_out_64_[0]),
		.chanx_out_65_(cbx_1__0__1_chanx_out_65_[0]),
		.chanx_out_66_(cbx_1__0__1_chanx_out_66_[0]),
		.chanx_out_67_(cbx_1__0__1_chanx_out_67_[0]),
		.chanx_out_68_(cbx_1__0__1_chanx_out_68_[0]),
		.chanx_out_69_(cbx_1__0__1_chanx_out_69_[0]),
		.chanx_out_70_(cbx_1__0__1_chanx_out_70_[0]),
		.chanx_out_71_(cbx_1__0__1_chanx_out_71_[0]),
		.chanx_out_72_(cbx_1__0__1_chanx_out_72_[0]),
		.chanx_out_73_(cbx_1__0__1_chanx_out_73_[0]),
		.chanx_out_74_(cbx_1__0__1_chanx_out_74_[0]),
		.chanx_out_75_(cbx_1__0__1_chanx_out_75_[0]),
		.chanx_out_76_(cbx_1__0__1_chanx_out_76_[0]),
		.chanx_out_77_(cbx_1__0__1_chanx_out_77_[0]),
		.chanx_out_78_(cbx_1__0__1_chanx_out_78_[0]),
		.chanx_out_79_(cbx_1__0__1_chanx_out_79_[0]),
		.chanx_out_80_(cbx_1__0__1_chanx_out_80_[0]),
		.chanx_out_81_(cbx_1__0__1_chanx_out_81_[0]),
		.chanx_out_82_(cbx_1__0__1_chanx_out_82_[0]),
		.chanx_out_83_(cbx_1__0__1_chanx_out_83_[0]),
		.chanx_out_84_(cbx_1__0__1_chanx_out_84_[0]),
		.chanx_out_85_(cbx_1__0__1_chanx_out_85_[0]),
		.chanx_out_86_(cbx_1__0__1_chanx_out_86_[0]),
		.chanx_out_87_(cbx_1__0__1_chanx_out_87_[0]),
		.chanx_out_88_(cbx_1__0__1_chanx_out_88_[0]),
		.chanx_out_89_(cbx_1__0__1_chanx_out_89_[0]),
		.chanx_out_90_(cbx_1__0__1_chanx_out_90_[0]),
		.chanx_out_91_(cbx_1__0__1_chanx_out_91_[0]),
		.chanx_out_92_(cbx_1__0__1_chanx_out_92_[0]),
		.chanx_out_93_(cbx_1__0__1_chanx_out_93_[0]),
		.chanx_out_94_(cbx_1__0__1_chanx_out_94_[0]),
		.chanx_out_95_(cbx_1__0__1_chanx_out_95_[0]),
		.chanx_out_96_(cbx_1__0__1_chanx_out_96_[0]),
		.chanx_out_97_(cbx_1__0__1_chanx_out_97_[0]),
		.chanx_out_98_(cbx_1__0__1_chanx_out_98_[0]),
		.chanx_out_99_(cbx_1__0__1_chanx_out_99_[0]),
		.chanx_out_100_(cbx_1__0__1_chanx_out_100_[0]),
		.chanx_out_101_(cbx_1__0__1_chanx_out_101_[0]),
		.chanx_out_102_(cbx_1__0__1_chanx_out_102_[0]),
		.chanx_out_103_(cbx_1__0__1_chanx_out_103_[0]),
		.chanx_out_104_(cbx_1__0__1_chanx_out_104_[0]),
		.chanx_out_105_(cbx_1__0__1_chanx_out_105_[0]),
		.chanx_out_106_(cbx_1__0__1_chanx_out_106_[0]),
		.chanx_out_107_(cbx_1__0__1_chanx_out_107_[0]),
		.chanx_out_108_(cbx_1__0__1_chanx_out_108_[0]),
		.chanx_out_109_(cbx_1__0__1_chanx_out_109_[0]),
		.chanx_out_110_(cbx_1__0__1_chanx_out_110_[0]),
		.chanx_out_111_(cbx_1__0__1_chanx_out_111_[0]),
		.chanx_out_112_(cbx_1__0__1_chanx_out_112_[0]),
		.chanx_out_113_(cbx_1__0__1_chanx_out_113_[0]),
		.chanx_out_114_(cbx_1__0__1_chanx_out_114_[0]),
		.chanx_out_115_(cbx_1__0__1_chanx_out_115_[0]),
		.chanx_out_116_(cbx_1__0__1_chanx_out_116_[0]),
		.chanx_out_117_(cbx_1__0__1_chanx_out_117_[0]),
		.chanx_out_118_(cbx_1__0__1_chanx_out_118_[0]),
		.chanx_out_119_(cbx_1__0__1_chanx_out_119_[0]),
		.chanx_out_120_(cbx_1__0__1_chanx_out_120_[0]),
		.chanx_out_121_(cbx_1__0__1_chanx_out_121_[0]),
		.chanx_out_122_(cbx_1__0__1_chanx_out_122_[0]),
		.chanx_out_123_(cbx_1__0__1_chanx_out_123_[0]),
		.chanx_out_124_(cbx_1__0__1_chanx_out_124_[0]),
		.chanx_out_125_(cbx_1__0__1_chanx_out_125_[0]),
		.chanx_out_126_(cbx_1__0__1_chanx_out_126_[0]),
		.chanx_out_127_(cbx_1__0__1_chanx_out_127_[0]),
		.chanx_out_128_(cbx_1__0__1_chanx_out_128_[0]),
		.chanx_out_129_(cbx_1__0__1_chanx_out_129_[0]),
		.chanx_out_130_(cbx_1__0__1_chanx_out_130_[0]),
		.chanx_out_131_(cbx_1__0__1_chanx_out_131_[0]),
		.chanx_out_132_(cbx_1__0__1_chanx_out_132_[0]),
		.chanx_out_133_(cbx_1__0__1_chanx_out_133_[0]),
		.chanx_out_134_(cbx_1__0__1_chanx_out_134_[0]),
		.chanx_out_135_(cbx_1__0__1_chanx_out_135_[0]),
		.chanx_out_136_(cbx_1__0__1_chanx_out_136_[0]),
		.chanx_out_137_(cbx_1__0__1_chanx_out_137_[0]),
		.chanx_out_138_(cbx_1__0__1_chanx_out_138_[0]),
		.chanx_out_139_(cbx_1__0__1_chanx_out_139_[0]),
		.chanx_out_140_(cbx_1__0__1_chanx_out_140_[0]),
		.chanx_out_141_(cbx_1__0__1_chanx_out_141_[0]),
		.chanx_out_142_(cbx_1__0__1_chanx_out_142_[0]),
		.chanx_out_143_(cbx_1__0__1_chanx_out_143_[0]),
		.chanx_out_144_(cbx_1__0__1_chanx_out_144_[0]),
		.chanx_out_145_(cbx_1__0__1_chanx_out_145_[0]),
		.chanx_out_146_(cbx_1__0__1_chanx_out_146_[0]),
		.chanx_out_147_(cbx_1__0__1_chanx_out_147_[0]),
		.chanx_out_148_(cbx_1__0__1_chanx_out_148_[0]),
		.chanx_out_149_(cbx_1__0__1_chanx_out_149_[0]),
		.chanx_out_150_(cbx_1__0__1_chanx_out_150_[0]),
		.chanx_out_151_(cbx_1__0__1_chanx_out_151_[0]),
		.chanx_out_152_(cbx_1__0__1_chanx_out_152_[0]),
		.chanx_out_153_(cbx_1__0__1_chanx_out_153_[0]),
		.chanx_out_154_(cbx_1__0__1_chanx_out_154_[0]),
		.chanx_out_155_(cbx_1__0__1_chanx_out_155_[0]),
		.chanx_out_156_(cbx_1__0__1_chanx_out_156_[0]),
		.chanx_out_157_(cbx_1__0__1_chanx_out_157_[0]),
		.chanx_out_158_(cbx_1__0__1_chanx_out_158_[0]),
		.chanx_out_159_(cbx_1__0__1_chanx_out_159_[0]),
		.chanx_out_160_(cbx_1__0__1_chanx_out_160_[0]),
		.chanx_out_161_(cbx_1__0__1_chanx_out_161_[0]),
		.chanx_out_162_(cbx_1__0__1_chanx_out_162_[0]),
		.chanx_out_163_(cbx_1__0__1_chanx_out_163_[0]),
		.chanx_out_164_(cbx_1__0__1_chanx_out_164_[0]),
		.chanx_out_165_(cbx_1__0__1_chanx_out_165_[0]),
		.chanx_out_166_(cbx_1__0__1_chanx_out_166_[0]),
		.chanx_out_167_(cbx_1__0__1_chanx_out_167_[0]),
		.chanx_out_168_(cbx_1__0__1_chanx_out_168_[0]),
		.chanx_out_169_(cbx_1__0__1_chanx_out_169_[0]),
		.chanx_out_170_(cbx_1__0__1_chanx_out_170_[0]),
		.chanx_out_171_(cbx_1__0__1_chanx_out_171_[0]),
		.chanx_out_172_(cbx_1__0__1_chanx_out_172_[0]),
		.chanx_out_173_(cbx_1__0__1_chanx_out_173_[0]),
		.chanx_out_174_(cbx_1__0__1_chanx_out_174_[0]),
		.chanx_out_175_(cbx_1__0__1_chanx_out_175_[0]),
		.chanx_out_176_(cbx_1__0__1_chanx_out_176_[0]),
		.chanx_out_177_(cbx_1__0__1_chanx_out_177_[0]),
		.chanx_out_178_(cbx_1__0__1_chanx_out_178_[0]),
		.chanx_out_179_(cbx_1__0__1_chanx_out_179_[0]),
		.chanx_out_180_(cbx_1__0__1_chanx_out_180_[0]),
		.chanx_out_181_(cbx_1__0__1_chanx_out_181_[0]),
		.chanx_out_182_(cbx_1__0__1_chanx_out_182_[0]),
		.chanx_out_183_(cbx_1__0__1_chanx_out_183_[0]),
		.chanx_out_184_(cbx_1__0__1_chanx_out_184_[0]),
		.chanx_out_185_(cbx_1__0__1_chanx_out_185_[0]),
		.chanx_out_186_(cbx_1__0__1_chanx_out_186_[0]),
		.chanx_out_187_(cbx_1__0__1_chanx_out_187_[0]),
		.chanx_out_188_(cbx_1__0__1_chanx_out_188_[0]),
		.chanx_out_189_(cbx_1__0__1_chanx_out_189_[0]),
		.chanx_out_190_(cbx_1__0__1_chanx_out_190_[0]),
		.chanx_out_191_(cbx_1__0__1_chanx_out_191_[0]),
		.chanx_out_192_(cbx_1__0__1_chanx_out_192_[0]),
		.chanx_out_193_(cbx_1__0__1_chanx_out_193_[0]),
		.chanx_out_194_(cbx_1__0__1_chanx_out_194_[0]),
		.chanx_out_195_(cbx_1__0__1_chanx_out_195_[0]),
		.chanx_out_196_(cbx_1__0__1_chanx_out_196_[0]),
		.chanx_out_197_(cbx_1__0__1_chanx_out_197_[0]),
		.chanx_out_198_(cbx_1__0__1_chanx_out_198_[0]),
		.chanx_out_199_(cbx_1__0__1_chanx_out_199_[0]),
		.top_grid_pin_20_(cbx_1__0__1_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__0__1_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__0__1_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__0__1_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__0__1_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__0__1_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__0__1_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__0__1_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__0__1_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__0__1_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__0__1_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__0__1_top_grid_pin_31_[0]),
		.top_grid_pin_32_(cbx_1__0__1_top_grid_pin_32_[0]),
		.top_grid_pin_33_(cbx_1__0__1_top_grid_pin_33_[0]),
		.top_grid_pin_34_(cbx_1__0__1_top_grid_pin_34_[0]),
		.top_grid_pin_35_(cbx_1__0__1_top_grid_pin_35_[0]),
		.top_grid_pin_36_(cbx_1__0__1_top_grid_pin_36_[0]),
		.top_grid_pin_37_(cbx_1__0__1_top_grid_pin_37_[0]),
		.top_grid_pin_38_(cbx_1__0__1_top_grid_pin_38_[0]),
		.top_grid_pin_39_(cbx_1__0__1_top_grid_pin_39_[0]),
		.bottom_grid_pin_0_(cbx_1__0__1_bottom_grid_pin_0_[0]),
		.ccff_tail(cbx_1__0__1_ccff_tail[0]));

	cbx_1__1_ cbx_1__1_ (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.chanx_in_0_(sb_0__1__0_chanx_right_out_0_[0]),
		.chanx_in_1_(sb_1__1__0_chanx_left_out_1_[0]),
		.chanx_in_2_(sb_0__1__0_chanx_right_out_2_[0]),
		.chanx_in_3_(sb_1__1__0_chanx_left_out_3_[0]),
		.chanx_in_4_(sb_0__1__0_chanx_right_out_4_[0]),
		.chanx_in_5_(sb_1__1__0_chanx_left_out_5_[0]),
		.chanx_in_6_(sb_0__1__0_chanx_right_out_6_[0]),
		.chanx_in_7_(sb_1__1__0_chanx_left_out_7_[0]),
		.chanx_in_8_(sb_0__1__0_chanx_right_out_8_[0]),
		.chanx_in_9_(sb_1__1__0_chanx_left_out_9_[0]),
		.chanx_in_10_(sb_0__1__0_chanx_right_out_10_[0]),
		.chanx_in_11_(sb_1__1__0_chanx_left_out_11_[0]),
		.chanx_in_12_(sb_0__1__0_chanx_right_out_12_[0]),
		.chanx_in_13_(sb_1__1__0_chanx_left_out_13_[0]),
		.chanx_in_14_(sb_0__1__0_chanx_right_out_14_[0]),
		.chanx_in_15_(sb_1__1__0_chanx_left_out_15_[0]),
		.chanx_in_16_(sb_0__1__0_chanx_right_out_16_[0]),
		.chanx_in_17_(sb_1__1__0_chanx_left_out_17_[0]),
		.chanx_in_18_(sb_0__1__0_chanx_right_out_18_[0]),
		.chanx_in_19_(sb_1__1__0_chanx_left_out_19_[0]),
		.chanx_in_20_(sb_0__1__0_chanx_right_out_20_[0]),
		.chanx_in_21_(sb_1__1__0_chanx_left_out_21_[0]),
		.chanx_in_22_(sb_0__1__0_chanx_right_out_22_[0]),
		.chanx_in_23_(sb_1__1__0_chanx_left_out_23_[0]),
		.chanx_in_24_(sb_0__1__0_chanx_right_out_24_[0]),
		.chanx_in_25_(sb_1__1__0_chanx_left_out_25_[0]),
		.chanx_in_26_(sb_0__1__0_chanx_right_out_26_[0]),
		.chanx_in_27_(sb_1__1__0_chanx_left_out_27_[0]),
		.chanx_in_28_(sb_0__1__0_chanx_right_out_28_[0]),
		.chanx_in_29_(sb_1__1__0_chanx_left_out_29_[0]),
		.chanx_in_30_(sb_0__1__0_chanx_right_out_30_[0]),
		.chanx_in_31_(sb_1__1__0_chanx_left_out_31_[0]),
		.chanx_in_32_(sb_0__1__0_chanx_right_out_32_[0]),
		.chanx_in_33_(sb_1__1__0_chanx_left_out_33_[0]),
		.chanx_in_34_(sb_0__1__0_chanx_right_out_34_[0]),
		.chanx_in_35_(sb_1__1__0_chanx_left_out_35_[0]),
		.chanx_in_36_(sb_0__1__0_chanx_right_out_36_[0]),
		.chanx_in_37_(sb_1__1__0_chanx_left_out_37_[0]),
		.chanx_in_38_(sb_0__1__0_chanx_right_out_38_[0]),
		.chanx_in_39_(sb_1__1__0_chanx_left_out_39_[0]),
		.chanx_in_40_(sb_0__1__0_chanx_right_out_40_[0]),
		.chanx_in_41_(sb_1__1__0_chanx_left_out_41_[0]),
		.chanx_in_42_(sb_0__1__0_chanx_right_out_42_[0]),
		.chanx_in_43_(sb_1__1__0_chanx_left_out_43_[0]),
		.chanx_in_44_(sb_0__1__0_chanx_right_out_44_[0]),
		.chanx_in_45_(sb_1__1__0_chanx_left_out_45_[0]),
		.chanx_in_46_(sb_0__1__0_chanx_right_out_46_[0]),
		.chanx_in_47_(sb_1__1__0_chanx_left_out_47_[0]),
		.chanx_in_48_(sb_0__1__0_chanx_right_out_48_[0]),
		.chanx_in_49_(sb_1__1__0_chanx_left_out_49_[0]),
		.chanx_in_50_(sb_0__1__0_chanx_right_out_50_[0]),
		.chanx_in_51_(sb_1__1__0_chanx_left_out_51_[0]),
		.chanx_in_52_(sb_0__1__0_chanx_right_out_52_[0]),
		.chanx_in_53_(sb_1__1__0_chanx_left_out_53_[0]),
		.chanx_in_54_(sb_0__1__0_chanx_right_out_54_[0]),
		.chanx_in_55_(sb_1__1__0_chanx_left_out_55_[0]),
		.chanx_in_56_(sb_0__1__0_chanx_right_out_56_[0]),
		.chanx_in_57_(sb_1__1__0_chanx_left_out_57_[0]),
		.chanx_in_58_(sb_0__1__0_chanx_right_out_58_[0]),
		.chanx_in_59_(sb_1__1__0_chanx_left_out_59_[0]),
		.chanx_in_60_(sb_0__1__0_chanx_right_out_60_[0]),
		.chanx_in_61_(sb_1__1__0_chanx_left_out_61_[0]),
		.chanx_in_62_(sb_0__1__0_chanx_right_out_62_[0]),
		.chanx_in_63_(sb_1__1__0_chanx_left_out_63_[0]),
		.chanx_in_64_(sb_0__1__0_chanx_right_out_64_[0]),
		.chanx_in_65_(sb_1__1__0_chanx_left_out_65_[0]),
		.chanx_in_66_(sb_0__1__0_chanx_right_out_66_[0]),
		.chanx_in_67_(sb_1__1__0_chanx_left_out_67_[0]),
		.chanx_in_68_(sb_0__1__0_chanx_right_out_68_[0]),
		.chanx_in_69_(sb_1__1__0_chanx_left_out_69_[0]),
		.chanx_in_70_(sb_0__1__0_chanx_right_out_70_[0]),
		.chanx_in_71_(sb_1__1__0_chanx_left_out_71_[0]),
		.chanx_in_72_(sb_0__1__0_chanx_right_out_72_[0]),
		.chanx_in_73_(sb_1__1__0_chanx_left_out_73_[0]),
		.chanx_in_74_(sb_0__1__0_chanx_right_out_74_[0]),
		.chanx_in_75_(sb_1__1__0_chanx_left_out_75_[0]),
		.chanx_in_76_(sb_0__1__0_chanx_right_out_76_[0]),
		.chanx_in_77_(sb_1__1__0_chanx_left_out_77_[0]),
		.chanx_in_78_(sb_0__1__0_chanx_right_out_78_[0]),
		.chanx_in_79_(sb_1__1__0_chanx_left_out_79_[0]),
		.chanx_in_80_(sb_0__1__0_chanx_right_out_80_[0]),
		.chanx_in_81_(sb_1__1__0_chanx_left_out_81_[0]),
		.chanx_in_82_(sb_0__1__0_chanx_right_out_82_[0]),
		.chanx_in_83_(sb_1__1__0_chanx_left_out_83_[0]),
		.chanx_in_84_(sb_0__1__0_chanx_right_out_84_[0]),
		.chanx_in_85_(sb_1__1__0_chanx_left_out_85_[0]),
		.chanx_in_86_(sb_0__1__0_chanx_right_out_86_[0]),
		.chanx_in_87_(sb_1__1__0_chanx_left_out_87_[0]),
		.chanx_in_88_(sb_0__1__0_chanx_right_out_88_[0]),
		.chanx_in_89_(sb_1__1__0_chanx_left_out_89_[0]),
		.chanx_in_90_(sb_0__1__0_chanx_right_out_90_[0]),
		.chanx_in_91_(sb_1__1__0_chanx_left_out_91_[0]),
		.chanx_in_92_(sb_0__1__0_chanx_right_out_92_[0]),
		.chanx_in_93_(sb_1__1__0_chanx_left_out_93_[0]),
		.chanx_in_94_(sb_0__1__0_chanx_right_out_94_[0]),
		.chanx_in_95_(sb_1__1__0_chanx_left_out_95_[0]),
		.chanx_in_96_(sb_0__1__0_chanx_right_out_96_[0]),
		.chanx_in_97_(sb_1__1__0_chanx_left_out_97_[0]),
		.chanx_in_98_(sb_0__1__0_chanx_right_out_98_[0]),
		.chanx_in_99_(sb_1__1__0_chanx_left_out_99_[0]),
		.chanx_in_100_(sb_0__1__0_chanx_right_out_100_[0]),
		.chanx_in_101_(sb_1__1__0_chanx_left_out_101_[0]),
		.chanx_in_102_(sb_0__1__0_chanx_right_out_102_[0]),
		.chanx_in_103_(sb_1__1__0_chanx_left_out_103_[0]),
		.chanx_in_104_(sb_0__1__0_chanx_right_out_104_[0]),
		.chanx_in_105_(sb_1__1__0_chanx_left_out_105_[0]),
		.chanx_in_106_(sb_0__1__0_chanx_right_out_106_[0]),
		.chanx_in_107_(sb_1__1__0_chanx_left_out_107_[0]),
		.chanx_in_108_(sb_0__1__0_chanx_right_out_108_[0]),
		.chanx_in_109_(sb_1__1__0_chanx_left_out_109_[0]),
		.chanx_in_110_(sb_0__1__0_chanx_right_out_110_[0]),
		.chanx_in_111_(sb_1__1__0_chanx_left_out_111_[0]),
		.chanx_in_112_(sb_0__1__0_chanx_right_out_112_[0]),
		.chanx_in_113_(sb_1__1__0_chanx_left_out_113_[0]),
		.chanx_in_114_(sb_0__1__0_chanx_right_out_114_[0]),
		.chanx_in_115_(sb_1__1__0_chanx_left_out_115_[0]),
		.chanx_in_116_(sb_0__1__0_chanx_right_out_116_[0]),
		.chanx_in_117_(sb_1__1__0_chanx_left_out_117_[0]),
		.chanx_in_118_(sb_0__1__0_chanx_right_out_118_[0]),
		.chanx_in_119_(sb_1__1__0_chanx_left_out_119_[0]),
		.chanx_in_120_(sb_0__1__0_chanx_right_out_120_[0]),
		.chanx_in_121_(sb_1__1__0_chanx_left_out_121_[0]),
		.chanx_in_122_(sb_0__1__0_chanx_right_out_122_[0]),
		.chanx_in_123_(sb_1__1__0_chanx_left_out_123_[0]),
		.chanx_in_124_(sb_0__1__0_chanx_right_out_124_[0]),
		.chanx_in_125_(sb_1__1__0_chanx_left_out_125_[0]),
		.chanx_in_126_(sb_0__1__0_chanx_right_out_126_[0]),
		.chanx_in_127_(sb_1__1__0_chanx_left_out_127_[0]),
		.chanx_in_128_(sb_0__1__0_chanx_right_out_128_[0]),
		.chanx_in_129_(sb_1__1__0_chanx_left_out_129_[0]),
		.chanx_in_130_(sb_0__1__0_chanx_right_out_130_[0]),
		.chanx_in_131_(sb_1__1__0_chanx_left_out_131_[0]),
		.chanx_in_132_(sb_0__1__0_chanx_right_out_132_[0]),
		.chanx_in_133_(sb_1__1__0_chanx_left_out_133_[0]),
		.chanx_in_134_(sb_0__1__0_chanx_right_out_134_[0]),
		.chanx_in_135_(sb_1__1__0_chanx_left_out_135_[0]),
		.chanx_in_136_(sb_0__1__0_chanx_right_out_136_[0]),
		.chanx_in_137_(sb_1__1__0_chanx_left_out_137_[0]),
		.chanx_in_138_(sb_0__1__0_chanx_right_out_138_[0]),
		.chanx_in_139_(sb_1__1__0_chanx_left_out_139_[0]),
		.chanx_in_140_(sb_0__1__0_chanx_right_out_140_[0]),
		.chanx_in_141_(sb_1__1__0_chanx_left_out_141_[0]),
		.chanx_in_142_(sb_0__1__0_chanx_right_out_142_[0]),
		.chanx_in_143_(sb_1__1__0_chanx_left_out_143_[0]),
		.chanx_in_144_(sb_0__1__0_chanx_right_out_144_[0]),
		.chanx_in_145_(sb_1__1__0_chanx_left_out_145_[0]),
		.chanx_in_146_(sb_0__1__0_chanx_right_out_146_[0]),
		.chanx_in_147_(sb_1__1__0_chanx_left_out_147_[0]),
		.chanx_in_148_(sb_0__1__0_chanx_right_out_148_[0]),
		.chanx_in_149_(sb_1__1__0_chanx_left_out_149_[0]),
		.chanx_in_150_(sb_0__1__0_chanx_right_out_150_[0]),
		.chanx_in_151_(sb_1__1__0_chanx_left_out_151_[0]),
		.chanx_in_152_(sb_0__1__0_chanx_right_out_152_[0]),
		.chanx_in_153_(sb_1__1__0_chanx_left_out_153_[0]),
		.chanx_in_154_(sb_0__1__0_chanx_right_out_154_[0]),
		.chanx_in_155_(sb_1__1__0_chanx_left_out_155_[0]),
		.chanx_in_156_(sb_0__1__0_chanx_right_out_156_[0]),
		.chanx_in_157_(sb_1__1__0_chanx_left_out_157_[0]),
		.chanx_in_158_(sb_0__1__0_chanx_right_out_158_[0]),
		.chanx_in_159_(sb_1__1__0_chanx_left_out_159_[0]),
		.chanx_in_160_(sb_0__1__0_chanx_right_out_160_[0]),
		.chanx_in_161_(sb_1__1__0_chanx_left_out_161_[0]),
		.chanx_in_162_(sb_0__1__0_chanx_right_out_162_[0]),
		.chanx_in_163_(sb_1__1__0_chanx_left_out_163_[0]),
		.chanx_in_164_(sb_0__1__0_chanx_right_out_164_[0]),
		.chanx_in_165_(sb_1__1__0_chanx_left_out_165_[0]),
		.chanx_in_166_(sb_0__1__0_chanx_right_out_166_[0]),
		.chanx_in_167_(sb_1__1__0_chanx_left_out_167_[0]),
		.chanx_in_168_(sb_0__1__0_chanx_right_out_168_[0]),
		.chanx_in_169_(sb_1__1__0_chanx_left_out_169_[0]),
		.chanx_in_170_(sb_0__1__0_chanx_right_out_170_[0]),
		.chanx_in_171_(sb_1__1__0_chanx_left_out_171_[0]),
		.chanx_in_172_(sb_0__1__0_chanx_right_out_172_[0]),
		.chanx_in_173_(sb_1__1__0_chanx_left_out_173_[0]),
		.chanx_in_174_(sb_0__1__0_chanx_right_out_174_[0]),
		.chanx_in_175_(sb_1__1__0_chanx_left_out_175_[0]),
		.chanx_in_176_(sb_0__1__0_chanx_right_out_176_[0]),
		.chanx_in_177_(sb_1__1__0_chanx_left_out_177_[0]),
		.chanx_in_178_(sb_0__1__0_chanx_right_out_178_[0]),
		.chanx_in_179_(sb_1__1__0_chanx_left_out_179_[0]),
		.chanx_in_180_(sb_0__1__0_chanx_right_out_180_[0]),
		.chanx_in_181_(sb_1__1__0_chanx_left_out_181_[0]),
		.chanx_in_182_(sb_0__1__0_chanx_right_out_182_[0]),
		.chanx_in_183_(sb_1__1__0_chanx_left_out_183_[0]),
		.chanx_in_184_(sb_0__1__0_chanx_right_out_184_[0]),
		.chanx_in_185_(sb_1__1__0_chanx_left_out_185_[0]),
		.chanx_in_186_(sb_0__1__0_chanx_right_out_186_[0]),
		.chanx_in_187_(sb_1__1__0_chanx_left_out_187_[0]),
		.chanx_in_188_(sb_0__1__0_chanx_right_out_188_[0]),
		.chanx_in_189_(sb_1__1__0_chanx_left_out_189_[0]),
		.chanx_in_190_(sb_0__1__0_chanx_right_out_190_[0]),
		.chanx_in_191_(sb_1__1__0_chanx_left_out_191_[0]),
		.chanx_in_192_(sb_0__1__0_chanx_right_out_192_[0]),
		.chanx_in_193_(sb_1__1__0_chanx_left_out_193_[0]),
		.chanx_in_194_(sb_0__1__0_chanx_right_out_194_[0]),
		.chanx_in_195_(sb_1__1__0_chanx_left_out_195_[0]),
		.chanx_in_196_(sb_0__1__0_chanx_right_out_196_[0]),
		.chanx_in_197_(sb_1__1__0_chanx_left_out_197_[0]),
		.chanx_in_198_(sb_0__1__0_chanx_right_out_198_[0]),
		.chanx_in_199_(sb_1__1__0_chanx_left_out_199_[0]),
		.ccff_head(sb_1__1__0_ccff_tail[0]),
		.chanx_out_0_(cbx_1__1__0_chanx_out_0_[0]),
		.chanx_out_1_(cbx_1__1__0_chanx_out_1_[0]),
		.chanx_out_2_(cbx_1__1__0_chanx_out_2_[0]),
		.chanx_out_3_(cbx_1__1__0_chanx_out_3_[0]),
		.chanx_out_4_(cbx_1__1__0_chanx_out_4_[0]),
		.chanx_out_5_(cbx_1__1__0_chanx_out_5_[0]),
		.chanx_out_6_(cbx_1__1__0_chanx_out_6_[0]),
		.chanx_out_7_(cbx_1__1__0_chanx_out_7_[0]),
		.chanx_out_8_(cbx_1__1__0_chanx_out_8_[0]),
		.chanx_out_9_(cbx_1__1__0_chanx_out_9_[0]),
		.chanx_out_10_(cbx_1__1__0_chanx_out_10_[0]),
		.chanx_out_11_(cbx_1__1__0_chanx_out_11_[0]),
		.chanx_out_12_(cbx_1__1__0_chanx_out_12_[0]),
		.chanx_out_13_(cbx_1__1__0_chanx_out_13_[0]),
		.chanx_out_14_(cbx_1__1__0_chanx_out_14_[0]),
		.chanx_out_15_(cbx_1__1__0_chanx_out_15_[0]),
		.chanx_out_16_(cbx_1__1__0_chanx_out_16_[0]),
		.chanx_out_17_(cbx_1__1__0_chanx_out_17_[0]),
		.chanx_out_18_(cbx_1__1__0_chanx_out_18_[0]),
		.chanx_out_19_(cbx_1__1__0_chanx_out_19_[0]),
		.chanx_out_20_(cbx_1__1__0_chanx_out_20_[0]),
		.chanx_out_21_(cbx_1__1__0_chanx_out_21_[0]),
		.chanx_out_22_(cbx_1__1__0_chanx_out_22_[0]),
		.chanx_out_23_(cbx_1__1__0_chanx_out_23_[0]),
		.chanx_out_24_(cbx_1__1__0_chanx_out_24_[0]),
		.chanx_out_25_(cbx_1__1__0_chanx_out_25_[0]),
		.chanx_out_26_(cbx_1__1__0_chanx_out_26_[0]),
		.chanx_out_27_(cbx_1__1__0_chanx_out_27_[0]),
		.chanx_out_28_(cbx_1__1__0_chanx_out_28_[0]),
		.chanx_out_29_(cbx_1__1__0_chanx_out_29_[0]),
		.chanx_out_30_(cbx_1__1__0_chanx_out_30_[0]),
		.chanx_out_31_(cbx_1__1__0_chanx_out_31_[0]),
		.chanx_out_32_(cbx_1__1__0_chanx_out_32_[0]),
		.chanx_out_33_(cbx_1__1__0_chanx_out_33_[0]),
		.chanx_out_34_(cbx_1__1__0_chanx_out_34_[0]),
		.chanx_out_35_(cbx_1__1__0_chanx_out_35_[0]),
		.chanx_out_36_(cbx_1__1__0_chanx_out_36_[0]),
		.chanx_out_37_(cbx_1__1__0_chanx_out_37_[0]),
		.chanx_out_38_(cbx_1__1__0_chanx_out_38_[0]),
		.chanx_out_39_(cbx_1__1__0_chanx_out_39_[0]),
		.chanx_out_40_(cbx_1__1__0_chanx_out_40_[0]),
		.chanx_out_41_(cbx_1__1__0_chanx_out_41_[0]),
		.chanx_out_42_(cbx_1__1__0_chanx_out_42_[0]),
		.chanx_out_43_(cbx_1__1__0_chanx_out_43_[0]),
		.chanx_out_44_(cbx_1__1__0_chanx_out_44_[0]),
		.chanx_out_45_(cbx_1__1__0_chanx_out_45_[0]),
		.chanx_out_46_(cbx_1__1__0_chanx_out_46_[0]),
		.chanx_out_47_(cbx_1__1__0_chanx_out_47_[0]),
		.chanx_out_48_(cbx_1__1__0_chanx_out_48_[0]),
		.chanx_out_49_(cbx_1__1__0_chanx_out_49_[0]),
		.chanx_out_50_(cbx_1__1__0_chanx_out_50_[0]),
		.chanx_out_51_(cbx_1__1__0_chanx_out_51_[0]),
		.chanx_out_52_(cbx_1__1__0_chanx_out_52_[0]),
		.chanx_out_53_(cbx_1__1__0_chanx_out_53_[0]),
		.chanx_out_54_(cbx_1__1__0_chanx_out_54_[0]),
		.chanx_out_55_(cbx_1__1__0_chanx_out_55_[0]),
		.chanx_out_56_(cbx_1__1__0_chanx_out_56_[0]),
		.chanx_out_57_(cbx_1__1__0_chanx_out_57_[0]),
		.chanx_out_58_(cbx_1__1__0_chanx_out_58_[0]),
		.chanx_out_59_(cbx_1__1__0_chanx_out_59_[0]),
		.chanx_out_60_(cbx_1__1__0_chanx_out_60_[0]),
		.chanx_out_61_(cbx_1__1__0_chanx_out_61_[0]),
		.chanx_out_62_(cbx_1__1__0_chanx_out_62_[0]),
		.chanx_out_63_(cbx_1__1__0_chanx_out_63_[0]),
		.chanx_out_64_(cbx_1__1__0_chanx_out_64_[0]),
		.chanx_out_65_(cbx_1__1__0_chanx_out_65_[0]),
		.chanx_out_66_(cbx_1__1__0_chanx_out_66_[0]),
		.chanx_out_67_(cbx_1__1__0_chanx_out_67_[0]),
		.chanx_out_68_(cbx_1__1__0_chanx_out_68_[0]),
		.chanx_out_69_(cbx_1__1__0_chanx_out_69_[0]),
		.chanx_out_70_(cbx_1__1__0_chanx_out_70_[0]),
		.chanx_out_71_(cbx_1__1__0_chanx_out_71_[0]),
		.chanx_out_72_(cbx_1__1__0_chanx_out_72_[0]),
		.chanx_out_73_(cbx_1__1__0_chanx_out_73_[0]),
		.chanx_out_74_(cbx_1__1__0_chanx_out_74_[0]),
		.chanx_out_75_(cbx_1__1__0_chanx_out_75_[0]),
		.chanx_out_76_(cbx_1__1__0_chanx_out_76_[0]),
		.chanx_out_77_(cbx_1__1__0_chanx_out_77_[0]),
		.chanx_out_78_(cbx_1__1__0_chanx_out_78_[0]),
		.chanx_out_79_(cbx_1__1__0_chanx_out_79_[0]),
		.chanx_out_80_(cbx_1__1__0_chanx_out_80_[0]),
		.chanx_out_81_(cbx_1__1__0_chanx_out_81_[0]),
		.chanx_out_82_(cbx_1__1__0_chanx_out_82_[0]),
		.chanx_out_83_(cbx_1__1__0_chanx_out_83_[0]),
		.chanx_out_84_(cbx_1__1__0_chanx_out_84_[0]),
		.chanx_out_85_(cbx_1__1__0_chanx_out_85_[0]),
		.chanx_out_86_(cbx_1__1__0_chanx_out_86_[0]),
		.chanx_out_87_(cbx_1__1__0_chanx_out_87_[0]),
		.chanx_out_88_(cbx_1__1__0_chanx_out_88_[0]),
		.chanx_out_89_(cbx_1__1__0_chanx_out_89_[0]),
		.chanx_out_90_(cbx_1__1__0_chanx_out_90_[0]),
		.chanx_out_91_(cbx_1__1__0_chanx_out_91_[0]),
		.chanx_out_92_(cbx_1__1__0_chanx_out_92_[0]),
		.chanx_out_93_(cbx_1__1__0_chanx_out_93_[0]),
		.chanx_out_94_(cbx_1__1__0_chanx_out_94_[0]),
		.chanx_out_95_(cbx_1__1__0_chanx_out_95_[0]),
		.chanx_out_96_(cbx_1__1__0_chanx_out_96_[0]),
		.chanx_out_97_(cbx_1__1__0_chanx_out_97_[0]),
		.chanx_out_98_(cbx_1__1__0_chanx_out_98_[0]),
		.chanx_out_99_(cbx_1__1__0_chanx_out_99_[0]),
		.chanx_out_100_(cbx_1__1__0_chanx_out_100_[0]),
		.chanx_out_101_(cbx_1__1__0_chanx_out_101_[0]),
		.chanx_out_102_(cbx_1__1__0_chanx_out_102_[0]),
		.chanx_out_103_(cbx_1__1__0_chanx_out_103_[0]),
		.chanx_out_104_(cbx_1__1__0_chanx_out_104_[0]),
		.chanx_out_105_(cbx_1__1__0_chanx_out_105_[0]),
		.chanx_out_106_(cbx_1__1__0_chanx_out_106_[0]),
		.chanx_out_107_(cbx_1__1__0_chanx_out_107_[0]),
		.chanx_out_108_(cbx_1__1__0_chanx_out_108_[0]),
		.chanx_out_109_(cbx_1__1__0_chanx_out_109_[0]),
		.chanx_out_110_(cbx_1__1__0_chanx_out_110_[0]),
		.chanx_out_111_(cbx_1__1__0_chanx_out_111_[0]),
		.chanx_out_112_(cbx_1__1__0_chanx_out_112_[0]),
		.chanx_out_113_(cbx_1__1__0_chanx_out_113_[0]),
		.chanx_out_114_(cbx_1__1__0_chanx_out_114_[0]),
		.chanx_out_115_(cbx_1__1__0_chanx_out_115_[0]),
		.chanx_out_116_(cbx_1__1__0_chanx_out_116_[0]),
		.chanx_out_117_(cbx_1__1__0_chanx_out_117_[0]),
		.chanx_out_118_(cbx_1__1__0_chanx_out_118_[0]),
		.chanx_out_119_(cbx_1__1__0_chanx_out_119_[0]),
		.chanx_out_120_(cbx_1__1__0_chanx_out_120_[0]),
		.chanx_out_121_(cbx_1__1__0_chanx_out_121_[0]),
		.chanx_out_122_(cbx_1__1__0_chanx_out_122_[0]),
		.chanx_out_123_(cbx_1__1__0_chanx_out_123_[0]),
		.chanx_out_124_(cbx_1__1__0_chanx_out_124_[0]),
		.chanx_out_125_(cbx_1__1__0_chanx_out_125_[0]),
		.chanx_out_126_(cbx_1__1__0_chanx_out_126_[0]),
		.chanx_out_127_(cbx_1__1__0_chanx_out_127_[0]),
		.chanx_out_128_(cbx_1__1__0_chanx_out_128_[0]),
		.chanx_out_129_(cbx_1__1__0_chanx_out_129_[0]),
		.chanx_out_130_(cbx_1__1__0_chanx_out_130_[0]),
		.chanx_out_131_(cbx_1__1__0_chanx_out_131_[0]),
		.chanx_out_132_(cbx_1__1__0_chanx_out_132_[0]),
		.chanx_out_133_(cbx_1__1__0_chanx_out_133_[0]),
		.chanx_out_134_(cbx_1__1__0_chanx_out_134_[0]),
		.chanx_out_135_(cbx_1__1__0_chanx_out_135_[0]),
		.chanx_out_136_(cbx_1__1__0_chanx_out_136_[0]),
		.chanx_out_137_(cbx_1__1__0_chanx_out_137_[0]),
		.chanx_out_138_(cbx_1__1__0_chanx_out_138_[0]),
		.chanx_out_139_(cbx_1__1__0_chanx_out_139_[0]),
		.chanx_out_140_(cbx_1__1__0_chanx_out_140_[0]),
		.chanx_out_141_(cbx_1__1__0_chanx_out_141_[0]),
		.chanx_out_142_(cbx_1__1__0_chanx_out_142_[0]),
		.chanx_out_143_(cbx_1__1__0_chanx_out_143_[0]),
		.chanx_out_144_(cbx_1__1__0_chanx_out_144_[0]),
		.chanx_out_145_(cbx_1__1__0_chanx_out_145_[0]),
		.chanx_out_146_(cbx_1__1__0_chanx_out_146_[0]),
		.chanx_out_147_(cbx_1__1__0_chanx_out_147_[0]),
		.chanx_out_148_(cbx_1__1__0_chanx_out_148_[0]),
		.chanx_out_149_(cbx_1__1__0_chanx_out_149_[0]),
		.chanx_out_150_(cbx_1__1__0_chanx_out_150_[0]),
		.chanx_out_151_(cbx_1__1__0_chanx_out_151_[0]),
		.chanx_out_152_(cbx_1__1__0_chanx_out_152_[0]),
		.chanx_out_153_(cbx_1__1__0_chanx_out_153_[0]),
		.chanx_out_154_(cbx_1__1__0_chanx_out_154_[0]),
		.chanx_out_155_(cbx_1__1__0_chanx_out_155_[0]),
		.chanx_out_156_(cbx_1__1__0_chanx_out_156_[0]),
		.chanx_out_157_(cbx_1__1__0_chanx_out_157_[0]),
		.chanx_out_158_(cbx_1__1__0_chanx_out_158_[0]),
		.chanx_out_159_(cbx_1__1__0_chanx_out_159_[0]),
		.chanx_out_160_(cbx_1__1__0_chanx_out_160_[0]),
		.chanx_out_161_(cbx_1__1__0_chanx_out_161_[0]),
		.chanx_out_162_(cbx_1__1__0_chanx_out_162_[0]),
		.chanx_out_163_(cbx_1__1__0_chanx_out_163_[0]),
		.chanx_out_164_(cbx_1__1__0_chanx_out_164_[0]),
		.chanx_out_165_(cbx_1__1__0_chanx_out_165_[0]),
		.chanx_out_166_(cbx_1__1__0_chanx_out_166_[0]),
		.chanx_out_167_(cbx_1__1__0_chanx_out_167_[0]),
		.chanx_out_168_(cbx_1__1__0_chanx_out_168_[0]),
		.chanx_out_169_(cbx_1__1__0_chanx_out_169_[0]),
		.chanx_out_170_(cbx_1__1__0_chanx_out_170_[0]),
		.chanx_out_171_(cbx_1__1__0_chanx_out_171_[0]),
		.chanx_out_172_(cbx_1__1__0_chanx_out_172_[0]),
		.chanx_out_173_(cbx_1__1__0_chanx_out_173_[0]),
		.chanx_out_174_(cbx_1__1__0_chanx_out_174_[0]),
		.chanx_out_175_(cbx_1__1__0_chanx_out_175_[0]),
		.chanx_out_176_(cbx_1__1__0_chanx_out_176_[0]),
		.chanx_out_177_(cbx_1__1__0_chanx_out_177_[0]),
		.chanx_out_178_(cbx_1__1__0_chanx_out_178_[0]),
		.chanx_out_179_(cbx_1__1__0_chanx_out_179_[0]),
		.chanx_out_180_(cbx_1__1__0_chanx_out_180_[0]),
		.chanx_out_181_(cbx_1__1__0_chanx_out_181_[0]),
		.chanx_out_182_(cbx_1__1__0_chanx_out_182_[0]),
		.chanx_out_183_(cbx_1__1__0_chanx_out_183_[0]),
		.chanx_out_184_(cbx_1__1__0_chanx_out_184_[0]),
		.chanx_out_185_(cbx_1__1__0_chanx_out_185_[0]),
		.chanx_out_186_(cbx_1__1__0_chanx_out_186_[0]),
		.chanx_out_187_(cbx_1__1__0_chanx_out_187_[0]),
		.chanx_out_188_(cbx_1__1__0_chanx_out_188_[0]),
		.chanx_out_189_(cbx_1__1__0_chanx_out_189_[0]),
		.chanx_out_190_(cbx_1__1__0_chanx_out_190_[0]),
		.chanx_out_191_(cbx_1__1__0_chanx_out_191_[0]),
		.chanx_out_192_(cbx_1__1__0_chanx_out_192_[0]),
		.chanx_out_193_(cbx_1__1__0_chanx_out_193_[0]),
		.chanx_out_194_(cbx_1__1__0_chanx_out_194_[0]),
		.chanx_out_195_(cbx_1__1__0_chanx_out_195_[0]),
		.chanx_out_196_(cbx_1__1__0_chanx_out_196_[0]),
		.chanx_out_197_(cbx_1__1__0_chanx_out_197_[0]),
		.chanx_out_198_(cbx_1__1__0_chanx_out_198_[0]),
		.chanx_out_199_(cbx_1__1__0_chanx_out_199_[0]),
		.top_grid_pin_20_(cbx_1__1__0_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__0_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__0_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__0_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__0_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__0_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__0_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__0_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__0_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__0_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__0_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__0_top_grid_pin_31_[0]),
		.top_grid_pin_32_(cbx_1__1__0_top_grid_pin_32_[0]),
		.top_grid_pin_33_(cbx_1__1__0_top_grid_pin_33_[0]),
		.top_grid_pin_34_(cbx_1__1__0_top_grid_pin_34_[0]),
		.top_grid_pin_35_(cbx_1__1__0_top_grid_pin_35_[0]),
		.top_grid_pin_36_(cbx_1__1__0_top_grid_pin_36_[0]),
		.top_grid_pin_37_(cbx_1__1__0_top_grid_pin_37_[0]),
		.top_grid_pin_38_(cbx_1__1__0_top_grid_pin_38_[0]),
		.top_grid_pin_39_(cbx_1__1__0_top_grid_pin_39_[0]),
		.bottom_grid_pin_42_(cbx_1__1__0_bottom_grid_pin_42_[0]),
		.bottom_grid_pin_43_(cbx_1__1__0_bottom_grid_pin_43_[0]),
		.bottom_grid_pin_69_(cbx_1__1__0_bottom_grid_pin_69_[0]),
		.ccff_tail(cbx_1__1__0_ccff_tail[0]));

	cbx_1__1_ cbx_2__1_ (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.chanx_in_0_(sb_1__1__0_chanx_right_out_0_[0]),
		.chanx_in_1_(sb_2__1__0_chanx_left_out_1_[0]),
		.chanx_in_2_(sb_1__1__0_chanx_right_out_2_[0]),
		.chanx_in_3_(sb_2__1__0_chanx_left_out_3_[0]),
		.chanx_in_4_(sb_1__1__0_chanx_right_out_4_[0]),
		.chanx_in_5_(sb_2__1__0_chanx_left_out_5_[0]),
		.chanx_in_6_(sb_1__1__0_chanx_right_out_6_[0]),
		.chanx_in_7_(sb_2__1__0_chanx_left_out_7_[0]),
		.chanx_in_8_(sb_1__1__0_chanx_right_out_8_[0]),
		.chanx_in_9_(sb_2__1__0_chanx_left_out_9_[0]),
		.chanx_in_10_(sb_1__1__0_chanx_right_out_10_[0]),
		.chanx_in_11_(sb_2__1__0_chanx_left_out_11_[0]),
		.chanx_in_12_(sb_1__1__0_chanx_right_out_12_[0]),
		.chanx_in_13_(sb_2__1__0_chanx_left_out_13_[0]),
		.chanx_in_14_(sb_1__1__0_chanx_right_out_14_[0]),
		.chanx_in_15_(sb_2__1__0_chanx_left_out_15_[0]),
		.chanx_in_16_(sb_1__1__0_chanx_right_out_16_[0]),
		.chanx_in_17_(sb_2__1__0_chanx_left_out_17_[0]),
		.chanx_in_18_(sb_1__1__0_chanx_right_out_18_[0]),
		.chanx_in_19_(sb_2__1__0_chanx_left_out_19_[0]),
		.chanx_in_20_(sb_1__1__0_chanx_right_out_20_[0]),
		.chanx_in_21_(sb_2__1__0_chanx_left_out_21_[0]),
		.chanx_in_22_(sb_1__1__0_chanx_right_out_22_[0]),
		.chanx_in_23_(sb_2__1__0_chanx_left_out_23_[0]),
		.chanx_in_24_(sb_1__1__0_chanx_right_out_24_[0]),
		.chanx_in_25_(sb_2__1__0_chanx_left_out_25_[0]),
		.chanx_in_26_(sb_1__1__0_chanx_right_out_26_[0]),
		.chanx_in_27_(sb_2__1__0_chanx_left_out_27_[0]),
		.chanx_in_28_(sb_1__1__0_chanx_right_out_28_[0]),
		.chanx_in_29_(sb_2__1__0_chanx_left_out_29_[0]),
		.chanx_in_30_(sb_1__1__0_chanx_right_out_30_[0]),
		.chanx_in_31_(sb_2__1__0_chanx_left_out_31_[0]),
		.chanx_in_32_(sb_1__1__0_chanx_right_out_32_[0]),
		.chanx_in_33_(sb_2__1__0_chanx_left_out_33_[0]),
		.chanx_in_34_(sb_1__1__0_chanx_right_out_34_[0]),
		.chanx_in_35_(sb_2__1__0_chanx_left_out_35_[0]),
		.chanx_in_36_(sb_1__1__0_chanx_right_out_36_[0]),
		.chanx_in_37_(sb_2__1__0_chanx_left_out_37_[0]),
		.chanx_in_38_(sb_1__1__0_chanx_right_out_38_[0]),
		.chanx_in_39_(sb_2__1__0_chanx_left_out_39_[0]),
		.chanx_in_40_(sb_1__1__0_chanx_right_out_40_[0]),
		.chanx_in_41_(sb_2__1__0_chanx_left_out_41_[0]),
		.chanx_in_42_(sb_1__1__0_chanx_right_out_42_[0]),
		.chanx_in_43_(sb_2__1__0_chanx_left_out_43_[0]),
		.chanx_in_44_(sb_1__1__0_chanx_right_out_44_[0]),
		.chanx_in_45_(sb_2__1__0_chanx_left_out_45_[0]),
		.chanx_in_46_(sb_1__1__0_chanx_right_out_46_[0]),
		.chanx_in_47_(sb_2__1__0_chanx_left_out_47_[0]),
		.chanx_in_48_(sb_1__1__0_chanx_right_out_48_[0]),
		.chanx_in_49_(sb_2__1__0_chanx_left_out_49_[0]),
		.chanx_in_50_(sb_1__1__0_chanx_right_out_50_[0]),
		.chanx_in_51_(sb_2__1__0_chanx_left_out_51_[0]),
		.chanx_in_52_(sb_1__1__0_chanx_right_out_52_[0]),
		.chanx_in_53_(sb_2__1__0_chanx_left_out_53_[0]),
		.chanx_in_54_(sb_1__1__0_chanx_right_out_54_[0]),
		.chanx_in_55_(sb_2__1__0_chanx_left_out_55_[0]),
		.chanx_in_56_(sb_1__1__0_chanx_right_out_56_[0]),
		.chanx_in_57_(sb_2__1__0_chanx_left_out_57_[0]),
		.chanx_in_58_(sb_1__1__0_chanx_right_out_58_[0]),
		.chanx_in_59_(sb_2__1__0_chanx_left_out_59_[0]),
		.chanx_in_60_(sb_1__1__0_chanx_right_out_60_[0]),
		.chanx_in_61_(sb_2__1__0_chanx_left_out_61_[0]),
		.chanx_in_62_(sb_1__1__0_chanx_right_out_62_[0]),
		.chanx_in_63_(sb_2__1__0_chanx_left_out_63_[0]),
		.chanx_in_64_(sb_1__1__0_chanx_right_out_64_[0]),
		.chanx_in_65_(sb_2__1__0_chanx_left_out_65_[0]),
		.chanx_in_66_(sb_1__1__0_chanx_right_out_66_[0]),
		.chanx_in_67_(sb_2__1__0_chanx_left_out_67_[0]),
		.chanx_in_68_(sb_1__1__0_chanx_right_out_68_[0]),
		.chanx_in_69_(sb_2__1__0_chanx_left_out_69_[0]),
		.chanx_in_70_(sb_1__1__0_chanx_right_out_70_[0]),
		.chanx_in_71_(sb_2__1__0_chanx_left_out_71_[0]),
		.chanx_in_72_(sb_1__1__0_chanx_right_out_72_[0]),
		.chanx_in_73_(sb_2__1__0_chanx_left_out_73_[0]),
		.chanx_in_74_(sb_1__1__0_chanx_right_out_74_[0]),
		.chanx_in_75_(sb_2__1__0_chanx_left_out_75_[0]),
		.chanx_in_76_(sb_1__1__0_chanx_right_out_76_[0]),
		.chanx_in_77_(sb_2__1__0_chanx_left_out_77_[0]),
		.chanx_in_78_(sb_1__1__0_chanx_right_out_78_[0]),
		.chanx_in_79_(sb_2__1__0_chanx_left_out_79_[0]),
		.chanx_in_80_(sb_1__1__0_chanx_right_out_80_[0]),
		.chanx_in_81_(sb_2__1__0_chanx_left_out_81_[0]),
		.chanx_in_82_(sb_1__1__0_chanx_right_out_82_[0]),
		.chanx_in_83_(sb_2__1__0_chanx_left_out_83_[0]),
		.chanx_in_84_(sb_1__1__0_chanx_right_out_84_[0]),
		.chanx_in_85_(sb_2__1__0_chanx_left_out_85_[0]),
		.chanx_in_86_(sb_1__1__0_chanx_right_out_86_[0]),
		.chanx_in_87_(sb_2__1__0_chanx_left_out_87_[0]),
		.chanx_in_88_(sb_1__1__0_chanx_right_out_88_[0]),
		.chanx_in_89_(sb_2__1__0_chanx_left_out_89_[0]),
		.chanx_in_90_(sb_1__1__0_chanx_right_out_90_[0]),
		.chanx_in_91_(sb_2__1__0_chanx_left_out_91_[0]),
		.chanx_in_92_(sb_1__1__0_chanx_right_out_92_[0]),
		.chanx_in_93_(sb_2__1__0_chanx_left_out_93_[0]),
		.chanx_in_94_(sb_1__1__0_chanx_right_out_94_[0]),
		.chanx_in_95_(sb_2__1__0_chanx_left_out_95_[0]),
		.chanx_in_96_(sb_1__1__0_chanx_right_out_96_[0]),
		.chanx_in_97_(sb_2__1__0_chanx_left_out_97_[0]),
		.chanx_in_98_(sb_1__1__0_chanx_right_out_98_[0]),
		.chanx_in_99_(sb_2__1__0_chanx_left_out_99_[0]),
		.chanx_in_100_(sb_1__1__0_chanx_right_out_100_[0]),
		.chanx_in_101_(sb_2__1__0_chanx_left_out_101_[0]),
		.chanx_in_102_(sb_1__1__0_chanx_right_out_102_[0]),
		.chanx_in_103_(sb_2__1__0_chanx_left_out_103_[0]),
		.chanx_in_104_(sb_1__1__0_chanx_right_out_104_[0]),
		.chanx_in_105_(sb_2__1__0_chanx_left_out_105_[0]),
		.chanx_in_106_(sb_1__1__0_chanx_right_out_106_[0]),
		.chanx_in_107_(sb_2__1__0_chanx_left_out_107_[0]),
		.chanx_in_108_(sb_1__1__0_chanx_right_out_108_[0]),
		.chanx_in_109_(sb_2__1__0_chanx_left_out_109_[0]),
		.chanx_in_110_(sb_1__1__0_chanx_right_out_110_[0]),
		.chanx_in_111_(sb_2__1__0_chanx_left_out_111_[0]),
		.chanx_in_112_(sb_1__1__0_chanx_right_out_112_[0]),
		.chanx_in_113_(sb_2__1__0_chanx_left_out_113_[0]),
		.chanx_in_114_(sb_1__1__0_chanx_right_out_114_[0]),
		.chanx_in_115_(sb_2__1__0_chanx_left_out_115_[0]),
		.chanx_in_116_(sb_1__1__0_chanx_right_out_116_[0]),
		.chanx_in_117_(sb_2__1__0_chanx_left_out_117_[0]),
		.chanx_in_118_(sb_1__1__0_chanx_right_out_118_[0]),
		.chanx_in_119_(sb_2__1__0_chanx_left_out_119_[0]),
		.chanx_in_120_(sb_1__1__0_chanx_right_out_120_[0]),
		.chanx_in_121_(sb_2__1__0_chanx_left_out_121_[0]),
		.chanx_in_122_(sb_1__1__0_chanx_right_out_122_[0]),
		.chanx_in_123_(sb_2__1__0_chanx_left_out_123_[0]),
		.chanx_in_124_(sb_1__1__0_chanx_right_out_124_[0]),
		.chanx_in_125_(sb_2__1__0_chanx_left_out_125_[0]),
		.chanx_in_126_(sb_1__1__0_chanx_right_out_126_[0]),
		.chanx_in_127_(sb_2__1__0_chanx_left_out_127_[0]),
		.chanx_in_128_(sb_1__1__0_chanx_right_out_128_[0]),
		.chanx_in_129_(sb_2__1__0_chanx_left_out_129_[0]),
		.chanx_in_130_(sb_1__1__0_chanx_right_out_130_[0]),
		.chanx_in_131_(sb_2__1__0_chanx_left_out_131_[0]),
		.chanx_in_132_(sb_1__1__0_chanx_right_out_132_[0]),
		.chanx_in_133_(sb_2__1__0_chanx_left_out_133_[0]),
		.chanx_in_134_(sb_1__1__0_chanx_right_out_134_[0]),
		.chanx_in_135_(sb_2__1__0_chanx_left_out_135_[0]),
		.chanx_in_136_(sb_1__1__0_chanx_right_out_136_[0]),
		.chanx_in_137_(sb_2__1__0_chanx_left_out_137_[0]),
		.chanx_in_138_(sb_1__1__0_chanx_right_out_138_[0]),
		.chanx_in_139_(sb_2__1__0_chanx_left_out_139_[0]),
		.chanx_in_140_(sb_1__1__0_chanx_right_out_140_[0]),
		.chanx_in_141_(sb_2__1__0_chanx_left_out_141_[0]),
		.chanx_in_142_(sb_1__1__0_chanx_right_out_142_[0]),
		.chanx_in_143_(sb_2__1__0_chanx_left_out_143_[0]),
		.chanx_in_144_(sb_1__1__0_chanx_right_out_144_[0]),
		.chanx_in_145_(sb_2__1__0_chanx_left_out_145_[0]),
		.chanx_in_146_(sb_1__1__0_chanx_right_out_146_[0]),
		.chanx_in_147_(sb_2__1__0_chanx_left_out_147_[0]),
		.chanx_in_148_(sb_1__1__0_chanx_right_out_148_[0]),
		.chanx_in_149_(sb_2__1__0_chanx_left_out_149_[0]),
		.chanx_in_150_(sb_1__1__0_chanx_right_out_150_[0]),
		.chanx_in_151_(sb_2__1__0_chanx_left_out_151_[0]),
		.chanx_in_152_(sb_1__1__0_chanx_right_out_152_[0]),
		.chanx_in_153_(sb_2__1__0_chanx_left_out_153_[0]),
		.chanx_in_154_(sb_1__1__0_chanx_right_out_154_[0]),
		.chanx_in_155_(sb_2__1__0_chanx_left_out_155_[0]),
		.chanx_in_156_(sb_1__1__0_chanx_right_out_156_[0]),
		.chanx_in_157_(sb_2__1__0_chanx_left_out_157_[0]),
		.chanx_in_158_(sb_1__1__0_chanx_right_out_158_[0]),
		.chanx_in_159_(sb_2__1__0_chanx_left_out_159_[0]),
		.chanx_in_160_(sb_1__1__0_chanx_right_out_160_[0]),
		.chanx_in_161_(sb_2__1__0_chanx_left_out_161_[0]),
		.chanx_in_162_(sb_1__1__0_chanx_right_out_162_[0]),
		.chanx_in_163_(sb_2__1__0_chanx_left_out_163_[0]),
		.chanx_in_164_(sb_1__1__0_chanx_right_out_164_[0]),
		.chanx_in_165_(sb_2__1__0_chanx_left_out_165_[0]),
		.chanx_in_166_(sb_1__1__0_chanx_right_out_166_[0]),
		.chanx_in_167_(sb_2__1__0_chanx_left_out_167_[0]),
		.chanx_in_168_(sb_1__1__0_chanx_right_out_168_[0]),
		.chanx_in_169_(sb_2__1__0_chanx_left_out_169_[0]),
		.chanx_in_170_(sb_1__1__0_chanx_right_out_170_[0]),
		.chanx_in_171_(sb_2__1__0_chanx_left_out_171_[0]),
		.chanx_in_172_(sb_1__1__0_chanx_right_out_172_[0]),
		.chanx_in_173_(sb_2__1__0_chanx_left_out_173_[0]),
		.chanx_in_174_(sb_1__1__0_chanx_right_out_174_[0]),
		.chanx_in_175_(sb_2__1__0_chanx_left_out_175_[0]),
		.chanx_in_176_(sb_1__1__0_chanx_right_out_176_[0]),
		.chanx_in_177_(sb_2__1__0_chanx_left_out_177_[0]),
		.chanx_in_178_(sb_1__1__0_chanx_right_out_178_[0]),
		.chanx_in_179_(sb_2__1__0_chanx_left_out_179_[0]),
		.chanx_in_180_(sb_1__1__0_chanx_right_out_180_[0]),
		.chanx_in_181_(sb_2__1__0_chanx_left_out_181_[0]),
		.chanx_in_182_(sb_1__1__0_chanx_right_out_182_[0]),
		.chanx_in_183_(sb_2__1__0_chanx_left_out_183_[0]),
		.chanx_in_184_(sb_1__1__0_chanx_right_out_184_[0]),
		.chanx_in_185_(sb_2__1__0_chanx_left_out_185_[0]),
		.chanx_in_186_(sb_1__1__0_chanx_right_out_186_[0]),
		.chanx_in_187_(sb_2__1__0_chanx_left_out_187_[0]),
		.chanx_in_188_(sb_1__1__0_chanx_right_out_188_[0]),
		.chanx_in_189_(sb_2__1__0_chanx_left_out_189_[0]),
		.chanx_in_190_(sb_1__1__0_chanx_right_out_190_[0]),
		.chanx_in_191_(sb_2__1__0_chanx_left_out_191_[0]),
		.chanx_in_192_(sb_1__1__0_chanx_right_out_192_[0]),
		.chanx_in_193_(sb_2__1__0_chanx_left_out_193_[0]),
		.chanx_in_194_(sb_1__1__0_chanx_right_out_194_[0]),
		.chanx_in_195_(sb_2__1__0_chanx_left_out_195_[0]),
		.chanx_in_196_(sb_1__1__0_chanx_right_out_196_[0]),
		.chanx_in_197_(sb_2__1__0_chanx_left_out_197_[0]),
		.chanx_in_198_(sb_1__1__0_chanx_right_out_198_[0]),
		.chanx_in_199_(sb_2__1__0_chanx_left_out_199_[0]),
		.ccff_head(sb_2__1__0_ccff_tail[0]),
		.chanx_out_0_(cbx_1__1__1_chanx_out_0_[0]),
		.chanx_out_1_(cbx_1__1__1_chanx_out_1_[0]),
		.chanx_out_2_(cbx_1__1__1_chanx_out_2_[0]),
		.chanx_out_3_(cbx_1__1__1_chanx_out_3_[0]),
		.chanx_out_4_(cbx_1__1__1_chanx_out_4_[0]),
		.chanx_out_5_(cbx_1__1__1_chanx_out_5_[0]),
		.chanx_out_6_(cbx_1__1__1_chanx_out_6_[0]),
		.chanx_out_7_(cbx_1__1__1_chanx_out_7_[0]),
		.chanx_out_8_(cbx_1__1__1_chanx_out_8_[0]),
		.chanx_out_9_(cbx_1__1__1_chanx_out_9_[0]),
		.chanx_out_10_(cbx_1__1__1_chanx_out_10_[0]),
		.chanx_out_11_(cbx_1__1__1_chanx_out_11_[0]),
		.chanx_out_12_(cbx_1__1__1_chanx_out_12_[0]),
		.chanx_out_13_(cbx_1__1__1_chanx_out_13_[0]),
		.chanx_out_14_(cbx_1__1__1_chanx_out_14_[0]),
		.chanx_out_15_(cbx_1__1__1_chanx_out_15_[0]),
		.chanx_out_16_(cbx_1__1__1_chanx_out_16_[0]),
		.chanx_out_17_(cbx_1__1__1_chanx_out_17_[0]),
		.chanx_out_18_(cbx_1__1__1_chanx_out_18_[0]),
		.chanx_out_19_(cbx_1__1__1_chanx_out_19_[0]),
		.chanx_out_20_(cbx_1__1__1_chanx_out_20_[0]),
		.chanx_out_21_(cbx_1__1__1_chanx_out_21_[0]),
		.chanx_out_22_(cbx_1__1__1_chanx_out_22_[0]),
		.chanx_out_23_(cbx_1__1__1_chanx_out_23_[0]),
		.chanx_out_24_(cbx_1__1__1_chanx_out_24_[0]),
		.chanx_out_25_(cbx_1__1__1_chanx_out_25_[0]),
		.chanx_out_26_(cbx_1__1__1_chanx_out_26_[0]),
		.chanx_out_27_(cbx_1__1__1_chanx_out_27_[0]),
		.chanx_out_28_(cbx_1__1__1_chanx_out_28_[0]),
		.chanx_out_29_(cbx_1__1__1_chanx_out_29_[0]),
		.chanx_out_30_(cbx_1__1__1_chanx_out_30_[0]),
		.chanx_out_31_(cbx_1__1__1_chanx_out_31_[0]),
		.chanx_out_32_(cbx_1__1__1_chanx_out_32_[0]),
		.chanx_out_33_(cbx_1__1__1_chanx_out_33_[0]),
		.chanx_out_34_(cbx_1__1__1_chanx_out_34_[0]),
		.chanx_out_35_(cbx_1__1__1_chanx_out_35_[0]),
		.chanx_out_36_(cbx_1__1__1_chanx_out_36_[0]),
		.chanx_out_37_(cbx_1__1__1_chanx_out_37_[0]),
		.chanx_out_38_(cbx_1__1__1_chanx_out_38_[0]),
		.chanx_out_39_(cbx_1__1__1_chanx_out_39_[0]),
		.chanx_out_40_(cbx_1__1__1_chanx_out_40_[0]),
		.chanx_out_41_(cbx_1__1__1_chanx_out_41_[0]),
		.chanx_out_42_(cbx_1__1__1_chanx_out_42_[0]),
		.chanx_out_43_(cbx_1__1__1_chanx_out_43_[0]),
		.chanx_out_44_(cbx_1__1__1_chanx_out_44_[0]),
		.chanx_out_45_(cbx_1__1__1_chanx_out_45_[0]),
		.chanx_out_46_(cbx_1__1__1_chanx_out_46_[0]),
		.chanx_out_47_(cbx_1__1__1_chanx_out_47_[0]),
		.chanx_out_48_(cbx_1__1__1_chanx_out_48_[0]),
		.chanx_out_49_(cbx_1__1__1_chanx_out_49_[0]),
		.chanx_out_50_(cbx_1__1__1_chanx_out_50_[0]),
		.chanx_out_51_(cbx_1__1__1_chanx_out_51_[0]),
		.chanx_out_52_(cbx_1__1__1_chanx_out_52_[0]),
		.chanx_out_53_(cbx_1__1__1_chanx_out_53_[0]),
		.chanx_out_54_(cbx_1__1__1_chanx_out_54_[0]),
		.chanx_out_55_(cbx_1__1__1_chanx_out_55_[0]),
		.chanx_out_56_(cbx_1__1__1_chanx_out_56_[0]),
		.chanx_out_57_(cbx_1__1__1_chanx_out_57_[0]),
		.chanx_out_58_(cbx_1__1__1_chanx_out_58_[0]),
		.chanx_out_59_(cbx_1__1__1_chanx_out_59_[0]),
		.chanx_out_60_(cbx_1__1__1_chanx_out_60_[0]),
		.chanx_out_61_(cbx_1__1__1_chanx_out_61_[0]),
		.chanx_out_62_(cbx_1__1__1_chanx_out_62_[0]),
		.chanx_out_63_(cbx_1__1__1_chanx_out_63_[0]),
		.chanx_out_64_(cbx_1__1__1_chanx_out_64_[0]),
		.chanx_out_65_(cbx_1__1__1_chanx_out_65_[0]),
		.chanx_out_66_(cbx_1__1__1_chanx_out_66_[0]),
		.chanx_out_67_(cbx_1__1__1_chanx_out_67_[0]),
		.chanx_out_68_(cbx_1__1__1_chanx_out_68_[0]),
		.chanx_out_69_(cbx_1__1__1_chanx_out_69_[0]),
		.chanx_out_70_(cbx_1__1__1_chanx_out_70_[0]),
		.chanx_out_71_(cbx_1__1__1_chanx_out_71_[0]),
		.chanx_out_72_(cbx_1__1__1_chanx_out_72_[0]),
		.chanx_out_73_(cbx_1__1__1_chanx_out_73_[0]),
		.chanx_out_74_(cbx_1__1__1_chanx_out_74_[0]),
		.chanx_out_75_(cbx_1__1__1_chanx_out_75_[0]),
		.chanx_out_76_(cbx_1__1__1_chanx_out_76_[0]),
		.chanx_out_77_(cbx_1__1__1_chanx_out_77_[0]),
		.chanx_out_78_(cbx_1__1__1_chanx_out_78_[0]),
		.chanx_out_79_(cbx_1__1__1_chanx_out_79_[0]),
		.chanx_out_80_(cbx_1__1__1_chanx_out_80_[0]),
		.chanx_out_81_(cbx_1__1__1_chanx_out_81_[0]),
		.chanx_out_82_(cbx_1__1__1_chanx_out_82_[0]),
		.chanx_out_83_(cbx_1__1__1_chanx_out_83_[0]),
		.chanx_out_84_(cbx_1__1__1_chanx_out_84_[0]),
		.chanx_out_85_(cbx_1__1__1_chanx_out_85_[0]),
		.chanx_out_86_(cbx_1__1__1_chanx_out_86_[0]),
		.chanx_out_87_(cbx_1__1__1_chanx_out_87_[0]),
		.chanx_out_88_(cbx_1__1__1_chanx_out_88_[0]),
		.chanx_out_89_(cbx_1__1__1_chanx_out_89_[0]),
		.chanx_out_90_(cbx_1__1__1_chanx_out_90_[0]),
		.chanx_out_91_(cbx_1__1__1_chanx_out_91_[0]),
		.chanx_out_92_(cbx_1__1__1_chanx_out_92_[0]),
		.chanx_out_93_(cbx_1__1__1_chanx_out_93_[0]),
		.chanx_out_94_(cbx_1__1__1_chanx_out_94_[0]),
		.chanx_out_95_(cbx_1__1__1_chanx_out_95_[0]),
		.chanx_out_96_(cbx_1__1__1_chanx_out_96_[0]),
		.chanx_out_97_(cbx_1__1__1_chanx_out_97_[0]),
		.chanx_out_98_(cbx_1__1__1_chanx_out_98_[0]),
		.chanx_out_99_(cbx_1__1__1_chanx_out_99_[0]),
		.chanx_out_100_(cbx_1__1__1_chanx_out_100_[0]),
		.chanx_out_101_(cbx_1__1__1_chanx_out_101_[0]),
		.chanx_out_102_(cbx_1__1__1_chanx_out_102_[0]),
		.chanx_out_103_(cbx_1__1__1_chanx_out_103_[0]),
		.chanx_out_104_(cbx_1__1__1_chanx_out_104_[0]),
		.chanx_out_105_(cbx_1__1__1_chanx_out_105_[0]),
		.chanx_out_106_(cbx_1__1__1_chanx_out_106_[0]),
		.chanx_out_107_(cbx_1__1__1_chanx_out_107_[0]),
		.chanx_out_108_(cbx_1__1__1_chanx_out_108_[0]),
		.chanx_out_109_(cbx_1__1__1_chanx_out_109_[0]),
		.chanx_out_110_(cbx_1__1__1_chanx_out_110_[0]),
		.chanx_out_111_(cbx_1__1__1_chanx_out_111_[0]),
		.chanx_out_112_(cbx_1__1__1_chanx_out_112_[0]),
		.chanx_out_113_(cbx_1__1__1_chanx_out_113_[0]),
		.chanx_out_114_(cbx_1__1__1_chanx_out_114_[0]),
		.chanx_out_115_(cbx_1__1__1_chanx_out_115_[0]),
		.chanx_out_116_(cbx_1__1__1_chanx_out_116_[0]),
		.chanx_out_117_(cbx_1__1__1_chanx_out_117_[0]),
		.chanx_out_118_(cbx_1__1__1_chanx_out_118_[0]),
		.chanx_out_119_(cbx_1__1__1_chanx_out_119_[0]),
		.chanx_out_120_(cbx_1__1__1_chanx_out_120_[0]),
		.chanx_out_121_(cbx_1__1__1_chanx_out_121_[0]),
		.chanx_out_122_(cbx_1__1__1_chanx_out_122_[0]),
		.chanx_out_123_(cbx_1__1__1_chanx_out_123_[0]),
		.chanx_out_124_(cbx_1__1__1_chanx_out_124_[0]),
		.chanx_out_125_(cbx_1__1__1_chanx_out_125_[0]),
		.chanx_out_126_(cbx_1__1__1_chanx_out_126_[0]),
		.chanx_out_127_(cbx_1__1__1_chanx_out_127_[0]),
		.chanx_out_128_(cbx_1__1__1_chanx_out_128_[0]),
		.chanx_out_129_(cbx_1__1__1_chanx_out_129_[0]),
		.chanx_out_130_(cbx_1__1__1_chanx_out_130_[0]),
		.chanx_out_131_(cbx_1__1__1_chanx_out_131_[0]),
		.chanx_out_132_(cbx_1__1__1_chanx_out_132_[0]),
		.chanx_out_133_(cbx_1__1__1_chanx_out_133_[0]),
		.chanx_out_134_(cbx_1__1__1_chanx_out_134_[0]),
		.chanx_out_135_(cbx_1__1__1_chanx_out_135_[0]),
		.chanx_out_136_(cbx_1__1__1_chanx_out_136_[0]),
		.chanx_out_137_(cbx_1__1__1_chanx_out_137_[0]),
		.chanx_out_138_(cbx_1__1__1_chanx_out_138_[0]),
		.chanx_out_139_(cbx_1__1__1_chanx_out_139_[0]),
		.chanx_out_140_(cbx_1__1__1_chanx_out_140_[0]),
		.chanx_out_141_(cbx_1__1__1_chanx_out_141_[0]),
		.chanx_out_142_(cbx_1__1__1_chanx_out_142_[0]),
		.chanx_out_143_(cbx_1__1__1_chanx_out_143_[0]),
		.chanx_out_144_(cbx_1__1__1_chanx_out_144_[0]),
		.chanx_out_145_(cbx_1__1__1_chanx_out_145_[0]),
		.chanx_out_146_(cbx_1__1__1_chanx_out_146_[0]),
		.chanx_out_147_(cbx_1__1__1_chanx_out_147_[0]),
		.chanx_out_148_(cbx_1__1__1_chanx_out_148_[0]),
		.chanx_out_149_(cbx_1__1__1_chanx_out_149_[0]),
		.chanx_out_150_(cbx_1__1__1_chanx_out_150_[0]),
		.chanx_out_151_(cbx_1__1__1_chanx_out_151_[0]),
		.chanx_out_152_(cbx_1__1__1_chanx_out_152_[0]),
		.chanx_out_153_(cbx_1__1__1_chanx_out_153_[0]),
		.chanx_out_154_(cbx_1__1__1_chanx_out_154_[0]),
		.chanx_out_155_(cbx_1__1__1_chanx_out_155_[0]),
		.chanx_out_156_(cbx_1__1__1_chanx_out_156_[0]),
		.chanx_out_157_(cbx_1__1__1_chanx_out_157_[0]),
		.chanx_out_158_(cbx_1__1__1_chanx_out_158_[0]),
		.chanx_out_159_(cbx_1__1__1_chanx_out_159_[0]),
		.chanx_out_160_(cbx_1__1__1_chanx_out_160_[0]),
		.chanx_out_161_(cbx_1__1__1_chanx_out_161_[0]),
		.chanx_out_162_(cbx_1__1__1_chanx_out_162_[0]),
		.chanx_out_163_(cbx_1__1__1_chanx_out_163_[0]),
		.chanx_out_164_(cbx_1__1__1_chanx_out_164_[0]),
		.chanx_out_165_(cbx_1__1__1_chanx_out_165_[0]),
		.chanx_out_166_(cbx_1__1__1_chanx_out_166_[0]),
		.chanx_out_167_(cbx_1__1__1_chanx_out_167_[0]),
		.chanx_out_168_(cbx_1__1__1_chanx_out_168_[0]),
		.chanx_out_169_(cbx_1__1__1_chanx_out_169_[0]),
		.chanx_out_170_(cbx_1__1__1_chanx_out_170_[0]),
		.chanx_out_171_(cbx_1__1__1_chanx_out_171_[0]),
		.chanx_out_172_(cbx_1__1__1_chanx_out_172_[0]),
		.chanx_out_173_(cbx_1__1__1_chanx_out_173_[0]),
		.chanx_out_174_(cbx_1__1__1_chanx_out_174_[0]),
		.chanx_out_175_(cbx_1__1__1_chanx_out_175_[0]),
		.chanx_out_176_(cbx_1__1__1_chanx_out_176_[0]),
		.chanx_out_177_(cbx_1__1__1_chanx_out_177_[0]),
		.chanx_out_178_(cbx_1__1__1_chanx_out_178_[0]),
		.chanx_out_179_(cbx_1__1__1_chanx_out_179_[0]),
		.chanx_out_180_(cbx_1__1__1_chanx_out_180_[0]),
		.chanx_out_181_(cbx_1__1__1_chanx_out_181_[0]),
		.chanx_out_182_(cbx_1__1__1_chanx_out_182_[0]),
		.chanx_out_183_(cbx_1__1__1_chanx_out_183_[0]),
		.chanx_out_184_(cbx_1__1__1_chanx_out_184_[0]),
		.chanx_out_185_(cbx_1__1__1_chanx_out_185_[0]),
		.chanx_out_186_(cbx_1__1__1_chanx_out_186_[0]),
		.chanx_out_187_(cbx_1__1__1_chanx_out_187_[0]),
		.chanx_out_188_(cbx_1__1__1_chanx_out_188_[0]),
		.chanx_out_189_(cbx_1__1__1_chanx_out_189_[0]),
		.chanx_out_190_(cbx_1__1__1_chanx_out_190_[0]),
		.chanx_out_191_(cbx_1__1__1_chanx_out_191_[0]),
		.chanx_out_192_(cbx_1__1__1_chanx_out_192_[0]),
		.chanx_out_193_(cbx_1__1__1_chanx_out_193_[0]),
		.chanx_out_194_(cbx_1__1__1_chanx_out_194_[0]),
		.chanx_out_195_(cbx_1__1__1_chanx_out_195_[0]),
		.chanx_out_196_(cbx_1__1__1_chanx_out_196_[0]),
		.chanx_out_197_(cbx_1__1__1_chanx_out_197_[0]),
		.chanx_out_198_(cbx_1__1__1_chanx_out_198_[0]),
		.chanx_out_199_(cbx_1__1__1_chanx_out_199_[0]),
		.top_grid_pin_20_(cbx_1__1__1_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__1_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__1_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__1_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__1_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__1_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__1_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__1_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__1_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__1_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__1_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__1_top_grid_pin_31_[0]),
		.top_grid_pin_32_(cbx_1__1__1_top_grid_pin_32_[0]),
		.top_grid_pin_33_(cbx_1__1__1_top_grid_pin_33_[0]),
		.top_grid_pin_34_(cbx_1__1__1_top_grid_pin_34_[0]),
		.top_grid_pin_35_(cbx_1__1__1_top_grid_pin_35_[0]),
		.top_grid_pin_36_(cbx_1__1__1_top_grid_pin_36_[0]),
		.top_grid_pin_37_(cbx_1__1__1_top_grid_pin_37_[0]),
		.top_grid_pin_38_(cbx_1__1__1_top_grid_pin_38_[0]),
		.top_grid_pin_39_(cbx_1__1__1_top_grid_pin_39_[0]),
		.bottom_grid_pin_42_(cbx_1__1__1_bottom_grid_pin_42_[0]),
		.bottom_grid_pin_43_(cbx_1__1__1_bottom_grid_pin_43_[0]),
		.bottom_grid_pin_69_(cbx_1__1__1_bottom_grid_pin_69_[0]),
		.ccff_tail(cbx_1__1__1_ccff_tail[0]));

	cbx_1__2_ cbx_1__2_ (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.chanx_in_0_(sb_0__2__0_chanx_right_out_0_[0]),
		.chanx_in_1_(sb_1__2__0_chanx_left_out_1_[0]),
		.chanx_in_2_(sb_0__2__0_chanx_right_out_2_[0]),
		.chanx_in_3_(sb_1__2__0_chanx_left_out_3_[0]),
		.chanx_in_4_(sb_0__2__0_chanx_right_out_4_[0]),
		.chanx_in_5_(sb_1__2__0_chanx_left_out_5_[0]),
		.chanx_in_6_(sb_0__2__0_chanx_right_out_6_[0]),
		.chanx_in_7_(sb_1__2__0_chanx_left_out_7_[0]),
		.chanx_in_8_(sb_0__2__0_chanx_right_out_8_[0]),
		.chanx_in_9_(sb_1__2__0_chanx_left_out_9_[0]),
		.chanx_in_10_(sb_0__2__0_chanx_right_out_10_[0]),
		.chanx_in_11_(sb_1__2__0_chanx_left_out_11_[0]),
		.chanx_in_12_(sb_0__2__0_chanx_right_out_12_[0]),
		.chanx_in_13_(sb_1__2__0_chanx_left_out_13_[0]),
		.chanx_in_14_(sb_0__2__0_chanx_right_out_14_[0]),
		.chanx_in_15_(sb_1__2__0_chanx_left_out_15_[0]),
		.chanx_in_16_(sb_0__2__0_chanx_right_out_16_[0]),
		.chanx_in_17_(sb_1__2__0_chanx_left_out_17_[0]),
		.chanx_in_18_(sb_0__2__0_chanx_right_out_18_[0]),
		.chanx_in_19_(sb_1__2__0_chanx_left_out_19_[0]),
		.chanx_in_20_(sb_0__2__0_chanx_right_out_20_[0]),
		.chanx_in_21_(sb_1__2__0_chanx_left_out_21_[0]),
		.chanx_in_22_(sb_0__2__0_chanx_right_out_22_[0]),
		.chanx_in_23_(sb_1__2__0_chanx_left_out_23_[0]),
		.chanx_in_24_(sb_0__2__0_chanx_right_out_24_[0]),
		.chanx_in_25_(sb_1__2__0_chanx_left_out_25_[0]),
		.chanx_in_26_(sb_0__2__0_chanx_right_out_26_[0]),
		.chanx_in_27_(sb_1__2__0_chanx_left_out_27_[0]),
		.chanx_in_28_(sb_0__2__0_chanx_right_out_28_[0]),
		.chanx_in_29_(sb_1__2__0_chanx_left_out_29_[0]),
		.chanx_in_30_(sb_0__2__0_chanx_right_out_30_[0]),
		.chanx_in_31_(sb_1__2__0_chanx_left_out_31_[0]),
		.chanx_in_32_(sb_0__2__0_chanx_right_out_32_[0]),
		.chanx_in_33_(sb_1__2__0_chanx_left_out_33_[0]),
		.chanx_in_34_(sb_0__2__0_chanx_right_out_34_[0]),
		.chanx_in_35_(sb_1__2__0_chanx_left_out_35_[0]),
		.chanx_in_36_(sb_0__2__0_chanx_right_out_36_[0]),
		.chanx_in_37_(sb_1__2__0_chanx_left_out_37_[0]),
		.chanx_in_38_(sb_0__2__0_chanx_right_out_38_[0]),
		.chanx_in_39_(sb_1__2__0_chanx_left_out_39_[0]),
		.chanx_in_40_(sb_0__2__0_chanx_right_out_40_[0]),
		.chanx_in_41_(sb_1__2__0_chanx_left_out_41_[0]),
		.chanx_in_42_(sb_0__2__0_chanx_right_out_42_[0]),
		.chanx_in_43_(sb_1__2__0_chanx_left_out_43_[0]),
		.chanx_in_44_(sb_0__2__0_chanx_right_out_44_[0]),
		.chanx_in_45_(sb_1__2__0_chanx_left_out_45_[0]),
		.chanx_in_46_(sb_0__2__0_chanx_right_out_46_[0]),
		.chanx_in_47_(sb_1__2__0_chanx_left_out_47_[0]),
		.chanx_in_48_(sb_0__2__0_chanx_right_out_48_[0]),
		.chanx_in_49_(sb_1__2__0_chanx_left_out_49_[0]),
		.chanx_in_50_(sb_0__2__0_chanx_right_out_50_[0]),
		.chanx_in_51_(sb_1__2__0_chanx_left_out_51_[0]),
		.chanx_in_52_(sb_0__2__0_chanx_right_out_52_[0]),
		.chanx_in_53_(sb_1__2__0_chanx_left_out_53_[0]),
		.chanx_in_54_(sb_0__2__0_chanx_right_out_54_[0]),
		.chanx_in_55_(sb_1__2__0_chanx_left_out_55_[0]),
		.chanx_in_56_(sb_0__2__0_chanx_right_out_56_[0]),
		.chanx_in_57_(sb_1__2__0_chanx_left_out_57_[0]),
		.chanx_in_58_(sb_0__2__0_chanx_right_out_58_[0]),
		.chanx_in_59_(sb_1__2__0_chanx_left_out_59_[0]),
		.chanx_in_60_(sb_0__2__0_chanx_right_out_60_[0]),
		.chanx_in_61_(sb_1__2__0_chanx_left_out_61_[0]),
		.chanx_in_62_(sb_0__2__0_chanx_right_out_62_[0]),
		.chanx_in_63_(sb_1__2__0_chanx_left_out_63_[0]),
		.chanx_in_64_(sb_0__2__0_chanx_right_out_64_[0]),
		.chanx_in_65_(sb_1__2__0_chanx_left_out_65_[0]),
		.chanx_in_66_(sb_0__2__0_chanx_right_out_66_[0]),
		.chanx_in_67_(sb_1__2__0_chanx_left_out_67_[0]),
		.chanx_in_68_(sb_0__2__0_chanx_right_out_68_[0]),
		.chanx_in_69_(sb_1__2__0_chanx_left_out_69_[0]),
		.chanx_in_70_(sb_0__2__0_chanx_right_out_70_[0]),
		.chanx_in_71_(sb_1__2__0_chanx_left_out_71_[0]),
		.chanx_in_72_(sb_0__2__0_chanx_right_out_72_[0]),
		.chanx_in_73_(sb_1__2__0_chanx_left_out_73_[0]),
		.chanx_in_74_(sb_0__2__0_chanx_right_out_74_[0]),
		.chanx_in_75_(sb_1__2__0_chanx_left_out_75_[0]),
		.chanx_in_76_(sb_0__2__0_chanx_right_out_76_[0]),
		.chanx_in_77_(sb_1__2__0_chanx_left_out_77_[0]),
		.chanx_in_78_(sb_0__2__0_chanx_right_out_78_[0]),
		.chanx_in_79_(sb_1__2__0_chanx_left_out_79_[0]),
		.chanx_in_80_(sb_0__2__0_chanx_right_out_80_[0]),
		.chanx_in_81_(sb_1__2__0_chanx_left_out_81_[0]),
		.chanx_in_82_(sb_0__2__0_chanx_right_out_82_[0]),
		.chanx_in_83_(sb_1__2__0_chanx_left_out_83_[0]),
		.chanx_in_84_(sb_0__2__0_chanx_right_out_84_[0]),
		.chanx_in_85_(sb_1__2__0_chanx_left_out_85_[0]),
		.chanx_in_86_(sb_0__2__0_chanx_right_out_86_[0]),
		.chanx_in_87_(sb_1__2__0_chanx_left_out_87_[0]),
		.chanx_in_88_(sb_0__2__0_chanx_right_out_88_[0]),
		.chanx_in_89_(sb_1__2__0_chanx_left_out_89_[0]),
		.chanx_in_90_(sb_0__2__0_chanx_right_out_90_[0]),
		.chanx_in_91_(sb_1__2__0_chanx_left_out_91_[0]),
		.chanx_in_92_(sb_0__2__0_chanx_right_out_92_[0]),
		.chanx_in_93_(sb_1__2__0_chanx_left_out_93_[0]),
		.chanx_in_94_(sb_0__2__0_chanx_right_out_94_[0]),
		.chanx_in_95_(sb_1__2__0_chanx_left_out_95_[0]),
		.chanx_in_96_(sb_0__2__0_chanx_right_out_96_[0]),
		.chanx_in_97_(sb_1__2__0_chanx_left_out_97_[0]),
		.chanx_in_98_(sb_0__2__0_chanx_right_out_98_[0]),
		.chanx_in_99_(sb_1__2__0_chanx_left_out_99_[0]),
		.chanx_in_100_(sb_0__2__0_chanx_right_out_100_[0]),
		.chanx_in_101_(sb_1__2__0_chanx_left_out_101_[0]),
		.chanx_in_102_(sb_0__2__0_chanx_right_out_102_[0]),
		.chanx_in_103_(sb_1__2__0_chanx_left_out_103_[0]),
		.chanx_in_104_(sb_0__2__0_chanx_right_out_104_[0]),
		.chanx_in_105_(sb_1__2__0_chanx_left_out_105_[0]),
		.chanx_in_106_(sb_0__2__0_chanx_right_out_106_[0]),
		.chanx_in_107_(sb_1__2__0_chanx_left_out_107_[0]),
		.chanx_in_108_(sb_0__2__0_chanx_right_out_108_[0]),
		.chanx_in_109_(sb_1__2__0_chanx_left_out_109_[0]),
		.chanx_in_110_(sb_0__2__0_chanx_right_out_110_[0]),
		.chanx_in_111_(sb_1__2__0_chanx_left_out_111_[0]),
		.chanx_in_112_(sb_0__2__0_chanx_right_out_112_[0]),
		.chanx_in_113_(sb_1__2__0_chanx_left_out_113_[0]),
		.chanx_in_114_(sb_0__2__0_chanx_right_out_114_[0]),
		.chanx_in_115_(sb_1__2__0_chanx_left_out_115_[0]),
		.chanx_in_116_(sb_0__2__0_chanx_right_out_116_[0]),
		.chanx_in_117_(sb_1__2__0_chanx_left_out_117_[0]),
		.chanx_in_118_(sb_0__2__0_chanx_right_out_118_[0]),
		.chanx_in_119_(sb_1__2__0_chanx_left_out_119_[0]),
		.chanx_in_120_(sb_0__2__0_chanx_right_out_120_[0]),
		.chanx_in_121_(sb_1__2__0_chanx_left_out_121_[0]),
		.chanx_in_122_(sb_0__2__0_chanx_right_out_122_[0]),
		.chanx_in_123_(sb_1__2__0_chanx_left_out_123_[0]),
		.chanx_in_124_(sb_0__2__0_chanx_right_out_124_[0]),
		.chanx_in_125_(sb_1__2__0_chanx_left_out_125_[0]),
		.chanx_in_126_(sb_0__2__0_chanx_right_out_126_[0]),
		.chanx_in_127_(sb_1__2__0_chanx_left_out_127_[0]),
		.chanx_in_128_(sb_0__2__0_chanx_right_out_128_[0]),
		.chanx_in_129_(sb_1__2__0_chanx_left_out_129_[0]),
		.chanx_in_130_(sb_0__2__0_chanx_right_out_130_[0]),
		.chanx_in_131_(sb_1__2__0_chanx_left_out_131_[0]),
		.chanx_in_132_(sb_0__2__0_chanx_right_out_132_[0]),
		.chanx_in_133_(sb_1__2__0_chanx_left_out_133_[0]),
		.chanx_in_134_(sb_0__2__0_chanx_right_out_134_[0]),
		.chanx_in_135_(sb_1__2__0_chanx_left_out_135_[0]),
		.chanx_in_136_(sb_0__2__0_chanx_right_out_136_[0]),
		.chanx_in_137_(sb_1__2__0_chanx_left_out_137_[0]),
		.chanx_in_138_(sb_0__2__0_chanx_right_out_138_[0]),
		.chanx_in_139_(sb_1__2__0_chanx_left_out_139_[0]),
		.chanx_in_140_(sb_0__2__0_chanx_right_out_140_[0]),
		.chanx_in_141_(sb_1__2__0_chanx_left_out_141_[0]),
		.chanx_in_142_(sb_0__2__0_chanx_right_out_142_[0]),
		.chanx_in_143_(sb_1__2__0_chanx_left_out_143_[0]),
		.chanx_in_144_(sb_0__2__0_chanx_right_out_144_[0]),
		.chanx_in_145_(sb_1__2__0_chanx_left_out_145_[0]),
		.chanx_in_146_(sb_0__2__0_chanx_right_out_146_[0]),
		.chanx_in_147_(sb_1__2__0_chanx_left_out_147_[0]),
		.chanx_in_148_(sb_0__2__0_chanx_right_out_148_[0]),
		.chanx_in_149_(sb_1__2__0_chanx_left_out_149_[0]),
		.chanx_in_150_(sb_0__2__0_chanx_right_out_150_[0]),
		.chanx_in_151_(sb_1__2__0_chanx_left_out_151_[0]),
		.chanx_in_152_(sb_0__2__0_chanx_right_out_152_[0]),
		.chanx_in_153_(sb_1__2__0_chanx_left_out_153_[0]),
		.chanx_in_154_(sb_0__2__0_chanx_right_out_154_[0]),
		.chanx_in_155_(sb_1__2__0_chanx_left_out_155_[0]),
		.chanx_in_156_(sb_0__2__0_chanx_right_out_156_[0]),
		.chanx_in_157_(sb_1__2__0_chanx_left_out_157_[0]),
		.chanx_in_158_(sb_0__2__0_chanx_right_out_158_[0]),
		.chanx_in_159_(sb_1__2__0_chanx_left_out_159_[0]),
		.chanx_in_160_(sb_0__2__0_chanx_right_out_160_[0]),
		.chanx_in_161_(sb_1__2__0_chanx_left_out_161_[0]),
		.chanx_in_162_(sb_0__2__0_chanx_right_out_162_[0]),
		.chanx_in_163_(sb_1__2__0_chanx_left_out_163_[0]),
		.chanx_in_164_(sb_0__2__0_chanx_right_out_164_[0]),
		.chanx_in_165_(sb_1__2__0_chanx_left_out_165_[0]),
		.chanx_in_166_(sb_0__2__0_chanx_right_out_166_[0]),
		.chanx_in_167_(sb_1__2__0_chanx_left_out_167_[0]),
		.chanx_in_168_(sb_0__2__0_chanx_right_out_168_[0]),
		.chanx_in_169_(sb_1__2__0_chanx_left_out_169_[0]),
		.chanx_in_170_(sb_0__2__0_chanx_right_out_170_[0]),
		.chanx_in_171_(sb_1__2__0_chanx_left_out_171_[0]),
		.chanx_in_172_(sb_0__2__0_chanx_right_out_172_[0]),
		.chanx_in_173_(sb_1__2__0_chanx_left_out_173_[0]),
		.chanx_in_174_(sb_0__2__0_chanx_right_out_174_[0]),
		.chanx_in_175_(sb_1__2__0_chanx_left_out_175_[0]),
		.chanx_in_176_(sb_0__2__0_chanx_right_out_176_[0]),
		.chanx_in_177_(sb_1__2__0_chanx_left_out_177_[0]),
		.chanx_in_178_(sb_0__2__0_chanx_right_out_178_[0]),
		.chanx_in_179_(sb_1__2__0_chanx_left_out_179_[0]),
		.chanx_in_180_(sb_0__2__0_chanx_right_out_180_[0]),
		.chanx_in_181_(sb_1__2__0_chanx_left_out_181_[0]),
		.chanx_in_182_(sb_0__2__0_chanx_right_out_182_[0]),
		.chanx_in_183_(sb_1__2__0_chanx_left_out_183_[0]),
		.chanx_in_184_(sb_0__2__0_chanx_right_out_184_[0]),
		.chanx_in_185_(sb_1__2__0_chanx_left_out_185_[0]),
		.chanx_in_186_(sb_0__2__0_chanx_right_out_186_[0]),
		.chanx_in_187_(sb_1__2__0_chanx_left_out_187_[0]),
		.chanx_in_188_(sb_0__2__0_chanx_right_out_188_[0]),
		.chanx_in_189_(sb_1__2__0_chanx_left_out_189_[0]),
		.chanx_in_190_(sb_0__2__0_chanx_right_out_190_[0]),
		.chanx_in_191_(sb_1__2__0_chanx_left_out_191_[0]),
		.chanx_in_192_(sb_0__2__0_chanx_right_out_192_[0]),
		.chanx_in_193_(sb_1__2__0_chanx_left_out_193_[0]),
		.chanx_in_194_(sb_0__2__0_chanx_right_out_194_[0]),
		.chanx_in_195_(sb_1__2__0_chanx_left_out_195_[0]),
		.chanx_in_196_(sb_0__2__0_chanx_right_out_196_[0]),
		.chanx_in_197_(sb_1__2__0_chanx_left_out_197_[0]),
		.chanx_in_198_(sb_0__2__0_chanx_right_out_198_[0]),
		.chanx_in_199_(sb_1__2__0_chanx_left_out_199_[0]),
		.ccff_head(sb_1__2__0_ccff_tail[0]),
		.chanx_out_0_(cbx_1__2__0_chanx_out_0_[0]),
		.chanx_out_1_(cbx_1__2__0_chanx_out_1_[0]),
		.chanx_out_2_(cbx_1__2__0_chanx_out_2_[0]),
		.chanx_out_3_(cbx_1__2__0_chanx_out_3_[0]),
		.chanx_out_4_(cbx_1__2__0_chanx_out_4_[0]),
		.chanx_out_5_(cbx_1__2__0_chanx_out_5_[0]),
		.chanx_out_6_(cbx_1__2__0_chanx_out_6_[0]),
		.chanx_out_7_(cbx_1__2__0_chanx_out_7_[0]),
		.chanx_out_8_(cbx_1__2__0_chanx_out_8_[0]),
		.chanx_out_9_(cbx_1__2__0_chanx_out_9_[0]),
		.chanx_out_10_(cbx_1__2__0_chanx_out_10_[0]),
		.chanx_out_11_(cbx_1__2__0_chanx_out_11_[0]),
		.chanx_out_12_(cbx_1__2__0_chanx_out_12_[0]),
		.chanx_out_13_(cbx_1__2__0_chanx_out_13_[0]),
		.chanx_out_14_(cbx_1__2__0_chanx_out_14_[0]),
		.chanx_out_15_(cbx_1__2__0_chanx_out_15_[0]),
		.chanx_out_16_(cbx_1__2__0_chanx_out_16_[0]),
		.chanx_out_17_(cbx_1__2__0_chanx_out_17_[0]),
		.chanx_out_18_(cbx_1__2__0_chanx_out_18_[0]),
		.chanx_out_19_(cbx_1__2__0_chanx_out_19_[0]),
		.chanx_out_20_(cbx_1__2__0_chanx_out_20_[0]),
		.chanx_out_21_(cbx_1__2__0_chanx_out_21_[0]),
		.chanx_out_22_(cbx_1__2__0_chanx_out_22_[0]),
		.chanx_out_23_(cbx_1__2__0_chanx_out_23_[0]),
		.chanx_out_24_(cbx_1__2__0_chanx_out_24_[0]),
		.chanx_out_25_(cbx_1__2__0_chanx_out_25_[0]),
		.chanx_out_26_(cbx_1__2__0_chanx_out_26_[0]),
		.chanx_out_27_(cbx_1__2__0_chanx_out_27_[0]),
		.chanx_out_28_(cbx_1__2__0_chanx_out_28_[0]),
		.chanx_out_29_(cbx_1__2__0_chanx_out_29_[0]),
		.chanx_out_30_(cbx_1__2__0_chanx_out_30_[0]),
		.chanx_out_31_(cbx_1__2__0_chanx_out_31_[0]),
		.chanx_out_32_(cbx_1__2__0_chanx_out_32_[0]),
		.chanx_out_33_(cbx_1__2__0_chanx_out_33_[0]),
		.chanx_out_34_(cbx_1__2__0_chanx_out_34_[0]),
		.chanx_out_35_(cbx_1__2__0_chanx_out_35_[0]),
		.chanx_out_36_(cbx_1__2__0_chanx_out_36_[0]),
		.chanx_out_37_(cbx_1__2__0_chanx_out_37_[0]),
		.chanx_out_38_(cbx_1__2__0_chanx_out_38_[0]),
		.chanx_out_39_(cbx_1__2__0_chanx_out_39_[0]),
		.chanx_out_40_(cbx_1__2__0_chanx_out_40_[0]),
		.chanx_out_41_(cbx_1__2__0_chanx_out_41_[0]),
		.chanx_out_42_(cbx_1__2__0_chanx_out_42_[0]),
		.chanx_out_43_(cbx_1__2__0_chanx_out_43_[0]),
		.chanx_out_44_(cbx_1__2__0_chanx_out_44_[0]),
		.chanx_out_45_(cbx_1__2__0_chanx_out_45_[0]),
		.chanx_out_46_(cbx_1__2__0_chanx_out_46_[0]),
		.chanx_out_47_(cbx_1__2__0_chanx_out_47_[0]),
		.chanx_out_48_(cbx_1__2__0_chanx_out_48_[0]),
		.chanx_out_49_(cbx_1__2__0_chanx_out_49_[0]),
		.chanx_out_50_(cbx_1__2__0_chanx_out_50_[0]),
		.chanx_out_51_(cbx_1__2__0_chanx_out_51_[0]),
		.chanx_out_52_(cbx_1__2__0_chanx_out_52_[0]),
		.chanx_out_53_(cbx_1__2__0_chanx_out_53_[0]),
		.chanx_out_54_(cbx_1__2__0_chanx_out_54_[0]),
		.chanx_out_55_(cbx_1__2__0_chanx_out_55_[0]),
		.chanx_out_56_(cbx_1__2__0_chanx_out_56_[0]),
		.chanx_out_57_(cbx_1__2__0_chanx_out_57_[0]),
		.chanx_out_58_(cbx_1__2__0_chanx_out_58_[0]),
		.chanx_out_59_(cbx_1__2__0_chanx_out_59_[0]),
		.chanx_out_60_(cbx_1__2__0_chanx_out_60_[0]),
		.chanx_out_61_(cbx_1__2__0_chanx_out_61_[0]),
		.chanx_out_62_(cbx_1__2__0_chanx_out_62_[0]),
		.chanx_out_63_(cbx_1__2__0_chanx_out_63_[0]),
		.chanx_out_64_(cbx_1__2__0_chanx_out_64_[0]),
		.chanx_out_65_(cbx_1__2__0_chanx_out_65_[0]),
		.chanx_out_66_(cbx_1__2__0_chanx_out_66_[0]),
		.chanx_out_67_(cbx_1__2__0_chanx_out_67_[0]),
		.chanx_out_68_(cbx_1__2__0_chanx_out_68_[0]),
		.chanx_out_69_(cbx_1__2__0_chanx_out_69_[0]),
		.chanx_out_70_(cbx_1__2__0_chanx_out_70_[0]),
		.chanx_out_71_(cbx_1__2__0_chanx_out_71_[0]),
		.chanx_out_72_(cbx_1__2__0_chanx_out_72_[0]),
		.chanx_out_73_(cbx_1__2__0_chanx_out_73_[0]),
		.chanx_out_74_(cbx_1__2__0_chanx_out_74_[0]),
		.chanx_out_75_(cbx_1__2__0_chanx_out_75_[0]),
		.chanx_out_76_(cbx_1__2__0_chanx_out_76_[0]),
		.chanx_out_77_(cbx_1__2__0_chanx_out_77_[0]),
		.chanx_out_78_(cbx_1__2__0_chanx_out_78_[0]),
		.chanx_out_79_(cbx_1__2__0_chanx_out_79_[0]),
		.chanx_out_80_(cbx_1__2__0_chanx_out_80_[0]),
		.chanx_out_81_(cbx_1__2__0_chanx_out_81_[0]),
		.chanx_out_82_(cbx_1__2__0_chanx_out_82_[0]),
		.chanx_out_83_(cbx_1__2__0_chanx_out_83_[0]),
		.chanx_out_84_(cbx_1__2__0_chanx_out_84_[0]),
		.chanx_out_85_(cbx_1__2__0_chanx_out_85_[0]),
		.chanx_out_86_(cbx_1__2__0_chanx_out_86_[0]),
		.chanx_out_87_(cbx_1__2__0_chanx_out_87_[0]),
		.chanx_out_88_(cbx_1__2__0_chanx_out_88_[0]),
		.chanx_out_89_(cbx_1__2__0_chanx_out_89_[0]),
		.chanx_out_90_(cbx_1__2__0_chanx_out_90_[0]),
		.chanx_out_91_(cbx_1__2__0_chanx_out_91_[0]),
		.chanx_out_92_(cbx_1__2__0_chanx_out_92_[0]),
		.chanx_out_93_(cbx_1__2__0_chanx_out_93_[0]),
		.chanx_out_94_(cbx_1__2__0_chanx_out_94_[0]),
		.chanx_out_95_(cbx_1__2__0_chanx_out_95_[0]),
		.chanx_out_96_(cbx_1__2__0_chanx_out_96_[0]),
		.chanx_out_97_(cbx_1__2__0_chanx_out_97_[0]),
		.chanx_out_98_(cbx_1__2__0_chanx_out_98_[0]),
		.chanx_out_99_(cbx_1__2__0_chanx_out_99_[0]),
		.chanx_out_100_(cbx_1__2__0_chanx_out_100_[0]),
		.chanx_out_101_(cbx_1__2__0_chanx_out_101_[0]),
		.chanx_out_102_(cbx_1__2__0_chanx_out_102_[0]),
		.chanx_out_103_(cbx_1__2__0_chanx_out_103_[0]),
		.chanx_out_104_(cbx_1__2__0_chanx_out_104_[0]),
		.chanx_out_105_(cbx_1__2__0_chanx_out_105_[0]),
		.chanx_out_106_(cbx_1__2__0_chanx_out_106_[0]),
		.chanx_out_107_(cbx_1__2__0_chanx_out_107_[0]),
		.chanx_out_108_(cbx_1__2__0_chanx_out_108_[0]),
		.chanx_out_109_(cbx_1__2__0_chanx_out_109_[0]),
		.chanx_out_110_(cbx_1__2__0_chanx_out_110_[0]),
		.chanx_out_111_(cbx_1__2__0_chanx_out_111_[0]),
		.chanx_out_112_(cbx_1__2__0_chanx_out_112_[0]),
		.chanx_out_113_(cbx_1__2__0_chanx_out_113_[0]),
		.chanx_out_114_(cbx_1__2__0_chanx_out_114_[0]),
		.chanx_out_115_(cbx_1__2__0_chanx_out_115_[0]),
		.chanx_out_116_(cbx_1__2__0_chanx_out_116_[0]),
		.chanx_out_117_(cbx_1__2__0_chanx_out_117_[0]),
		.chanx_out_118_(cbx_1__2__0_chanx_out_118_[0]),
		.chanx_out_119_(cbx_1__2__0_chanx_out_119_[0]),
		.chanx_out_120_(cbx_1__2__0_chanx_out_120_[0]),
		.chanx_out_121_(cbx_1__2__0_chanx_out_121_[0]),
		.chanx_out_122_(cbx_1__2__0_chanx_out_122_[0]),
		.chanx_out_123_(cbx_1__2__0_chanx_out_123_[0]),
		.chanx_out_124_(cbx_1__2__0_chanx_out_124_[0]),
		.chanx_out_125_(cbx_1__2__0_chanx_out_125_[0]),
		.chanx_out_126_(cbx_1__2__0_chanx_out_126_[0]),
		.chanx_out_127_(cbx_1__2__0_chanx_out_127_[0]),
		.chanx_out_128_(cbx_1__2__0_chanx_out_128_[0]),
		.chanx_out_129_(cbx_1__2__0_chanx_out_129_[0]),
		.chanx_out_130_(cbx_1__2__0_chanx_out_130_[0]),
		.chanx_out_131_(cbx_1__2__0_chanx_out_131_[0]),
		.chanx_out_132_(cbx_1__2__0_chanx_out_132_[0]),
		.chanx_out_133_(cbx_1__2__0_chanx_out_133_[0]),
		.chanx_out_134_(cbx_1__2__0_chanx_out_134_[0]),
		.chanx_out_135_(cbx_1__2__0_chanx_out_135_[0]),
		.chanx_out_136_(cbx_1__2__0_chanx_out_136_[0]),
		.chanx_out_137_(cbx_1__2__0_chanx_out_137_[0]),
		.chanx_out_138_(cbx_1__2__0_chanx_out_138_[0]),
		.chanx_out_139_(cbx_1__2__0_chanx_out_139_[0]),
		.chanx_out_140_(cbx_1__2__0_chanx_out_140_[0]),
		.chanx_out_141_(cbx_1__2__0_chanx_out_141_[0]),
		.chanx_out_142_(cbx_1__2__0_chanx_out_142_[0]),
		.chanx_out_143_(cbx_1__2__0_chanx_out_143_[0]),
		.chanx_out_144_(cbx_1__2__0_chanx_out_144_[0]),
		.chanx_out_145_(cbx_1__2__0_chanx_out_145_[0]),
		.chanx_out_146_(cbx_1__2__0_chanx_out_146_[0]),
		.chanx_out_147_(cbx_1__2__0_chanx_out_147_[0]),
		.chanx_out_148_(cbx_1__2__0_chanx_out_148_[0]),
		.chanx_out_149_(cbx_1__2__0_chanx_out_149_[0]),
		.chanx_out_150_(cbx_1__2__0_chanx_out_150_[0]),
		.chanx_out_151_(cbx_1__2__0_chanx_out_151_[0]),
		.chanx_out_152_(cbx_1__2__0_chanx_out_152_[0]),
		.chanx_out_153_(cbx_1__2__0_chanx_out_153_[0]),
		.chanx_out_154_(cbx_1__2__0_chanx_out_154_[0]),
		.chanx_out_155_(cbx_1__2__0_chanx_out_155_[0]),
		.chanx_out_156_(cbx_1__2__0_chanx_out_156_[0]),
		.chanx_out_157_(cbx_1__2__0_chanx_out_157_[0]),
		.chanx_out_158_(cbx_1__2__0_chanx_out_158_[0]),
		.chanx_out_159_(cbx_1__2__0_chanx_out_159_[0]),
		.chanx_out_160_(cbx_1__2__0_chanx_out_160_[0]),
		.chanx_out_161_(cbx_1__2__0_chanx_out_161_[0]),
		.chanx_out_162_(cbx_1__2__0_chanx_out_162_[0]),
		.chanx_out_163_(cbx_1__2__0_chanx_out_163_[0]),
		.chanx_out_164_(cbx_1__2__0_chanx_out_164_[0]),
		.chanx_out_165_(cbx_1__2__0_chanx_out_165_[0]),
		.chanx_out_166_(cbx_1__2__0_chanx_out_166_[0]),
		.chanx_out_167_(cbx_1__2__0_chanx_out_167_[0]),
		.chanx_out_168_(cbx_1__2__0_chanx_out_168_[0]),
		.chanx_out_169_(cbx_1__2__0_chanx_out_169_[0]),
		.chanx_out_170_(cbx_1__2__0_chanx_out_170_[0]),
		.chanx_out_171_(cbx_1__2__0_chanx_out_171_[0]),
		.chanx_out_172_(cbx_1__2__0_chanx_out_172_[0]),
		.chanx_out_173_(cbx_1__2__0_chanx_out_173_[0]),
		.chanx_out_174_(cbx_1__2__0_chanx_out_174_[0]),
		.chanx_out_175_(cbx_1__2__0_chanx_out_175_[0]),
		.chanx_out_176_(cbx_1__2__0_chanx_out_176_[0]),
		.chanx_out_177_(cbx_1__2__0_chanx_out_177_[0]),
		.chanx_out_178_(cbx_1__2__0_chanx_out_178_[0]),
		.chanx_out_179_(cbx_1__2__0_chanx_out_179_[0]),
		.chanx_out_180_(cbx_1__2__0_chanx_out_180_[0]),
		.chanx_out_181_(cbx_1__2__0_chanx_out_181_[0]),
		.chanx_out_182_(cbx_1__2__0_chanx_out_182_[0]),
		.chanx_out_183_(cbx_1__2__0_chanx_out_183_[0]),
		.chanx_out_184_(cbx_1__2__0_chanx_out_184_[0]),
		.chanx_out_185_(cbx_1__2__0_chanx_out_185_[0]),
		.chanx_out_186_(cbx_1__2__0_chanx_out_186_[0]),
		.chanx_out_187_(cbx_1__2__0_chanx_out_187_[0]),
		.chanx_out_188_(cbx_1__2__0_chanx_out_188_[0]),
		.chanx_out_189_(cbx_1__2__0_chanx_out_189_[0]),
		.chanx_out_190_(cbx_1__2__0_chanx_out_190_[0]),
		.chanx_out_191_(cbx_1__2__0_chanx_out_191_[0]),
		.chanx_out_192_(cbx_1__2__0_chanx_out_192_[0]),
		.chanx_out_193_(cbx_1__2__0_chanx_out_193_[0]),
		.chanx_out_194_(cbx_1__2__0_chanx_out_194_[0]),
		.chanx_out_195_(cbx_1__2__0_chanx_out_195_[0]),
		.chanx_out_196_(cbx_1__2__0_chanx_out_196_[0]),
		.chanx_out_197_(cbx_1__2__0_chanx_out_197_[0]),
		.chanx_out_198_(cbx_1__2__0_chanx_out_198_[0]),
		.chanx_out_199_(cbx_1__2__0_chanx_out_199_[0]),
		.top_grid_pin_0_(cbx_1__2__0_top_grid_pin_0_[0]),
		.bottom_grid_pin_42_(cbx_1__2__0_bottom_grid_pin_42_[0]),
		.bottom_grid_pin_43_(cbx_1__2__0_bottom_grid_pin_43_[0]),
		.bottom_grid_pin_68_(cbx_1__2__0_bottom_grid_pin_68_[0]),
		.ccff_tail(cbx_1__2__0_ccff_tail[0]));

	cbx_1__2_ cbx_2__2_ (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.chanx_in_0_(sb_1__2__0_chanx_right_out_0_[0]),
		.chanx_in_1_(sb_2__2__0_chanx_left_out_1_[0]),
		.chanx_in_2_(sb_1__2__0_chanx_right_out_2_[0]),
		.chanx_in_3_(sb_2__2__0_chanx_left_out_3_[0]),
		.chanx_in_4_(sb_1__2__0_chanx_right_out_4_[0]),
		.chanx_in_5_(sb_2__2__0_chanx_left_out_5_[0]),
		.chanx_in_6_(sb_1__2__0_chanx_right_out_6_[0]),
		.chanx_in_7_(sb_2__2__0_chanx_left_out_7_[0]),
		.chanx_in_8_(sb_1__2__0_chanx_right_out_8_[0]),
		.chanx_in_9_(sb_2__2__0_chanx_left_out_9_[0]),
		.chanx_in_10_(sb_1__2__0_chanx_right_out_10_[0]),
		.chanx_in_11_(sb_2__2__0_chanx_left_out_11_[0]),
		.chanx_in_12_(sb_1__2__0_chanx_right_out_12_[0]),
		.chanx_in_13_(sb_2__2__0_chanx_left_out_13_[0]),
		.chanx_in_14_(sb_1__2__0_chanx_right_out_14_[0]),
		.chanx_in_15_(sb_2__2__0_chanx_left_out_15_[0]),
		.chanx_in_16_(sb_1__2__0_chanx_right_out_16_[0]),
		.chanx_in_17_(sb_2__2__0_chanx_left_out_17_[0]),
		.chanx_in_18_(sb_1__2__0_chanx_right_out_18_[0]),
		.chanx_in_19_(sb_2__2__0_chanx_left_out_19_[0]),
		.chanx_in_20_(sb_1__2__0_chanx_right_out_20_[0]),
		.chanx_in_21_(sb_2__2__0_chanx_left_out_21_[0]),
		.chanx_in_22_(sb_1__2__0_chanx_right_out_22_[0]),
		.chanx_in_23_(sb_2__2__0_chanx_left_out_23_[0]),
		.chanx_in_24_(sb_1__2__0_chanx_right_out_24_[0]),
		.chanx_in_25_(sb_2__2__0_chanx_left_out_25_[0]),
		.chanx_in_26_(sb_1__2__0_chanx_right_out_26_[0]),
		.chanx_in_27_(sb_2__2__0_chanx_left_out_27_[0]),
		.chanx_in_28_(sb_1__2__0_chanx_right_out_28_[0]),
		.chanx_in_29_(sb_2__2__0_chanx_left_out_29_[0]),
		.chanx_in_30_(sb_1__2__0_chanx_right_out_30_[0]),
		.chanx_in_31_(sb_2__2__0_chanx_left_out_31_[0]),
		.chanx_in_32_(sb_1__2__0_chanx_right_out_32_[0]),
		.chanx_in_33_(sb_2__2__0_chanx_left_out_33_[0]),
		.chanx_in_34_(sb_1__2__0_chanx_right_out_34_[0]),
		.chanx_in_35_(sb_2__2__0_chanx_left_out_35_[0]),
		.chanx_in_36_(sb_1__2__0_chanx_right_out_36_[0]),
		.chanx_in_37_(sb_2__2__0_chanx_left_out_37_[0]),
		.chanx_in_38_(sb_1__2__0_chanx_right_out_38_[0]),
		.chanx_in_39_(sb_2__2__0_chanx_left_out_39_[0]),
		.chanx_in_40_(sb_1__2__0_chanx_right_out_40_[0]),
		.chanx_in_41_(sb_2__2__0_chanx_left_out_41_[0]),
		.chanx_in_42_(sb_1__2__0_chanx_right_out_42_[0]),
		.chanx_in_43_(sb_2__2__0_chanx_left_out_43_[0]),
		.chanx_in_44_(sb_1__2__0_chanx_right_out_44_[0]),
		.chanx_in_45_(sb_2__2__0_chanx_left_out_45_[0]),
		.chanx_in_46_(sb_1__2__0_chanx_right_out_46_[0]),
		.chanx_in_47_(sb_2__2__0_chanx_left_out_47_[0]),
		.chanx_in_48_(sb_1__2__0_chanx_right_out_48_[0]),
		.chanx_in_49_(sb_2__2__0_chanx_left_out_49_[0]),
		.chanx_in_50_(sb_1__2__0_chanx_right_out_50_[0]),
		.chanx_in_51_(sb_2__2__0_chanx_left_out_51_[0]),
		.chanx_in_52_(sb_1__2__0_chanx_right_out_52_[0]),
		.chanx_in_53_(sb_2__2__0_chanx_left_out_53_[0]),
		.chanx_in_54_(sb_1__2__0_chanx_right_out_54_[0]),
		.chanx_in_55_(sb_2__2__0_chanx_left_out_55_[0]),
		.chanx_in_56_(sb_1__2__0_chanx_right_out_56_[0]),
		.chanx_in_57_(sb_2__2__0_chanx_left_out_57_[0]),
		.chanx_in_58_(sb_1__2__0_chanx_right_out_58_[0]),
		.chanx_in_59_(sb_2__2__0_chanx_left_out_59_[0]),
		.chanx_in_60_(sb_1__2__0_chanx_right_out_60_[0]),
		.chanx_in_61_(sb_2__2__0_chanx_left_out_61_[0]),
		.chanx_in_62_(sb_1__2__0_chanx_right_out_62_[0]),
		.chanx_in_63_(sb_2__2__0_chanx_left_out_63_[0]),
		.chanx_in_64_(sb_1__2__0_chanx_right_out_64_[0]),
		.chanx_in_65_(sb_2__2__0_chanx_left_out_65_[0]),
		.chanx_in_66_(sb_1__2__0_chanx_right_out_66_[0]),
		.chanx_in_67_(sb_2__2__0_chanx_left_out_67_[0]),
		.chanx_in_68_(sb_1__2__0_chanx_right_out_68_[0]),
		.chanx_in_69_(sb_2__2__0_chanx_left_out_69_[0]),
		.chanx_in_70_(sb_1__2__0_chanx_right_out_70_[0]),
		.chanx_in_71_(sb_2__2__0_chanx_left_out_71_[0]),
		.chanx_in_72_(sb_1__2__0_chanx_right_out_72_[0]),
		.chanx_in_73_(sb_2__2__0_chanx_left_out_73_[0]),
		.chanx_in_74_(sb_1__2__0_chanx_right_out_74_[0]),
		.chanx_in_75_(sb_2__2__0_chanx_left_out_75_[0]),
		.chanx_in_76_(sb_1__2__0_chanx_right_out_76_[0]),
		.chanx_in_77_(sb_2__2__0_chanx_left_out_77_[0]),
		.chanx_in_78_(sb_1__2__0_chanx_right_out_78_[0]),
		.chanx_in_79_(sb_2__2__0_chanx_left_out_79_[0]),
		.chanx_in_80_(sb_1__2__0_chanx_right_out_80_[0]),
		.chanx_in_81_(sb_2__2__0_chanx_left_out_81_[0]),
		.chanx_in_82_(sb_1__2__0_chanx_right_out_82_[0]),
		.chanx_in_83_(sb_2__2__0_chanx_left_out_83_[0]),
		.chanx_in_84_(sb_1__2__0_chanx_right_out_84_[0]),
		.chanx_in_85_(sb_2__2__0_chanx_left_out_85_[0]),
		.chanx_in_86_(sb_1__2__0_chanx_right_out_86_[0]),
		.chanx_in_87_(sb_2__2__0_chanx_left_out_87_[0]),
		.chanx_in_88_(sb_1__2__0_chanx_right_out_88_[0]),
		.chanx_in_89_(sb_2__2__0_chanx_left_out_89_[0]),
		.chanx_in_90_(sb_1__2__0_chanx_right_out_90_[0]),
		.chanx_in_91_(sb_2__2__0_chanx_left_out_91_[0]),
		.chanx_in_92_(sb_1__2__0_chanx_right_out_92_[0]),
		.chanx_in_93_(sb_2__2__0_chanx_left_out_93_[0]),
		.chanx_in_94_(sb_1__2__0_chanx_right_out_94_[0]),
		.chanx_in_95_(sb_2__2__0_chanx_left_out_95_[0]),
		.chanx_in_96_(sb_1__2__0_chanx_right_out_96_[0]),
		.chanx_in_97_(sb_2__2__0_chanx_left_out_97_[0]),
		.chanx_in_98_(sb_1__2__0_chanx_right_out_98_[0]),
		.chanx_in_99_(sb_2__2__0_chanx_left_out_99_[0]),
		.chanx_in_100_(sb_1__2__0_chanx_right_out_100_[0]),
		.chanx_in_101_(sb_2__2__0_chanx_left_out_101_[0]),
		.chanx_in_102_(sb_1__2__0_chanx_right_out_102_[0]),
		.chanx_in_103_(sb_2__2__0_chanx_left_out_103_[0]),
		.chanx_in_104_(sb_1__2__0_chanx_right_out_104_[0]),
		.chanx_in_105_(sb_2__2__0_chanx_left_out_105_[0]),
		.chanx_in_106_(sb_1__2__0_chanx_right_out_106_[0]),
		.chanx_in_107_(sb_2__2__0_chanx_left_out_107_[0]),
		.chanx_in_108_(sb_1__2__0_chanx_right_out_108_[0]),
		.chanx_in_109_(sb_2__2__0_chanx_left_out_109_[0]),
		.chanx_in_110_(sb_1__2__0_chanx_right_out_110_[0]),
		.chanx_in_111_(sb_2__2__0_chanx_left_out_111_[0]),
		.chanx_in_112_(sb_1__2__0_chanx_right_out_112_[0]),
		.chanx_in_113_(sb_2__2__0_chanx_left_out_113_[0]),
		.chanx_in_114_(sb_1__2__0_chanx_right_out_114_[0]),
		.chanx_in_115_(sb_2__2__0_chanx_left_out_115_[0]),
		.chanx_in_116_(sb_1__2__0_chanx_right_out_116_[0]),
		.chanx_in_117_(sb_2__2__0_chanx_left_out_117_[0]),
		.chanx_in_118_(sb_1__2__0_chanx_right_out_118_[0]),
		.chanx_in_119_(sb_2__2__0_chanx_left_out_119_[0]),
		.chanx_in_120_(sb_1__2__0_chanx_right_out_120_[0]),
		.chanx_in_121_(sb_2__2__0_chanx_left_out_121_[0]),
		.chanx_in_122_(sb_1__2__0_chanx_right_out_122_[0]),
		.chanx_in_123_(sb_2__2__0_chanx_left_out_123_[0]),
		.chanx_in_124_(sb_1__2__0_chanx_right_out_124_[0]),
		.chanx_in_125_(sb_2__2__0_chanx_left_out_125_[0]),
		.chanx_in_126_(sb_1__2__0_chanx_right_out_126_[0]),
		.chanx_in_127_(sb_2__2__0_chanx_left_out_127_[0]),
		.chanx_in_128_(sb_1__2__0_chanx_right_out_128_[0]),
		.chanx_in_129_(sb_2__2__0_chanx_left_out_129_[0]),
		.chanx_in_130_(sb_1__2__0_chanx_right_out_130_[0]),
		.chanx_in_131_(sb_2__2__0_chanx_left_out_131_[0]),
		.chanx_in_132_(sb_1__2__0_chanx_right_out_132_[0]),
		.chanx_in_133_(sb_2__2__0_chanx_left_out_133_[0]),
		.chanx_in_134_(sb_1__2__0_chanx_right_out_134_[0]),
		.chanx_in_135_(sb_2__2__0_chanx_left_out_135_[0]),
		.chanx_in_136_(sb_1__2__0_chanx_right_out_136_[0]),
		.chanx_in_137_(sb_2__2__0_chanx_left_out_137_[0]),
		.chanx_in_138_(sb_1__2__0_chanx_right_out_138_[0]),
		.chanx_in_139_(sb_2__2__0_chanx_left_out_139_[0]),
		.chanx_in_140_(sb_1__2__0_chanx_right_out_140_[0]),
		.chanx_in_141_(sb_2__2__0_chanx_left_out_141_[0]),
		.chanx_in_142_(sb_1__2__0_chanx_right_out_142_[0]),
		.chanx_in_143_(sb_2__2__0_chanx_left_out_143_[0]),
		.chanx_in_144_(sb_1__2__0_chanx_right_out_144_[0]),
		.chanx_in_145_(sb_2__2__0_chanx_left_out_145_[0]),
		.chanx_in_146_(sb_1__2__0_chanx_right_out_146_[0]),
		.chanx_in_147_(sb_2__2__0_chanx_left_out_147_[0]),
		.chanx_in_148_(sb_1__2__0_chanx_right_out_148_[0]),
		.chanx_in_149_(sb_2__2__0_chanx_left_out_149_[0]),
		.chanx_in_150_(sb_1__2__0_chanx_right_out_150_[0]),
		.chanx_in_151_(sb_2__2__0_chanx_left_out_151_[0]),
		.chanx_in_152_(sb_1__2__0_chanx_right_out_152_[0]),
		.chanx_in_153_(sb_2__2__0_chanx_left_out_153_[0]),
		.chanx_in_154_(sb_1__2__0_chanx_right_out_154_[0]),
		.chanx_in_155_(sb_2__2__0_chanx_left_out_155_[0]),
		.chanx_in_156_(sb_1__2__0_chanx_right_out_156_[0]),
		.chanx_in_157_(sb_2__2__0_chanx_left_out_157_[0]),
		.chanx_in_158_(sb_1__2__0_chanx_right_out_158_[0]),
		.chanx_in_159_(sb_2__2__0_chanx_left_out_159_[0]),
		.chanx_in_160_(sb_1__2__0_chanx_right_out_160_[0]),
		.chanx_in_161_(sb_2__2__0_chanx_left_out_161_[0]),
		.chanx_in_162_(sb_1__2__0_chanx_right_out_162_[0]),
		.chanx_in_163_(sb_2__2__0_chanx_left_out_163_[0]),
		.chanx_in_164_(sb_1__2__0_chanx_right_out_164_[0]),
		.chanx_in_165_(sb_2__2__0_chanx_left_out_165_[0]),
		.chanx_in_166_(sb_1__2__0_chanx_right_out_166_[0]),
		.chanx_in_167_(sb_2__2__0_chanx_left_out_167_[0]),
		.chanx_in_168_(sb_1__2__0_chanx_right_out_168_[0]),
		.chanx_in_169_(sb_2__2__0_chanx_left_out_169_[0]),
		.chanx_in_170_(sb_1__2__0_chanx_right_out_170_[0]),
		.chanx_in_171_(sb_2__2__0_chanx_left_out_171_[0]),
		.chanx_in_172_(sb_1__2__0_chanx_right_out_172_[0]),
		.chanx_in_173_(sb_2__2__0_chanx_left_out_173_[0]),
		.chanx_in_174_(sb_1__2__0_chanx_right_out_174_[0]),
		.chanx_in_175_(sb_2__2__0_chanx_left_out_175_[0]),
		.chanx_in_176_(sb_1__2__0_chanx_right_out_176_[0]),
		.chanx_in_177_(sb_2__2__0_chanx_left_out_177_[0]),
		.chanx_in_178_(sb_1__2__0_chanx_right_out_178_[0]),
		.chanx_in_179_(sb_2__2__0_chanx_left_out_179_[0]),
		.chanx_in_180_(sb_1__2__0_chanx_right_out_180_[0]),
		.chanx_in_181_(sb_2__2__0_chanx_left_out_181_[0]),
		.chanx_in_182_(sb_1__2__0_chanx_right_out_182_[0]),
		.chanx_in_183_(sb_2__2__0_chanx_left_out_183_[0]),
		.chanx_in_184_(sb_1__2__0_chanx_right_out_184_[0]),
		.chanx_in_185_(sb_2__2__0_chanx_left_out_185_[0]),
		.chanx_in_186_(sb_1__2__0_chanx_right_out_186_[0]),
		.chanx_in_187_(sb_2__2__0_chanx_left_out_187_[0]),
		.chanx_in_188_(sb_1__2__0_chanx_right_out_188_[0]),
		.chanx_in_189_(sb_2__2__0_chanx_left_out_189_[0]),
		.chanx_in_190_(sb_1__2__0_chanx_right_out_190_[0]),
		.chanx_in_191_(sb_2__2__0_chanx_left_out_191_[0]),
		.chanx_in_192_(sb_1__2__0_chanx_right_out_192_[0]),
		.chanx_in_193_(sb_2__2__0_chanx_left_out_193_[0]),
		.chanx_in_194_(sb_1__2__0_chanx_right_out_194_[0]),
		.chanx_in_195_(sb_2__2__0_chanx_left_out_195_[0]),
		.chanx_in_196_(sb_1__2__0_chanx_right_out_196_[0]),
		.chanx_in_197_(sb_2__2__0_chanx_left_out_197_[0]),
		.chanx_in_198_(sb_1__2__0_chanx_right_out_198_[0]),
		.chanx_in_199_(sb_2__2__0_chanx_left_out_199_[0]),
		.ccff_head(sb_2__2__0_ccff_tail[0]),
		.chanx_out_0_(cbx_1__2__1_chanx_out_0_[0]),
		.chanx_out_1_(cbx_1__2__1_chanx_out_1_[0]),
		.chanx_out_2_(cbx_1__2__1_chanx_out_2_[0]),
		.chanx_out_3_(cbx_1__2__1_chanx_out_3_[0]),
		.chanx_out_4_(cbx_1__2__1_chanx_out_4_[0]),
		.chanx_out_5_(cbx_1__2__1_chanx_out_5_[0]),
		.chanx_out_6_(cbx_1__2__1_chanx_out_6_[0]),
		.chanx_out_7_(cbx_1__2__1_chanx_out_7_[0]),
		.chanx_out_8_(cbx_1__2__1_chanx_out_8_[0]),
		.chanx_out_9_(cbx_1__2__1_chanx_out_9_[0]),
		.chanx_out_10_(cbx_1__2__1_chanx_out_10_[0]),
		.chanx_out_11_(cbx_1__2__1_chanx_out_11_[0]),
		.chanx_out_12_(cbx_1__2__1_chanx_out_12_[0]),
		.chanx_out_13_(cbx_1__2__1_chanx_out_13_[0]),
		.chanx_out_14_(cbx_1__2__1_chanx_out_14_[0]),
		.chanx_out_15_(cbx_1__2__1_chanx_out_15_[0]),
		.chanx_out_16_(cbx_1__2__1_chanx_out_16_[0]),
		.chanx_out_17_(cbx_1__2__1_chanx_out_17_[0]),
		.chanx_out_18_(cbx_1__2__1_chanx_out_18_[0]),
		.chanx_out_19_(cbx_1__2__1_chanx_out_19_[0]),
		.chanx_out_20_(cbx_1__2__1_chanx_out_20_[0]),
		.chanx_out_21_(cbx_1__2__1_chanx_out_21_[0]),
		.chanx_out_22_(cbx_1__2__1_chanx_out_22_[0]),
		.chanx_out_23_(cbx_1__2__1_chanx_out_23_[0]),
		.chanx_out_24_(cbx_1__2__1_chanx_out_24_[0]),
		.chanx_out_25_(cbx_1__2__1_chanx_out_25_[0]),
		.chanx_out_26_(cbx_1__2__1_chanx_out_26_[0]),
		.chanx_out_27_(cbx_1__2__1_chanx_out_27_[0]),
		.chanx_out_28_(cbx_1__2__1_chanx_out_28_[0]),
		.chanx_out_29_(cbx_1__2__1_chanx_out_29_[0]),
		.chanx_out_30_(cbx_1__2__1_chanx_out_30_[0]),
		.chanx_out_31_(cbx_1__2__1_chanx_out_31_[0]),
		.chanx_out_32_(cbx_1__2__1_chanx_out_32_[0]),
		.chanx_out_33_(cbx_1__2__1_chanx_out_33_[0]),
		.chanx_out_34_(cbx_1__2__1_chanx_out_34_[0]),
		.chanx_out_35_(cbx_1__2__1_chanx_out_35_[0]),
		.chanx_out_36_(cbx_1__2__1_chanx_out_36_[0]),
		.chanx_out_37_(cbx_1__2__1_chanx_out_37_[0]),
		.chanx_out_38_(cbx_1__2__1_chanx_out_38_[0]),
		.chanx_out_39_(cbx_1__2__1_chanx_out_39_[0]),
		.chanx_out_40_(cbx_1__2__1_chanx_out_40_[0]),
		.chanx_out_41_(cbx_1__2__1_chanx_out_41_[0]),
		.chanx_out_42_(cbx_1__2__1_chanx_out_42_[0]),
		.chanx_out_43_(cbx_1__2__1_chanx_out_43_[0]),
		.chanx_out_44_(cbx_1__2__1_chanx_out_44_[0]),
		.chanx_out_45_(cbx_1__2__1_chanx_out_45_[0]),
		.chanx_out_46_(cbx_1__2__1_chanx_out_46_[0]),
		.chanx_out_47_(cbx_1__2__1_chanx_out_47_[0]),
		.chanx_out_48_(cbx_1__2__1_chanx_out_48_[0]),
		.chanx_out_49_(cbx_1__2__1_chanx_out_49_[0]),
		.chanx_out_50_(cbx_1__2__1_chanx_out_50_[0]),
		.chanx_out_51_(cbx_1__2__1_chanx_out_51_[0]),
		.chanx_out_52_(cbx_1__2__1_chanx_out_52_[0]),
		.chanx_out_53_(cbx_1__2__1_chanx_out_53_[0]),
		.chanx_out_54_(cbx_1__2__1_chanx_out_54_[0]),
		.chanx_out_55_(cbx_1__2__1_chanx_out_55_[0]),
		.chanx_out_56_(cbx_1__2__1_chanx_out_56_[0]),
		.chanx_out_57_(cbx_1__2__1_chanx_out_57_[0]),
		.chanx_out_58_(cbx_1__2__1_chanx_out_58_[0]),
		.chanx_out_59_(cbx_1__2__1_chanx_out_59_[0]),
		.chanx_out_60_(cbx_1__2__1_chanx_out_60_[0]),
		.chanx_out_61_(cbx_1__2__1_chanx_out_61_[0]),
		.chanx_out_62_(cbx_1__2__1_chanx_out_62_[0]),
		.chanx_out_63_(cbx_1__2__1_chanx_out_63_[0]),
		.chanx_out_64_(cbx_1__2__1_chanx_out_64_[0]),
		.chanx_out_65_(cbx_1__2__1_chanx_out_65_[0]),
		.chanx_out_66_(cbx_1__2__1_chanx_out_66_[0]),
		.chanx_out_67_(cbx_1__2__1_chanx_out_67_[0]),
		.chanx_out_68_(cbx_1__2__1_chanx_out_68_[0]),
		.chanx_out_69_(cbx_1__2__1_chanx_out_69_[0]),
		.chanx_out_70_(cbx_1__2__1_chanx_out_70_[0]),
		.chanx_out_71_(cbx_1__2__1_chanx_out_71_[0]),
		.chanx_out_72_(cbx_1__2__1_chanx_out_72_[0]),
		.chanx_out_73_(cbx_1__2__1_chanx_out_73_[0]),
		.chanx_out_74_(cbx_1__2__1_chanx_out_74_[0]),
		.chanx_out_75_(cbx_1__2__1_chanx_out_75_[0]),
		.chanx_out_76_(cbx_1__2__1_chanx_out_76_[0]),
		.chanx_out_77_(cbx_1__2__1_chanx_out_77_[0]),
		.chanx_out_78_(cbx_1__2__1_chanx_out_78_[0]),
		.chanx_out_79_(cbx_1__2__1_chanx_out_79_[0]),
		.chanx_out_80_(cbx_1__2__1_chanx_out_80_[0]),
		.chanx_out_81_(cbx_1__2__1_chanx_out_81_[0]),
		.chanx_out_82_(cbx_1__2__1_chanx_out_82_[0]),
		.chanx_out_83_(cbx_1__2__1_chanx_out_83_[0]),
		.chanx_out_84_(cbx_1__2__1_chanx_out_84_[0]),
		.chanx_out_85_(cbx_1__2__1_chanx_out_85_[0]),
		.chanx_out_86_(cbx_1__2__1_chanx_out_86_[0]),
		.chanx_out_87_(cbx_1__2__1_chanx_out_87_[0]),
		.chanx_out_88_(cbx_1__2__1_chanx_out_88_[0]),
		.chanx_out_89_(cbx_1__2__1_chanx_out_89_[0]),
		.chanx_out_90_(cbx_1__2__1_chanx_out_90_[0]),
		.chanx_out_91_(cbx_1__2__1_chanx_out_91_[0]),
		.chanx_out_92_(cbx_1__2__1_chanx_out_92_[0]),
		.chanx_out_93_(cbx_1__2__1_chanx_out_93_[0]),
		.chanx_out_94_(cbx_1__2__1_chanx_out_94_[0]),
		.chanx_out_95_(cbx_1__2__1_chanx_out_95_[0]),
		.chanx_out_96_(cbx_1__2__1_chanx_out_96_[0]),
		.chanx_out_97_(cbx_1__2__1_chanx_out_97_[0]),
		.chanx_out_98_(cbx_1__2__1_chanx_out_98_[0]),
		.chanx_out_99_(cbx_1__2__1_chanx_out_99_[0]),
		.chanx_out_100_(cbx_1__2__1_chanx_out_100_[0]),
		.chanx_out_101_(cbx_1__2__1_chanx_out_101_[0]),
		.chanx_out_102_(cbx_1__2__1_chanx_out_102_[0]),
		.chanx_out_103_(cbx_1__2__1_chanx_out_103_[0]),
		.chanx_out_104_(cbx_1__2__1_chanx_out_104_[0]),
		.chanx_out_105_(cbx_1__2__1_chanx_out_105_[0]),
		.chanx_out_106_(cbx_1__2__1_chanx_out_106_[0]),
		.chanx_out_107_(cbx_1__2__1_chanx_out_107_[0]),
		.chanx_out_108_(cbx_1__2__1_chanx_out_108_[0]),
		.chanx_out_109_(cbx_1__2__1_chanx_out_109_[0]),
		.chanx_out_110_(cbx_1__2__1_chanx_out_110_[0]),
		.chanx_out_111_(cbx_1__2__1_chanx_out_111_[0]),
		.chanx_out_112_(cbx_1__2__1_chanx_out_112_[0]),
		.chanx_out_113_(cbx_1__2__1_chanx_out_113_[0]),
		.chanx_out_114_(cbx_1__2__1_chanx_out_114_[0]),
		.chanx_out_115_(cbx_1__2__1_chanx_out_115_[0]),
		.chanx_out_116_(cbx_1__2__1_chanx_out_116_[0]),
		.chanx_out_117_(cbx_1__2__1_chanx_out_117_[0]),
		.chanx_out_118_(cbx_1__2__1_chanx_out_118_[0]),
		.chanx_out_119_(cbx_1__2__1_chanx_out_119_[0]),
		.chanx_out_120_(cbx_1__2__1_chanx_out_120_[0]),
		.chanx_out_121_(cbx_1__2__1_chanx_out_121_[0]),
		.chanx_out_122_(cbx_1__2__1_chanx_out_122_[0]),
		.chanx_out_123_(cbx_1__2__1_chanx_out_123_[0]),
		.chanx_out_124_(cbx_1__2__1_chanx_out_124_[0]),
		.chanx_out_125_(cbx_1__2__1_chanx_out_125_[0]),
		.chanx_out_126_(cbx_1__2__1_chanx_out_126_[0]),
		.chanx_out_127_(cbx_1__2__1_chanx_out_127_[0]),
		.chanx_out_128_(cbx_1__2__1_chanx_out_128_[0]),
		.chanx_out_129_(cbx_1__2__1_chanx_out_129_[0]),
		.chanx_out_130_(cbx_1__2__1_chanx_out_130_[0]),
		.chanx_out_131_(cbx_1__2__1_chanx_out_131_[0]),
		.chanx_out_132_(cbx_1__2__1_chanx_out_132_[0]),
		.chanx_out_133_(cbx_1__2__1_chanx_out_133_[0]),
		.chanx_out_134_(cbx_1__2__1_chanx_out_134_[0]),
		.chanx_out_135_(cbx_1__2__1_chanx_out_135_[0]),
		.chanx_out_136_(cbx_1__2__1_chanx_out_136_[0]),
		.chanx_out_137_(cbx_1__2__1_chanx_out_137_[0]),
		.chanx_out_138_(cbx_1__2__1_chanx_out_138_[0]),
		.chanx_out_139_(cbx_1__2__1_chanx_out_139_[0]),
		.chanx_out_140_(cbx_1__2__1_chanx_out_140_[0]),
		.chanx_out_141_(cbx_1__2__1_chanx_out_141_[0]),
		.chanx_out_142_(cbx_1__2__1_chanx_out_142_[0]),
		.chanx_out_143_(cbx_1__2__1_chanx_out_143_[0]),
		.chanx_out_144_(cbx_1__2__1_chanx_out_144_[0]),
		.chanx_out_145_(cbx_1__2__1_chanx_out_145_[0]),
		.chanx_out_146_(cbx_1__2__1_chanx_out_146_[0]),
		.chanx_out_147_(cbx_1__2__1_chanx_out_147_[0]),
		.chanx_out_148_(cbx_1__2__1_chanx_out_148_[0]),
		.chanx_out_149_(cbx_1__2__1_chanx_out_149_[0]),
		.chanx_out_150_(cbx_1__2__1_chanx_out_150_[0]),
		.chanx_out_151_(cbx_1__2__1_chanx_out_151_[0]),
		.chanx_out_152_(cbx_1__2__1_chanx_out_152_[0]),
		.chanx_out_153_(cbx_1__2__1_chanx_out_153_[0]),
		.chanx_out_154_(cbx_1__2__1_chanx_out_154_[0]),
		.chanx_out_155_(cbx_1__2__1_chanx_out_155_[0]),
		.chanx_out_156_(cbx_1__2__1_chanx_out_156_[0]),
		.chanx_out_157_(cbx_1__2__1_chanx_out_157_[0]),
		.chanx_out_158_(cbx_1__2__1_chanx_out_158_[0]),
		.chanx_out_159_(cbx_1__2__1_chanx_out_159_[0]),
		.chanx_out_160_(cbx_1__2__1_chanx_out_160_[0]),
		.chanx_out_161_(cbx_1__2__1_chanx_out_161_[0]),
		.chanx_out_162_(cbx_1__2__1_chanx_out_162_[0]),
		.chanx_out_163_(cbx_1__2__1_chanx_out_163_[0]),
		.chanx_out_164_(cbx_1__2__1_chanx_out_164_[0]),
		.chanx_out_165_(cbx_1__2__1_chanx_out_165_[0]),
		.chanx_out_166_(cbx_1__2__1_chanx_out_166_[0]),
		.chanx_out_167_(cbx_1__2__1_chanx_out_167_[0]),
		.chanx_out_168_(cbx_1__2__1_chanx_out_168_[0]),
		.chanx_out_169_(cbx_1__2__1_chanx_out_169_[0]),
		.chanx_out_170_(cbx_1__2__1_chanx_out_170_[0]),
		.chanx_out_171_(cbx_1__2__1_chanx_out_171_[0]),
		.chanx_out_172_(cbx_1__2__1_chanx_out_172_[0]),
		.chanx_out_173_(cbx_1__2__1_chanx_out_173_[0]),
		.chanx_out_174_(cbx_1__2__1_chanx_out_174_[0]),
		.chanx_out_175_(cbx_1__2__1_chanx_out_175_[0]),
		.chanx_out_176_(cbx_1__2__1_chanx_out_176_[0]),
		.chanx_out_177_(cbx_1__2__1_chanx_out_177_[0]),
		.chanx_out_178_(cbx_1__2__1_chanx_out_178_[0]),
		.chanx_out_179_(cbx_1__2__1_chanx_out_179_[0]),
		.chanx_out_180_(cbx_1__2__1_chanx_out_180_[0]),
		.chanx_out_181_(cbx_1__2__1_chanx_out_181_[0]),
		.chanx_out_182_(cbx_1__2__1_chanx_out_182_[0]),
		.chanx_out_183_(cbx_1__2__1_chanx_out_183_[0]),
		.chanx_out_184_(cbx_1__2__1_chanx_out_184_[0]),
		.chanx_out_185_(cbx_1__2__1_chanx_out_185_[0]),
		.chanx_out_186_(cbx_1__2__1_chanx_out_186_[0]),
		.chanx_out_187_(cbx_1__2__1_chanx_out_187_[0]),
		.chanx_out_188_(cbx_1__2__1_chanx_out_188_[0]),
		.chanx_out_189_(cbx_1__2__1_chanx_out_189_[0]),
		.chanx_out_190_(cbx_1__2__1_chanx_out_190_[0]),
		.chanx_out_191_(cbx_1__2__1_chanx_out_191_[0]),
		.chanx_out_192_(cbx_1__2__1_chanx_out_192_[0]),
		.chanx_out_193_(cbx_1__2__1_chanx_out_193_[0]),
		.chanx_out_194_(cbx_1__2__1_chanx_out_194_[0]),
		.chanx_out_195_(cbx_1__2__1_chanx_out_195_[0]),
		.chanx_out_196_(cbx_1__2__1_chanx_out_196_[0]),
		.chanx_out_197_(cbx_1__2__1_chanx_out_197_[0]),
		.chanx_out_198_(cbx_1__2__1_chanx_out_198_[0]),
		.chanx_out_199_(cbx_1__2__1_chanx_out_199_[0]),
		.top_grid_pin_0_(cbx_1__2__1_top_grid_pin_0_[0]),
		.bottom_grid_pin_42_(cbx_1__2__1_bottom_grid_pin_42_[0]),
		.bottom_grid_pin_43_(cbx_1__2__1_bottom_grid_pin_43_[0]),
		.bottom_grid_pin_68_(cbx_1__2__1_bottom_grid_pin_68_[0]),
		.ccff_tail(cbx_1__2__1_ccff_tail[0]));

	cby_0__1_ cby_0__1_ (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.chany_in_0_(sb_0__0__0_chany_top_out_0_[0]),
		.chany_in_1_(sb_0__1__0_chany_bottom_out_1_[0]),
		.chany_in_2_(sb_0__0__0_chany_top_out_2_[0]),
		.chany_in_3_(sb_0__1__0_chany_bottom_out_3_[0]),
		.chany_in_4_(sb_0__0__0_chany_top_out_4_[0]),
		.chany_in_5_(sb_0__1__0_chany_bottom_out_5_[0]),
		.chany_in_6_(sb_0__0__0_chany_top_out_6_[0]),
		.chany_in_7_(sb_0__1__0_chany_bottom_out_7_[0]),
		.chany_in_8_(sb_0__0__0_chany_top_out_8_[0]),
		.chany_in_9_(sb_0__1__0_chany_bottom_out_9_[0]),
		.chany_in_10_(sb_0__0__0_chany_top_out_10_[0]),
		.chany_in_11_(sb_0__1__0_chany_bottom_out_11_[0]),
		.chany_in_12_(sb_0__0__0_chany_top_out_12_[0]),
		.chany_in_13_(sb_0__1__0_chany_bottom_out_13_[0]),
		.chany_in_14_(sb_0__0__0_chany_top_out_14_[0]),
		.chany_in_15_(sb_0__1__0_chany_bottom_out_15_[0]),
		.chany_in_16_(sb_0__0__0_chany_top_out_16_[0]),
		.chany_in_17_(sb_0__1__0_chany_bottom_out_17_[0]),
		.chany_in_18_(sb_0__0__0_chany_top_out_18_[0]),
		.chany_in_19_(sb_0__1__0_chany_bottom_out_19_[0]),
		.chany_in_20_(sb_0__0__0_chany_top_out_20_[0]),
		.chany_in_21_(sb_0__1__0_chany_bottom_out_21_[0]),
		.chany_in_22_(sb_0__0__0_chany_top_out_22_[0]),
		.chany_in_23_(sb_0__1__0_chany_bottom_out_23_[0]),
		.chany_in_24_(sb_0__0__0_chany_top_out_24_[0]),
		.chany_in_25_(sb_0__1__0_chany_bottom_out_25_[0]),
		.chany_in_26_(sb_0__0__0_chany_top_out_26_[0]),
		.chany_in_27_(sb_0__1__0_chany_bottom_out_27_[0]),
		.chany_in_28_(sb_0__0__0_chany_top_out_28_[0]),
		.chany_in_29_(sb_0__1__0_chany_bottom_out_29_[0]),
		.chany_in_30_(sb_0__0__0_chany_top_out_30_[0]),
		.chany_in_31_(sb_0__1__0_chany_bottom_out_31_[0]),
		.chany_in_32_(sb_0__0__0_chany_top_out_32_[0]),
		.chany_in_33_(sb_0__1__0_chany_bottom_out_33_[0]),
		.chany_in_34_(sb_0__0__0_chany_top_out_34_[0]),
		.chany_in_35_(sb_0__1__0_chany_bottom_out_35_[0]),
		.chany_in_36_(sb_0__0__0_chany_top_out_36_[0]),
		.chany_in_37_(sb_0__1__0_chany_bottom_out_37_[0]),
		.chany_in_38_(sb_0__0__0_chany_top_out_38_[0]),
		.chany_in_39_(sb_0__1__0_chany_bottom_out_39_[0]),
		.chany_in_40_(sb_0__0__0_chany_top_out_40_[0]),
		.chany_in_41_(sb_0__1__0_chany_bottom_out_41_[0]),
		.chany_in_42_(sb_0__0__0_chany_top_out_42_[0]),
		.chany_in_43_(sb_0__1__0_chany_bottom_out_43_[0]),
		.chany_in_44_(sb_0__0__0_chany_top_out_44_[0]),
		.chany_in_45_(sb_0__1__0_chany_bottom_out_45_[0]),
		.chany_in_46_(sb_0__0__0_chany_top_out_46_[0]),
		.chany_in_47_(sb_0__1__0_chany_bottom_out_47_[0]),
		.chany_in_48_(sb_0__0__0_chany_top_out_48_[0]),
		.chany_in_49_(sb_0__1__0_chany_bottom_out_49_[0]),
		.chany_in_50_(sb_0__0__0_chany_top_out_50_[0]),
		.chany_in_51_(sb_0__1__0_chany_bottom_out_51_[0]),
		.chany_in_52_(sb_0__0__0_chany_top_out_52_[0]),
		.chany_in_53_(sb_0__1__0_chany_bottom_out_53_[0]),
		.chany_in_54_(sb_0__0__0_chany_top_out_54_[0]),
		.chany_in_55_(sb_0__1__0_chany_bottom_out_55_[0]),
		.chany_in_56_(sb_0__0__0_chany_top_out_56_[0]),
		.chany_in_57_(sb_0__1__0_chany_bottom_out_57_[0]),
		.chany_in_58_(sb_0__0__0_chany_top_out_58_[0]),
		.chany_in_59_(sb_0__1__0_chany_bottom_out_59_[0]),
		.chany_in_60_(sb_0__0__0_chany_top_out_60_[0]),
		.chany_in_61_(sb_0__1__0_chany_bottom_out_61_[0]),
		.chany_in_62_(sb_0__0__0_chany_top_out_62_[0]),
		.chany_in_63_(sb_0__1__0_chany_bottom_out_63_[0]),
		.chany_in_64_(sb_0__0__0_chany_top_out_64_[0]),
		.chany_in_65_(sb_0__1__0_chany_bottom_out_65_[0]),
		.chany_in_66_(sb_0__0__0_chany_top_out_66_[0]),
		.chany_in_67_(sb_0__1__0_chany_bottom_out_67_[0]),
		.chany_in_68_(sb_0__0__0_chany_top_out_68_[0]),
		.chany_in_69_(sb_0__1__0_chany_bottom_out_69_[0]),
		.chany_in_70_(sb_0__0__0_chany_top_out_70_[0]),
		.chany_in_71_(sb_0__1__0_chany_bottom_out_71_[0]),
		.chany_in_72_(sb_0__0__0_chany_top_out_72_[0]),
		.chany_in_73_(sb_0__1__0_chany_bottom_out_73_[0]),
		.chany_in_74_(sb_0__0__0_chany_top_out_74_[0]),
		.chany_in_75_(sb_0__1__0_chany_bottom_out_75_[0]),
		.chany_in_76_(sb_0__0__0_chany_top_out_76_[0]),
		.chany_in_77_(sb_0__1__0_chany_bottom_out_77_[0]),
		.chany_in_78_(sb_0__0__0_chany_top_out_78_[0]),
		.chany_in_79_(sb_0__1__0_chany_bottom_out_79_[0]),
		.chany_in_80_(sb_0__0__0_chany_top_out_80_[0]),
		.chany_in_81_(sb_0__1__0_chany_bottom_out_81_[0]),
		.chany_in_82_(sb_0__0__0_chany_top_out_82_[0]),
		.chany_in_83_(sb_0__1__0_chany_bottom_out_83_[0]),
		.chany_in_84_(sb_0__0__0_chany_top_out_84_[0]),
		.chany_in_85_(sb_0__1__0_chany_bottom_out_85_[0]),
		.chany_in_86_(sb_0__0__0_chany_top_out_86_[0]),
		.chany_in_87_(sb_0__1__0_chany_bottom_out_87_[0]),
		.chany_in_88_(sb_0__0__0_chany_top_out_88_[0]),
		.chany_in_89_(sb_0__1__0_chany_bottom_out_89_[0]),
		.chany_in_90_(sb_0__0__0_chany_top_out_90_[0]),
		.chany_in_91_(sb_0__1__0_chany_bottom_out_91_[0]),
		.chany_in_92_(sb_0__0__0_chany_top_out_92_[0]),
		.chany_in_93_(sb_0__1__0_chany_bottom_out_93_[0]),
		.chany_in_94_(sb_0__0__0_chany_top_out_94_[0]),
		.chany_in_95_(sb_0__1__0_chany_bottom_out_95_[0]),
		.chany_in_96_(sb_0__0__0_chany_top_out_96_[0]),
		.chany_in_97_(sb_0__1__0_chany_bottom_out_97_[0]),
		.chany_in_98_(sb_0__0__0_chany_top_out_98_[0]),
		.chany_in_99_(sb_0__1__0_chany_bottom_out_99_[0]),
		.chany_in_100_(sb_0__0__0_chany_top_out_100_[0]),
		.chany_in_101_(sb_0__1__0_chany_bottom_out_101_[0]),
		.chany_in_102_(sb_0__0__0_chany_top_out_102_[0]),
		.chany_in_103_(sb_0__1__0_chany_bottom_out_103_[0]),
		.chany_in_104_(sb_0__0__0_chany_top_out_104_[0]),
		.chany_in_105_(sb_0__1__0_chany_bottom_out_105_[0]),
		.chany_in_106_(sb_0__0__0_chany_top_out_106_[0]),
		.chany_in_107_(sb_0__1__0_chany_bottom_out_107_[0]),
		.chany_in_108_(sb_0__0__0_chany_top_out_108_[0]),
		.chany_in_109_(sb_0__1__0_chany_bottom_out_109_[0]),
		.chany_in_110_(sb_0__0__0_chany_top_out_110_[0]),
		.chany_in_111_(sb_0__1__0_chany_bottom_out_111_[0]),
		.chany_in_112_(sb_0__0__0_chany_top_out_112_[0]),
		.chany_in_113_(sb_0__1__0_chany_bottom_out_113_[0]),
		.chany_in_114_(sb_0__0__0_chany_top_out_114_[0]),
		.chany_in_115_(sb_0__1__0_chany_bottom_out_115_[0]),
		.chany_in_116_(sb_0__0__0_chany_top_out_116_[0]),
		.chany_in_117_(sb_0__1__0_chany_bottom_out_117_[0]),
		.chany_in_118_(sb_0__0__0_chany_top_out_118_[0]),
		.chany_in_119_(sb_0__1__0_chany_bottom_out_119_[0]),
		.chany_in_120_(sb_0__0__0_chany_top_out_120_[0]),
		.chany_in_121_(sb_0__1__0_chany_bottom_out_121_[0]),
		.chany_in_122_(sb_0__0__0_chany_top_out_122_[0]),
		.chany_in_123_(sb_0__1__0_chany_bottom_out_123_[0]),
		.chany_in_124_(sb_0__0__0_chany_top_out_124_[0]),
		.chany_in_125_(sb_0__1__0_chany_bottom_out_125_[0]),
		.chany_in_126_(sb_0__0__0_chany_top_out_126_[0]),
		.chany_in_127_(sb_0__1__0_chany_bottom_out_127_[0]),
		.chany_in_128_(sb_0__0__0_chany_top_out_128_[0]),
		.chany_in_129_(sb_0__1__0_chany_bottom_out_129_[0]),
		.chany_in_130_(sb_0__0__0_chany_top_out_130_[0]),
		.chany_in_131_(sb_0__1__0_chany_bottom_out_131_[0]),
		.chany_in_132_(sb_0__0__0_chany_top_out_132_[0]),
		.chany_in_133_(sb_0__1__0_chany_bottom_out_133_[0]),
		.chany_in_134_(sb_0__0__0_chany_top_out_134_[0]),
		.chany_in_135_(sb_0__1__0_chany_bottom_out_135_[0]),
		.chany_in_136_(sb_0__0__0_chany_top_out_136_[0]),
		.chany_in_137_(sb_0__1__0_chany_bottom_out_137_[0]),
		.chany_in_138_(sb_0__0__0_chany_top_out_138_[0]),
		.chany_in_139_(sb_0__1__0_chany_bottom_out_139_[0]),
		.chany_in_140_(sb_0__0__0_chany_top_out_140_[0]),
		.chany_in_141_(sb_0__1__0_chany_bottom_out_141_[0]),
		.chany_in_142_(sb_0__0__0_chany_top_out_142_[0]),
		.chany_in_143_(sb_0__1__0_chany_bottom_out_143_[0]),
		.chany_in_144_(sb_0__0__0_chany_top_out_144_[0]),
		.chany_in_145_(sb_0__1__0_chany_bottom_out_145_[0]),
		.chany_in_146_(sb_0__0__0_chany_top_out_146_[0]),
		.chany_in_147_(sb_0__1__0_chany_bottom_out_147_[0]),
		.chany_in_148_(sb_0__0__0_chany_top_out_148_[0]),
		.chany_in_149_(sb_0__1__0_chany_bottom_out_149_[0]),
		.chany_in_150_(sb_0__0__0_chany_top_out_150_[0]),
		.chany_in_151_(sb_0__1__0_chany_bottom_out_151_[0]),
		.chany_in_152_(sb_0__0__0_chany_top_out_152_[0]),
		.chany_in_153_(sb_0__1__0_chany_bottom_out_153_[0]),
		.chany_in_154_(sb_0__0__0_chany_top_out_154_[0]),
		.chany_in_155_(sb_0__1__0_chany_bottom_out_155_[0]),
		.chany_in_156_(sb_0__0__0_chany_top_out_156_[0]),
		.chany_in_157_(sb_0__1__0_chany_bottom_out_157_[0]),
		.chany_in_158_(sb_0__0__0_chany_top_out_158_[0]),
		.chany_in_159_(sb_0__1__0_chany_bottom_out_159_[0]),
		.chany_in_160_(sb_0__0__0_chany_top_out_160_[0]),
		.chany_in_161_(sb_0__1__0_chany_bottom_out_161_[0]),
		.chany_in_162_(sb_0__0__0_chany_top_out_162_[0]),
		.chany_in_163_(sb_0__1__0_chany_bottom_out_163_[0]),
		.chany_in_164_(sb_0__0__0_chany_top_out_164_[0]),
		.chany_in_165_(sb_0__1__0_chany_bottom_out_165_[0]),
		.chany_in_166_(sb_0__0__0_chany_top_out_166_[0]),
		.chany_in_167_(sb_0__1__0_chany_bottom_out_167_[0]),
		.chany_in_168_(sb_0__0__0_chany_top_out_168_[0]),
		.chany_in_169_(sb_0__1__0_chany_bottom_out_169_[0]),
		.chany_in_170_(sb_0__0__0_chany_top_out_170_[0]),
		.chany_in_171_(sb_0__1__0_chany_bottom_out_171_[0]),
		.chany_in_172_(sb_0__0__0_chany_top_out_172_[0]),
		.chany_in_173_(sb_0__1__0_chany_bottom_out_173_[0]),
		.chany_in_174_(sb_0__0__0_chany_top_out_174_[0]),
		.chany_in_175_(sb_0__1__0_chany_bottom_out_175_[0]),
		.chany_in_176_(sb_0__0__0_chany_top_out_176_[0]),
		.chany_in_177_(sb_0__1__0_chany_bottom_out_177_[0]),
		.chany_in_178_(sb_0__0__0_chany_top_out_178_[0]),
		.chany_in_179_(sb_0__1__0_chany_bottom_out_179_[0]),
		.chany_in_180_(sb_0__0__0_chany_top_out_180_[0]),
		.chany_in_181_(sb_0__1__0_chany_bottom_out_181_[0]),
		.chany_in_182_(sb_0__0__0_chany_top_out_182_[0]),
		.chany_in_183_(sb_0__1__0_chany_bottom_out_183_[0]),
		.chany_in_184_(sb_0__0__0_chany_top_out_184_[0]),
		.chany_in_185_(sb_0__1__0_chany_bottom_out_185_[0]),
		.chany_in_186_(sb_0__0__0_chany_top_out_186_[0]),
		.chany_in_187_(sb_0__1__0_chany_bottom_out_187_[0]),
		.chany_in_188_(sb_0__0__0_chany_top_out_188_[0]),
		.chany_in_189_(sb_0__1__0_chany_bottom_out_189_[0]),
		.chany_in_190_(sb_0__0__0_chany_top_out_190_[0]),
		.chany_in_191_(sb_0__1__0_chany_bottom_out_191_[0]),
		.chany_in_192_(sb_0__0__0_chany_top_out_192_[0]),
		.chany_in_193_(sb_0__1__0_chany_bottom_out_193_[0]),
		.chany_in_194_(sb_0__0__0_chany_top_out_194_[0]),
		.chany_in_195_(sb_0__1__0_chany_bottom_out_195_[0]),
		.chany_in_196_(sb_0__0__0_chany_top_out_196_[0]),
		.chany_in_197_(sb_0__1__0_chany_bottom_out_197_[0]),
		.chany_in_198_(sb_0__0__0_chany_top_out_198_[0]),
		.chany_in_199_(sb_0__1__0_chany_bottom_out_199_[0]),
		.ccff_head(sb_0__0__0_ccff_tail[0]),
		.chany_out_0_(cby_0__1__0_chany_out_0_[0]),
		.chany_out_1_(cby_0__1__0_chany_out_1_[0]),
		.chany_out_2_(cby_0__1__0_chany_out_2_[0]),
		.chany_out_3_(cby_0__1__0_chany_out_3_[0]),
		.chany_out_4_(cby_0__1__0_chany_out_4_[0]),
		.chany_out_5_(cby_0__1__0_chany_out_5_[0]),
		.chany_out_6_(cby_0__1__0_chany_out_6_[0]),
		.chany_out_7_(cby_0__1__0_chany_out_7_[0]),
		.chany_out_8_(cby_0__1__0_chany_out_8_[0]),
		.chany_out_9_(cby_0__1__0_chany_out_9_[0]),
		.chany_out_10_(cby_0__1__0_chany_out_10_[0]),
		.chany_out_11_(cby_0__1__0_chany_out_11_[0]),
		.chany_out_12_(cby_0__1__0_chany_out_12_[0]),
		.chany_out_13_(cby_0__1__0_chany_out_13_[0]),
		.chany_out_14_(cby_0__1__0_chany_out_14_[0]),
		.chany_out_15_(cby_0__1__0_chany_out_15_[0]),
		.chany_out_16_(cby_0__1__0_chany_out_16_[0]),
		.chany_out_17_(cby_0__1__0_chany_out_17_[0]),
		.chany_out_18_(cby_0__1__0_chany_out_18_[0]),
		.chany_out_19_(cby_0__1__0_chany_out_19_[0]),
		.chany_out_20_(cby_0__1__0_chany_out_20_[0]),
		.chany_out_21_(cby_0__1__0_chany_out_21_[0]),
		.chany_out_22_(cby_0__1__0_chany_out_22_[0]),
		.chany_out_23_(cby_0__1__0_chany_out_23_[0]),
		.chany_out_24_(cby_0__1__0_chany_out_24_[0]),
		.chany_out_25_(cby_0__1__0_chany_out_25_[0]),
		.chany_out_26_(cby_0__1__0_chany_out_26_[0]),
		.chany_out_27_(cby_0__1__0_chany_out_27_[0]),
		.chany_out_28_(cby_0__1__0_chany_out_28_[0]),
		.chany_out_29_(cby_0__1__0_chany_out_29_[0]),
		.chany_out_30_(cby_0__1__0_chany_out_30_[0]),
		.chany_out_31_(cby_0__1__0_chany_out_31_[0]),
		.chany_out_32_(cby_0__1__0_chany_out_32_[0]),
		.chany_out_33_(cby_0__1__0_chany_out_33_[0]),
		.chany_out_34_(cby_0__1__0_chany_out_34_[0]),
		.chany_out_35_(cby_0__1__0_chany_out_35_[0]),
		.chany_out_36_(cby_0__1__0_chany_out_36_[0]),
		.chany_out_37_(cby_0__1__0_chany_out_37_[0]),
		.chany_out_38_(cby_0__1__0_chany_out_38_[0]),
		.chany_out_39_(cby_0__1__0_chany_out_39_[0]),
		.chany_out_40_(cby_0__1__0_chany_out_40_[0]),
		.chany_out_41_(cby_0__1__0_chany_out_41_[0]),
		.chany_out_42_(cby_0__1__0_chany_out_42_[0]),
		.chany_out_43_(cby_0__1__0_chany_out_43_[0]),
		.chany_out_44_(cby_0__1__0_chany_out_44_[0]),
		.chany_out_45_(cby_0__1__0_chany_out_45_[0]),
		.chany_out_46_(cby_0__1__0_chany_out_46_[0]),
		.chany_out_47_(cby_0__1__0_chany_out_47_[0]),
		.chany_out_48_(cby_0__1__0_chany_out_48_[0]),
		.chany_out_49_(cby_0__1__0_chany_out_49_[0]),
		.chany_out_50_(cby_0__1__0_chany_out_50_[0]),
		.chany_out_51_(cby_0__1__0_chany_out_51_[0]),
		.chany_out_52_(cby_0__1__0_chany_out_52_[0]),
		.chany_out_53_(cby_0__1__0_chany_out_53_[0]),
		.chany_out_54_(cby_0__1__0_chany_out_54_[0]),
		.chany_out_55_(cby_0__1__0_chany_out_55_[0]),
		.chany_out_56_(cby_0__1__0_chany_out_56_[0]),
		.chany_out_57_(cby_0__1__0_chany_out_57_[0]),
		.chany_out_58_(cby_0__1__0_chany_out_58_[0]),
		.chany_out_59_(cby_0__1__0_chany_out_59_[0]),
		.chany_out_60_(cby_0__1__0_chany_out_60_[0]),
		.chany_out_61_(cby_0__1__0_chany_out_61_[0]),
		.chany_out_62_(cby_0__1__0_chany_out_62_[0]),
		.chany_out_63_(cby_0__1__0_chany_out_63_[0]),
		.chany_out_64_(cby_0__1__0_chany_out_64_[0]),
		.chany_out_65_(cby_0__1__0_chany_out_65_[0]),
		.chany_out_66_(cby_0__1__0_chany_out_66_[0]),
		.chany_out_67_(cby_0__1__0_chany_out_67_[0]),
		.chany_out_68_(cby_0__1__0_chany_out_68_[0]),
		.chany_out_69_(cby_0__1__0_chany_out_69_[0]),
		.chany_out_70_(cby_0__1__0_chany_out_70_[0]),
		.chany_out_71_(cby_0__1__0_chany_out_71_[0]),
		.chany_out_72_(cby_0__1__0_chany_out_72_[0]),
		.chany_out_73_(cby_0__1__0_chany_out_73_[0]),
		.chany_out_74_(cby_0__1__0_chany_out_74_[0]),
		.chany_out_75_(cby_0__1__0_chany_out_75_[0]),
		.chany_out_76_(cby_0__1__0_chany_out_76_[0]),
		.chany_out_77_(cby_0__1__0_chany_out_77_[0]),
		.chany_out_78_(cby_0__1__0_chany_out_78_[0]),
		.chany_out_79_(cby_0__1__0_chany_out_79_[0]),
		.chany_out_80_(cby_0__1__0_chany_out_80_[0]),
		.chany_out_81_(cby_0__1__0_chany_out_81_[0]),
		.chany_out_82_(cby_0__1__0_chany_out_82_[0]),
		.chany_out_83_(cby_0__1__0_chany_out_83_[0]),
		.chany_out_84_(cby_0__1__0_chany_out_84_[0]),
		.chany_out_85_(cby_0__1__0_chany_out_85_[0]),
		.chany_out_86_(cby_0__1__0_chany_out_86_[0]),
		.chany_out_87_(cby_0__1__0_chany_out_87_[0]),
		.chany_out_88_(cby_0__1__0_chany_out_88_[0]),
		.chany_out_89_(cby_0__1__0_chany_out_89_[0]),
		.chany_out_90_(cby_0__1__0_chany_out_90_[0]),
		.chany_out_91_(cby_0__1__0_chany_out_91_[0]),
		.chany_out_92_(cby_0__1__0_chany_out_92_[0]),
		.chany_out_93_(cby_0__1__0_chany_out_93_[0]),
		.chany_out_94_(cby_0__1__0_chany_out_94_[0]),
		.chany_out_95_(cby_0__1__0_chany_out_95_[0]),
		.chany_out_96_(cby_0__1__0_chany_out_96_[0]),
		.chany_out_97_(cby_0__1__0_chany_out_97_[0]),
		.chany_out_98_(cby_0__1__0_chany_out_98_[0]),
		.chany_out_99_(cby_0__1__0_chany_out_99_[0]),
		.chany_out_100_(cby_0__1__0_chany_out_100_[0]),
		.chany_out_101_(cby_0__1__0_chany_out_101_[0]),
		.chany_out_102_(cby_0__1__0_chany_out_102_[0]),
		.chany_out_103_(cby_0__1__0_chany_out_103_[0]),
		.chany_out_104_(cby_0__1__0_chany_out_104_[0]),
		.chany_out_105_(cby_0__1__0_chany_out_105_[0]),
		.chany_out_106_(cby_0__1__0_chany_out_106_[0]),
		.chany_out_107_(cby_0__1__0_chany_out_107_[0]),
		.chany_out_108_(cby_0__1__0_chany_out_108_[0]),
		.chany_out_109_(cby_0__1__0_chany_out_109_[0]),
		.chany_out_110_(cby_0__1__0_chany_out_110_[0]),
		.chany_out_111_(cby_0__1__0_chany_out_111_[0]),
		.chany_out_112_(cby_0__1__0_chany_out_112_[0]),
		.chany_out_113_(cby_0__1__0_chany_out_113_[0]),
		.chany_out_114_(cby_0__1__0_chany_out_114_[0]),
		.chany_out_115_(cby_0__1__0_chany_out_115_[0]),
		.chany_out_116_(cby_0__1__0_chany_out_116_[0]),
		.chany_out_117_(cby_0__1__0_chany_out_117_[0]),
		.chany_out_118_(cby_0__1__0_chany_out_118_[0]),
		.chany_out_119_(cby_0__1__0_chany_out_119_[0]),
		.chany_out_120_(cby_0__1__0_chany_out_120_[0]),
		.chany_out_121_(cby_0__1__0_chany_out_121_[0]),
		.chany_out_122_(cby_0__1__0_chany_out_122_[0]),
		.chany_out_123_(cby_0__1__0_chany_out_123_[0]),
		.chany_out_124_(cby_0__1__0_chany_out_124_[0]),
		.chany_out_125_(cby_0__1__0_chany_out_125_[0]),
		.chany_out_126_(cby_0__1__0_chany_out_126_[0]),
		.chany_out_127_(cby_0__1__0_chany_out_127_[0]),
		.chany_out_128_(cby_0__1__0_chany_out_128_[0]),
		.chany_out_129_(cby_0__1__0_chany_out_129_[0]),
		.chany_out_130_(cby_0__1__0_chany_out_130_[0]),
		.chany_out_131_(cby_0__1__0_chany_out_131_[0]),
		.chany_out_132_(cby_0__1__0_chany_out_132_[0]),
		.chany_out_133_(cby_0__1__0_chany_out_133_[0]),
		.chany_out_134_(cby_0__1__0_chany_out_134_[0]),
		.chany_out_135_(cby_0__1__0_chany_out_135_[0]),
		.chany_out_136_(cby_0__1__0_chany_out_136_[0]),
		.chany_out_137_(cby_0__1__0_chany_out_137_[0]),
		.chany_out_138_(cby_0__1__0_chany_out_138_[0]),
		.chany_out_139_(cby_0__1__0_chany_out_139_[0]),
		.chany_out_140_(cby_0__1__0_chany_out_140_[0]),
		.chany_out_141_(cby_0__1__0_chany_out_141_[0]),
		.chany_out_142_(cby_0__1__0_chany_out_142_[0]),
		.chany_out_143_(cby_0__1__0_chany_out_143_[0]),
		.chany_out_144_(cby_0__1__0_chany_out_144_[0]),
		.chany_out_145_(cby_0__1__0_chany_out_145_[0]),
		.chany_out_146_(cby_0__1__0_chany_out_146_[0]),
		.chany_out_147_(cby_0__1__0_chany_out_147_[0]),
		.chany_out_148_(cby_0__1__0_chany_out_148_[0]),
		.chany_out_149_(cby_0__1__0_chany_out_149_[0]),
		.chany_out_150_(cby_0__1__0_chany_out_150_[0]),
		.chany_out_151_(cby_0__1__0_chany_out_151_[0]),
		.chany_out_152_(cby_0__1__0_chany_out_152_[0]),
		.chany_out_153_(cby_0__1__0_chany_out_153_[0]),
		.chany_out_154_(cby_0__1__0_chany_out_154_[0]),
		.chany_out_155_(cby_0__1__0_chany_out_155_[0]),
		.chany_out_156_(cby_0__1__0_chany_out_156_[0]),
		.chany_out_157_(cby_0__1__0_chany_out_157_[0]),
		.chany_out_158_(cby_0__1__0_chany_out_158_[0]),
		.chany_out_159_(cby_0__1__0_chany_out_159_[0]),
		.chany_out_160_(cby_0__1__0_chany_out_160_[0]),
		.chany_out_161_(cby_0__1__0_chany_out_161_[0]),
		.chany_out_162_(cby_0__1__0_chany_out_162_[0]),
		.chany_out_163_(cby_0__1__0_chany_out_163_[0]),
		.chany_out_164_(cby_0__1__0_chany_out_164_[0]),
		.chany_out_165_(cby_0__1__0_chany_out_165_[0]),
		.chany_out_166_(cby_0__1__0_chany_out_166_[0]),
		.chany_out_167_(cby_0__1__0_chany_out_167_[0]),
		.chany_out_168_(cby_0__1__0_chany_out_168_[0]),
		.chany_out_169_(cby_0__1__0_chany_out_169_[0]),
		.chany_out_170_(cby_0__1__0_chany_out_170_[0]),
		.chany_out_171_(cby_0__1__0_chany_out_171_[0]),
		.chany_out_172_(cby_0__1__0_chany_out_172_[0]),
		.chany_out_173_(cby_0__1__0_chany_out_173_[0]),
		.chany_out_174_(cby_0__1__0_chany_out_174_[0]),
		.chany_out_175_(cby_0__1__0_chany_out_175_[0]),
		.chany_out_176_(cby_0__1__0_chany_out_176_[0]),
		.chany_out_177_(cby_0__1__0_chany_out_177_[0]),
		.chany_out_178_(cby_0__1__0_chany_out_178_[0]),
		.chany_out_179_(cby_0__1__0_chany_out_179_[0]),
		.chany_out_180_(cby_0__1__0_chany_out_180_[0]),
		.chany_out_181_(cby_0__1__0_chany_out_181_[0]),
		.chany_out_182_(cby_0__1__0_chany_out_182_[0]),
		.chany_out_183_(cby_0__1__0_chany_out_183_[0]),
		.chany_out_184_(cby_0__1__0_chany_out_184_[0]),
		.chany_out_185_(cby_0__1__0_chany_out_185_[0]),
		.chany_out_186_(cby_0__1__0_chany_out_186_[0]),
		.chany_out_187_(cby_0__1__0_chany_out_187_[0]),
		.chany_out_188_(cby_0__1__0_chany_out_188_[0]),
		.chany_out_189_(cby_0__1__0_chany_out_189_[0]),
		.chany_out_190_(cby_0__1__0_chany_out_190_[0]),
		.chany_out_191_(cby_0__1__0_chany_out_191_[0]),
		.chany_out_192_(cby_0__1__0_chany_out_192_[0]),
		.chany_out_193_(cby_0__1__0_chany_out_193_[0]),
		.chany_out_194_(cby_0__1__0_chany_out_194_[0]),
		.chany_out_195_(cby_0__1__0_chany_out_195_[0]),
		.chany_out_196_(cby_0__1__0_chany_out_196_[0]),
		.chany_out_197_(cby_0__1__0_chany_out_197_[0]),
		.chany_out_198_(cby_0__1__0_chany_out_198_[0]),
		.chany_out_199_(cby_0__1__0_chany_out_199_[0]),
		.left_grid_pin_0_(cby_0__1__0_left_grid_pin_0_[0]),
		.ccff_tail(cby_0__1__0_ccff_tail[0]));

	cby_0__1_ cby_0__2_ (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.chany_in_0_(sb_0__1__0_chany_top_out_0_[0]),
		.chany_in_1_(sb_0__2__0_chany_bottom_out_1_[0]),
		.chany_in_2_(sb_0__1__0_chany_top_out_2_[0]),
		.chany_in_3_(sb_0__2__0_chany_bottom_out_3_[0]),
		.chany_in_4_(sb_0__1__0_chany_top_out_4_[0]),
		.chany_in_5_(sb_0__2__0_chany_bottom_out_5_[0]),
		.chany_in_6_(sb_0__1__0_chany_top_out_6_[0]),
		.chany_in_7_(sb_0__2__0_chany_bottom_out_7_[0]),
		.chany_in_8_(sb_0__1__0_chany_top_out_8_[0]),
		.chany_in_9_(sb_0__2__0_chany_bottom_out_9_[0]),
		.chany_in_10_(sb_0__1__0_chany_top_out_10_[0]),
		.chany_in_11_(sb_0__2__0_chany_bottom_out_11_[0]),
		.chany_in_12_(sb_0__1__0_chany_top_out_12_[0]),
		.chany_in_13_(sb_0__2__0_chany_bottom_out_13_[0]),
		.chany_in_14_(sb_0__1__0_chany_top_out_14_[0]),
		.chany_in_15_(sb_0__2__0_chany_bottom_out_15_[0]),
		.chany_in_16_(sb_0__1__0_chany_top_out_16_[0]),
		.chany_in_17_(sb_0__2__0_chany_bottom_out_17_[0]),
		.chany_in_18_(sb_0__1__0_chany_top_out_18_[0]),
		.chany_in_19_(sb_0__2__0_chany_bottom_out_19_[0]),
		.chany_in_20_(sb_0__1__0_chany_top_out_20_[0]),
		.chany_in_21_(sb_0__2__0_chany_bottom_out_21_[0]),
		.chany_in_22_(sb_0__1__0_chany_top_out_22_[0]),
		.chany_in_23_(sb_0__2__0_chany_bottom_out_23_[0]),
		.chany_in_24_(sb_0__1__0_chany_top_out_24_[0]),
		.chany_in_25_(sb_0__2__0_chany_bottom_out_25_[0]),
		.chany_in_26_(sb_0__1__0_chany_top_out_26_[0]),
		.chany_in_27_(sb_0__2__0_chany_bottom_out_27_[0]),
		.chany_in_28_(sb_0__1__0_chany_top_out_28_[0]),
		.chany_in_29_(sb_0__2__0_chany_bottom_out_29_[0]),
		.chany_in_30_(sb_0__1__0_chany_top_out_30_[0]),
		.chany_in_31_(sb_0__2__0_chany_bottom_out_31_[0]),
		.chany_in_32_(sb_0__1__0_chany_top_out_32_[0]),
		.chany_in_33_(sb_0__2__0_chany_bottom_out_33_[0]),
		.chany_in_34_(sb_0__1__0_chany_top_out_34_[0]),
		.chany_in_35_(sb_0__2__0_chany_bottom_out_35_[0]),
		.chany_in_36_(sb_0__1__0_chany_top_out_36_[0]),
		.chany_in_37_(sb_0__2__0_chany_bottom_out_37_[0]),
		.chany_in_38_(sb_0__1__0_chany_top_out_38_[0]),
		.chany_in_39_(sb_0__2__0_chany_bottom_out_39_[0]),
		.chany_in_40_(sb_0__1__0_chany_top_out_40_[0]),
		.chany_in_41_(sb_0__2__0_chany_bottom_out_41_[0]),
		.chany_in_42_(sb_0__1__0_chany_top_out_42_[0]),
		.chany_in_43_(sb_0__2__0_chany_bottom_out_43_[0]),
		.chany_in_44_(sb_0__1__0_chany_top_out_44_[0]),
		.chany_in_45_(sb_0__2__0_chany_bottom_out_45_[0]),
		.chany_in_46_(sb_0__1__0_chany_top_out_46_[0]),
		.chany_in_47_(sb_0__2__0_chany_bottom_out_47_[0]),
		.chany_in_48_(sb_0__1__0_chany_top_out_48_[0]),
		.chany_in_49_(sb_0__2__0_chany_bottom_out_49_[0]),
		.chany_in_50_(sb_0__1__0_chany_top_out_50_[0]),
		.chany_in_51_(sb_0__2__0_chany_bottom_out_51_[0]),
		.chany_in_52_(sb_0__1__0_chany_top_out_52_[0]),
		.chany_in_53_(sb_0__2__0_chany_bottom_out_53_[0]),
		.chany_in_54_(sb_0__1__0_chany_top_out_54_[0]),
		.chany_in_55_(sb_0__2__0_chany_bottom_out_55_[0]),
		.chany_in_56_(sb_0__1__0_chany_top_out_56_[0]),
		.chany_in_57_(sb_0__2__0_chany_bottom_out_57_[0]),
		.chany_in_58_(sb_0__1__0_chany_top_out_58_[0]),
		.chany_in_59_(sb_0__2__0_chany_bottom_out_59_[0]),
		.chany_in_60_(sb_0__1__0_chany_top_out_60_[0]),
		.chany_in_61_(sb_0__2__0_chany_bottom_out_61_[0]),
		.chany_in_62_(sb_0__1__0_chany_top_out_62_[0]),
		.chany_in_63_(sb_0__2__0_chany_bottom_out_63_[0]),
		.chany_in_64_(sb_0__1__0_chany_top_out_64_[0]),
		.chany_in_65_(sb_0__2__0_chany_bottom_out_65_[0]),
		.chany_in_66_(sb_0__1__0_chany_top_out_66_[0]),
		.chany_in_67_(sb_0__2__0_chany_bottom_out_67_[0]),
		.chany_in_68_(sb_0__1__0_chany_top_out_68_[0]),
		.chany_in_69_(sb_0__2__0_chany_bottom_out_69_[0]),
		.chany_in_70_(sb_0__1__0_chany_top_out_70_[0]),
		.chany_in_71_(sb_0__2__0_chany_bottom_out_71_[0]),
		.chany_in_72_(sb_0__1__0_chany_top_out_72_[0]),
		.chany_in_73_(sb_0__2__0_chany_bottom_out_73_[0]),
		.chany_in_74_(sb_0__1__0_chany_top_out_74_[0]),
		.chany_in_75_(sb_0__2__0_chany_bottom_out_75_[0]),
		.chany_in_76_(sb_0__1__0_chany_top_out_76_[0]),
		.chany_in_77_(sb_0__2__0_chany_bottom_out_77_[0]),
		.chany_in_78_(sb_0__1__0_chany_top_out_78_[0]),
		.chany_in_79_(sb_0__2__0_chany_bottom_out_79_[0]),
		.chany_in_80_(sb_0__1__0_chany_top_out_80_[0]),
		.chany_in_81_(sb_0__2__0_chany_bottom_out_81_[0]),
		.chany_in_82_(sb_0__1__0_chany_top_out_82_[0]),
		.chany_in_83_(sb_0__2__0_chany_bottom_out_83_[0]),
		.chany_in_84_(sb_0__1__0_chany_top_out_84_[0]),
		.chany_in_85_(sb_0__2__0_chany_bottom_out_85_[0]),
		.chany_in_86_(sb_0__1__0_chany_top_out_86_[0]),
		.chany_in_87_(sb_0__2__0_chany_bottom_out_87_[0]),
		.chany_in_88_(sb_0__1__0_chany_top_out_88_[0]),
		.chany_in_89_(sb_0__2__0_chany_bottom_out_89_[0]),
		.chany_in_90_(sb_0__1__0_chany_top_out_90_[0]),
		.chany_in_91_(sb_0__2__0_chany_bottom_out_91_[0]),
		.chany_in_92_(sb_0__1__0_chany_top_out_92_[0]),
		.chany_in_93_(sb_0__2__0_chany_bottom_out_93_[0]),
		.chany_in_94_(sb_0__1__0_chany_top_out_94_[0]),
		.chany_in_95_(sb_0__2__0_chany_bottom_out_95_[0]),
		.chany_in_96_(sb_0__1__0_chany_top_out_96_[0]),
		.chany_in_97_(sb_0__2__0_chany_bottom_out_97_[0]),
		.chany_in_98_(sb_0__1__0_chany_top_out_98_[0]),
		.chany_in_99_(sb_0__2__0_chany_bottom_out_99_[0]),
		.chany_in_100_(sb_0__1__0_chany_top_out_100_[0]),
		.chany_in_101_(sb_0__2__0_chany_bottom_out_101_[0]),
		.chany_in_102_(sb_0__1__0_chany_top_out_102_[0]),
		.chany_in_103_(sb_0__2__0_chany_bottom_out_103_[0]),
		.chany_in_104_(sb_0__1__0_chany_top_out_104_[0]),
		.chany_in_105_(sb_0__2__0_chany_bottom_out_105_[0]),
		.chany_in_106_(sb_0__1__0_chany_top_out_106_[0]),
		.chany_in_107_(sb_0__2__0_chany_bottom_out_107_[0]),
		.chany_in_108_(sb_0__1__0_chany_top_out_108_[0]),
		.chany_in_109_(sb_0__2__0_chany_bottom_out_109_[0]),
		.chany_in_110_(sb_0__1__0_chany_top_out_110_[0]),
		.chany_in_111_(sb_0__2__0_chany_bottom_out_111_[0]),
		.chany_in_112_(sb_0__1__0_chany_top_out_112_[0]),
		.chany_in_113_(sb_0__2__0_chany_bottom_out_113_[0]),
		.chany_in_114_(sb_0__1__0_chany_top_out_114_[0]),
		.chany_in_115_(sb_0__2__0_chany_bottom_out_115_[0]),
		.chany_in_116_(sb_0__1__0_chany_top_out_116_[0]),
		.chany_in_117_(sb_0__2__0_chany_bottom_out_117_[0]),
		.chany_in_118_(sb_0__1__0_chany_top_out_118_[0]),
		.chany_in_119_(sb_0__2__0_chany_bottom_out_119_[0]),
		.chany_in_120_(sb_0__1__0_chany_top_out_120_[0]),
		.chany_in_121_(sb_0__2__0_chany_bottom_out_121_[0]),
		.chany_in_122_(sb_0__1__0_chany_top_out_122_[0]),
		.chany_in_123_(sb_0__2__0_chany_bottom_out_123_[0]),
		.chany_in_124_(sb_0__1__0_chany_top_out_124_[0]),
		.chany_in_125_(sb_0__2__0_chany_bottom_out_125_[0]),
		.chany_in_126_(sb_0__1__0_chany_top_out_126_[0]),
		.chany_in_127_(sb_0__2__0_chany_bottom_out_127_[0]),
		.chany_in_128_(sb_0__1__0_chany_top_out_128_[0]),
		.chany_in_129_(sb_0__2__0_chany_bottom_out_129_[0]),
		.chany_in_130_(sb_0__1__0_chany_top_out_130_[0]),
		.chany_in_131_(sb_0__2__0_chany_bottom_out_131_[0]),
		.chany_in_132_(sb_0__1__0_chany_top_out_132_[0]),
		.chany_in_133_(sb_0__2__0_chany_bottom_out_133_[0]),
		.chany_in_134_(sb_0__1__0_chany_top_out_134_[0]),
		.chany_in_135_(sb_0__2__0_chany_bottom_out_135_[0]),
		.chany_in_136_(sb_0__1__0_chany_top_out_136_[0]),
		.chany_in_137_(sb_0__2__0_chany_bottom_out_137_[0]),
		.chany_in_138_(sb_0__1__0_chany_top_out_138_[0]),
		.chany_in_139_(sb_0__2__0_chany_bottom_out_139_[0]),
		.chany_in_140_(sb_0__1__0_chany_top_out_140_[0]),
		.chany_in_141_(sb_0__2__0_chany_bottom_out_141_[0]),
		.chany_in_142_(sb_0__1__0_chany_top_out_142_[0]),
		.chany_in_143_(sb_0__2__0_chany_bottom_out_143_[0]),
		.chany_in_144_(sb_0__1__0_chany_top_out_144_[0]),
		.chany_in_145_(sb_0__2__0_chany_bottom_out_145_[0]),
		.chany_in_146_(sb_0__1__0_chany_top_out_146_[0]),
		.chany_in_147_(sb_0__2__0_chany_bottom_out_147_[0]),
		.chany_in_148_(sb_0__1__0_chany_top_out_148_[0]),
		.chany_in_149_(sb_0__2__0_chany_bottom_out_149_[0]),
		.chany_in_150_(sb_0__1__0_chany_top_out_150_[0]),
		.chany_in_151_(sb_0__2__0_chany_bottom_out_151_[0]),
		.chany_in_152_(sb_0__1__0_chany_top_out_152_[0]),
		.chany_in_153_(sb_0__2__0_chany_bottom_out_153_[0]),
		.chany_in_154_(sb_0__1__0_chany_top_out_154_[0]),
		.chany_in_155_(sb_0__2__0_chany_bottom_out_155_[0]),
		.chany_in_156_(sb_0__1__0_chany_top_out_156_[0]),
		.chany_in_157_(sb_0__2__0_chany_bottom_out_157_[0]),
		.chany_in_158_(sb_0__1__0_chany_top_out_158_[0]),
		.chany_in_159_(sb_0__2__0_chany_bottom_out_159_[0]),
		.chany_in_160_(sb_0__1__0_chany_top_out_160_[0]),
		.chany_in_161_(sb_0__2__0_chany_bottom_out_161_[0]),
		.chany_in_162_(sb_0__1__0_chany_top_out_162_[0]),
		.chany_in_163_(sb_0__2__0_chany_bottom_out_163_[0]),
		.chany_in_164_(sb_0__1__0_chany_top_out_164_[0]),
		.chany_in_165_(sb_0__2__0_chany_bottom_out_165_[0]),
		.chany_in_166_(sb_0__1__0_chany_top_out_166_[0]),
		.chany_in_167_(sb_0__2__0_chany_bottom_out_167_[0]),
		.chany_in_168_(sb_0__1__0_chany_top_out_168_[0]),
		.chany_in_169_(sb_0__2__0_chany_bottom_out_169_[0]),
		.chany_in_170_(sb_0__1__0_chany_top_out_170_[0]),
		.chany_in_171_(sb_0__2__0_chany_bottom_out_171_[0]),
		.chany_in_172_(sb_0__1__0_chany_top_out_172_[0]),
		.chany_in_173_(sb_0__2__0_chany_bottom_out_173_[0]),
		.chany_in_174_(sb_0__1__0_chany_top_out_174_[0]),
		.chany_in_175_(sb_0__2__0_chany_bottom_out_175_[0]),
		.chany_in_176_(sb_0__1__0_chany_top_out_176_[0]),
		.chany_in_177_(sb_0__2__0_chany_bottom_out_177_[0]),
		.chany_in_178_(sb_0__1__0_chany_top_out_178_[0]),
		.chany_in_179_(sb_0__2__0_chany_bottom_out_179_[0]),
		.chany_in_180_(sb_0__1__0_chany_top_out_180_[0]),
		.chany_in_181_(sb_0__2__0_chany_bottom_out_181_[0]),
		.chany_in_182_(sb_0__1__0_chany_top_out_182_[0]),
		.chany_in_183_(sb_0__2__0_chany_bottom_out_183_[0]),
		.chany_in_184_(sb_0__1__0_chany_top_out_184_[0]),
		.chany_in_185_(sb_0__2__0_chany_bottom_out_185_[0]),
		.chany_in_186_(sb_0__1__0_chany_top_out_186_[0]),
		.chany_in_187_(sb_0__2__0_chany_bottom_out_187_[0]),
		.chany_in_188_(sb_0__1__0_chany_top_out_188_[0]),
		.chany_in_189_(sb_0__2__0_chany_bottom_out_189_[0]),
		.chany_in_190_(sb_0__1__0_chany_top_out_190_[0]),
		.chany_in_191_(sb_0__2__0_chany_bottom_out_191_[0]),
		.chany_in_192_(sb_0__1__0_chany_top_out_192_[0]),
		.chany_in_193_(sb_0__2__0_chany_bottom_out_193_[0]),
		.chany_in_194_(sb_0__1__0_chany_top_out_194_[0]),
		.chany_in_195_(sb_0__2__0_chany_bottom_out_195_[0]),
		.chany_in_196_(sb_0__1__0_chany_top_out_196_[0]),
		.chany_in_197_(sb_0__2__0_chany_bottom_out_197_[0]),
		.chany_in_198_(sb_0__1__0_chany_top_out_198_[0]),
		.chany_in_199_(sb_0__2__0_chany_bottom_out_199_[0]),
		.ccff_head(sb_0__1__0_ccff_tail[0]),
		.chany_out_0_(cby_0__1__1_chany_out_0_[0]),
		.chany_out_1_(cby_0__1__1_chany_out_1_[0]),
		.chany_out_2_(cby_0__1__1_chany_out_2_[0]),
		.chany_out_3_(cby_0__1__1_chany_out_3_[0]),
		.chany_out_4_(cby_0__1__1_chany_out_4_[0]),
		.chany_out_5_(cby_0__1__1_chany_out_5_[0]),
		.chany_out_6_(cby_0__1__1_chany_out_6_[0]),
		.chany_out_7_(cby_0__1__1_chany_out_7_[0]),
		.chany_out_8_(cby_0__1__1_chany_out_8_[0]),
		.chany_out_9_(cby_0__1__1_chany_out_9_[0]),
		.chany_out_10_(cby_0__1__1_chany_out_10_[0]),
		.chany_out_11_(cby_0__1__1_chany_out_11_[0]),
		.chany_out_12_(cby_0__1__1_chany_out_12_[0]),
		.chany_out_13_(cby_0__1__1_chany_out_13_[0]),
		.chany_out_14_(cby_0__1__1_chany_out_14_[0]),
		.chany_out_15_(cby_0__1__1_chany_out_15_[0]),
		.chany_out_16_(cby_0__1__1_chany_out_16_[0]),
		.chany_out_17_(cby_0__1__1_chany_out_17_[0]),
		.chany_out_18_(cby_0__1__1_chany_out_18_[0]),
		.chany_out_19_(cby_0__1__1_chany_out_19_[0]),
		.chany_out_20_(cby_0__1__1_chany_out_20_[0]),
		.chany_out_21_(cby_0__1__1_chany_out_21_[0]),
		.chany_out_22_(cby_0__1__1_chany_out_22_[0]),
		.chany_out_23_(cby_0__1__1_chany_out_23_[0]),
		.chany_out_24_(cby_0__1__1_chany_out_24_[0]),
		.chany_out_25_(cby_0__1__1_chany_out_25_[0]),
		.chany_out_26_(cby_0__1__1_chany_out_26_[0]),
		.chany_out_27_(cby_0__1__1_chany_out_27_[0]),
		.chany_out_28_(cby_0__1__1_chany_out_28_[0]),
		.chany_out_29_(cby_0__1__1_chany_out_29_[0]),
		.chany_out_30_(cby_0__1__1_chany_out_30_[0]),
		.chany_out_31_(cby_0__1__1_chany_out_31_[0]),
		.chany_out_32_(cby_0__1__1_chany_out_32_[0]),
		.chany_out_33_(cby_0__1__1_chany_out_33_[0]),
		.chany_out_34_(cby_0__1__1_chany_out_34_[0]),
		.chany_out_35_(cby_0__1__1_chany_out_35_[0]),
		.chany_out_36_(cby_0__1__1_chany_out_36_[0]),
		.chany_out_37_(cby_0__1__1_chany_out_37_[0]),
		.chany_out_38_(cby_0__1__1_chany_out_38_[0]),
		.chany_out_39_(cby_0__1__1_chany_out_39_[0]),
		.chany_out_40_(cby_0__1__1_chany_out_40_[0]),
		.chany_out_41_(cby_0__1__1_chany_out_41_[0]),
		.chany_out_42_(cby_0__1__1_chany_out_42_[0]),
		.chany_out_43_(cby_0__1__1_chany_out_43_[0]),
		.chany_out_44_(cby_0__1__1_chany_out_44_[0]),
		.chany_out_45_(cby_0__1__1_chany_out_45_[0]),
		.chany_out_46_(cby_0__1__1_chany_out_46_[0]),
		.chany_out_47_(cby_0__1__1_chany_out_47_[0]),
		.chany_out_48_(cby_0__1__1_chany_out_48_[0]),
		.chany_out_49_(cby_0__1__1_chany_out_49_[0]),
		.chany_out_50_(cby_0__1__1_chany_out_50_[0]),
		.chany_out_51_(cby_0__1__1_chany_out_51_[0]),
		.chany_out_52_(cby_0__1__1_chany_out_52_[0]),
		.chany_out_53_(cby_0__1__1_chany_out_53_[0]),
		.chany_out_54_(cby_0__1__1_chany_out_54_[0]),
		.chany_out_55_(cby_0__1__1_chany_out_55_[0]),
		.chany_out_56_(cby_0__1__1_chany_out_56_[0]),
		.chany_out_57_(cby_0__1__1_chany_out_57_[0]),
		.chany_out_58_(cby_0__1__1_chany_out_58_[0]),
		.chany_out_59_(cby_0__1__1_chany_out_59_[0]),
		.chany_out_60_(cby_0__1__1_chany_out_60_[0]),
		.chany_out_61_(cby_0__1__1_chany_out_61_[0]),
		.chany_out_62_(cby_0__1__1_chany_out_62_[0]),
		.chany_out_63_(cby_0__1__1_chany_out_63_[0]),
		.chany_out_64_(cby_0__1__1_chany_out_64_[0]),
		.chany_out_65_(cby_0__1__1_chany_out_65_[0]),
		.chany_out_66_(cby_0__1__1_chany_out_66_[0]),
		.chany_out_67_(cby_0__1__1_chany_out_67_[0]),
		.chany_out_68_(cby_0__1__1_chany_out_68_[0]),
		.chany_out_69_(cby_0__1__1_chany_out_69_[0]),
		.chany_out_70_(cby_0__1__1_chany_out_70_[0]),
		.chany_out_71_(cby_0__1__1_chany_out_71_[0]),
		.chany_out_72_(cby_0__1__1_chany_out_72_[0]),
		.chany_out_73_(cby_0__1__1_chany_out_73_[0]),
		.chany_out_74_(cby_0__1__1_chany_out_74_[0]),
		.chany_out_75_(cby_0__1__1_chany_out_75_[0]),
		.chany_out_76_(cby_0__1__1_chany_out_76_[0]),
		.chany_out_77_(cby_0__1__1_chany_out_77_[0]),
		.chany_out_78_(cby_0__1__1_chany_out_78_[0]),
		.chany_out_79_(cby_0__1__1_chany_out_79_[0]),
		.chany_out_80_(cby_0__1__1_chany_out_80_[0]),
		.chany_out_81_(cby_0__1__1_chany_out_81_[0]),
		.chany_out_82_(cby_0__1__1_chany_out_82_[0]),
		.chany_out_83_(cby_0__1__1_chany_out_83_[0]),
		.chany_out_84_(cby_0__1__1_chany_out_84_[0]),
		.chany_out_85_(cby_0__1__1_chany_out_85_[0]),
		.chany_out_86_(cby_0__1__1_chany_out_86_[0]),
		.chany_out_87_(cby_0__1__1_chany_out_87_[0]),
		.chany_out_88_(cby_0__1__1_chany_out_88_[0]),
		.chany_out_89_(cby_0__1__1_chany_out_89_[0]),
		.chany_out_90_(cby_0__1__1_chany_out_90_[0]),
		.chany_out_91_(cby_0__1__1_chany_out_91_[0]),
		.chany_out_92_(cby_0__1__1_chany_out_92_[0]),
		.chany_out_93_(cby_0__1__1_chany_out_93_[0]),
		.chany_out_94_(cby_0__1__1_chany_out_94_[0]),
		.chany_out_95_(cby_0__1__1_chany_out_95_[0]),
		.chany_out_96_(cby_0__1__1_chany_out_96_[0]),
		.chany_out_97_(cby_0__1__1_chany_out_97_[0]),
		.chany_out_98_(cby_0__1__1_chany_out_98_[0]),
		.chany_out_99_(cby_0__1__1_chany_out_99_[0]),
		.chany_out_100_(cby_0__1__1_chany_out_100_[0]),
		.chany_out_101_(cby_0__1__1_chany_out_101_[0]),
		.chany_out_102_(cby_0__1__1_chany_out_102_[0]),
		.chany_out_103_(cby_0__1__1_chany_out_103_[0]),
		.chany_out_104_(cby_0__1__1_chany_out_104_[0]),
		.chany_out_105_(cby_0__1__1_chany_out_105_[0]),
		.chany_out_106_(cby_0__1__1_chany_out_106_[0]),
		.chany_out_107_(cby_0__1__1_chany_out_107_[0]),
		.chany_out_108_(cby_0__1__1_chany_out_108_[0]),
		.chany_out_109_(cby_0__1__1_chany_out_109_[0]),
		.chany_out_110_(cby_0__1__1_chany_out_110_[0]),
		.chany_out_111_(cby_0__1__1_chany_out_111_[0]),
		.chany_out_112_(cby_0__1__1_chany_out_112_[0]),
		.chany_out_113_(cby_0__1__1_chany_out_113_[0]),
		.chany_out_114_(cby_0__1__1_chany_out_114_[0]),
		.chany_out_115_(cby_0__1__1_chany_out_115_[0]),
		.chany_out_116_(cby_0__1__1_chany_out_116_[0]),
		.chany_out_117_(cby_0__1__1_chany_out_117_[0]),
		.chany_out_118_(cby_0__1__1_chany_out_118_[0]),
		.chany_out_119_(cby_0__1__1_chany_out_119_[0]),
		.chany_out_120_(cby_0__1__1_chany_out_120_[0]),
		.chany_out_121_(cby_0__1__1_chany_out_121_[0]),
		.chany_out_122_(cby_0__1__1_chany_out_122_[0]),
		.chany_out_123_(cby_0__1__1_chany_out_123_[0]),
		.chany_out_124_(cby_0__1__1_chany_out_124_[0]),
		.chany_out_125_(cby_0__1__1_chany_out_125_[0]),
		.chany_out_126_(cby_0__1__1_chany_out_126_[0]),
		.chany_out_127_(cby_0__1__1_chany_out_127_[0]),
		.chany_out_128_(cby_0__1__1_chany_out_128_[0]),
		.chany_out_129_(cby_0__1__1_chany_out_129_[0]),
		.chany_out_130_(cby_0__1__1_chany_out_130_[0]),
		.chany_out_131_(cby_0__1__1_chany_out_131_[0]),
		.chany_out_132_(cby_0__1__1_chany_out_132_[0]),
		.chany_out_133_(cby_0__1__1_chany_out_133_[0]),
		.chany_out_134_(cby_0__1__1_chany_out_134_[0]),
		.chany_out_135_(cby_0__1__1_chany_out_135_[0]),
		.chany_out_136_(cby_0__1__1_chany_out_136_[0]),
		.chany_out_137_(cby_0__1__1_chany_out_137_[0]),
		.chany_out_138_(cby_0__1__1_chany_out_138_[0]),
		.chany_out_139_(cby_0__1__1_chany_out_139_[0]),
		.chany_out_140_(cby_0__1__1_chany_out_140_[0]),
		.chany_out_141_(cby_0__1__1_chany_out_141_[0]),
		.chany_out_142_(cby_0__1__1_chany_out_142_[0]),
		.chany_out_143_(cby_0__1__1_chany_out_143_[0]),
		.chany_out_144_(cby_0__1__1_chany_out_144_[0]),
		.chany_out_145_(cby_0__1__1_chany_out_145_[0]),
		.chany_out_146_(cby_0__1__1_chany_out_146_[0]),
		.chany_out_147_(cby_0__1__1_chany_out_147_[0]),
		.chany_out_148_(cby_0__1__1_chany_out_148_[0]),
		.chany_out_149_(cby_0__1__1_chany_out_149_[0]),
		.chany_out_150_(cby_0__1__1_chany_out_150_[0]),
		.chany_out_151_(cby_0__1__1_chany_out_151_[0]),
		.chany_out_152_(cby_0__1__1_chany_out_152_[0]),
		.chany_out_153_(cby_0__1__1_chany_out_153_[0]),
		.chany_out_154_(cby_0__1__1_chany_out_154_[0]),
		.chany_out_155_(cby_0__1__1_chany_out_155_[0]),
		.chany_out_156_(cby_0__1__1_chany_out_156_[0]),
		.chany_out_157_(cby_0__1__1_chany_out_157_[0]),
		.chany_out_158_(cby_0__1__1_chany_out_158_[0]),
		.chany_out_159_(cby_0__1__1_chany_out_159_[0]),
		.chany_out_160_(cby_0__1__1_chany_out_160_[0]),
		.chany_out_161_(cby_0__1__1_chany_out_161_[0]),
		.chany_out_162_(cby_0__1__1_chany_out_162_[0]),
		.chany_out_163_(cby_0__1__1_chany_out_163_[0]),
		.chany_out_164_(cby_0__1__1_chany_out_164_[0]),
		.chany_out_165_(cby_0__1__1_chany_out_165_[0]),
		.chany_out_166_(cby_0__1__1_chany_out_166_[0]),
		.chany_out_167_(cby_0__1__1_chany_out_167_[0]),
		.chany_out_168_(cby_0__1__1_chany_out_168_[0]),
		.chany_out_169_(cby_0__1__1_chany_out_169_[0]),
		.chany_out_170_(cby_0__1__1_chany_out_170_[0]),
		.chany_out_171_(cby_0__1__1_chany_out_171_[0]),
		.chany_out_172_(cby_0__1__1_chany_out_172_[0]),
		.chany_out_173_(cby_0__1__1_chany_out_173_[0]),
		.chany_out_174_(cby_0__1__1_chany_out_174_[0]),
		.chany_out_175_(cby_0__1__1_chany_out_175_[0]),
		.chany_out_176_(cby_0__1__1_chany_out_176_[0]),
		.chany_out_177_(cby_0__1__1_chany_out_177_[0]),
		.chany_out_178_(cby_0__1__1_chany_out_178_[0]),
		.chany_out_179_(cby_0__1__1_chany_out_179_[0]),
		.chany_out_180_(cby_0__1__1_chany_out_180_[0]),
		.chany_out_181_(cby_0__1__1_chany_out_181_[0]),
		.chany_out_182_(cby_0__1__1_chany_out_182_[0]),
		.chany_out_183_(cby_0__1__1_chany_out_183_[0]),
		.chany_out_184_(cby_0__1__1_chany_out_184_[0]),
		.chany_out_185_(cby_0__1__1_chany_out_185_[0]),
		.chany_out_186_(cby_0__1__1_chany_out_186_[0]),
		.chany_out_187_(cby_0__1__1_chany_out_187_[0]),
		.chany_out_188_(cby_0__1__1_chany_out_188_[0]),
		.chany_out_189_(cby_0__1__1_chany_out_189_[0]),
		.chany_out_190_(cby_0__1__1_chany_out_190_[0]),
		.chany_out_191_(cby_0__1__1_chany_out_191_[0]),
		.chany_out_192_(cby_0__1__1_chany_out_192_[0]),
		.chany_out_193_(cby_0__1__1_chany_out_193_[0]),
		.chany_out_194_(cby_0__1__1_chany_out_194_[0]),
		.chany_out_195_(cby_0__1__1_chany_out_195_[0]),
		.chany_out_196_(cby_0__1__1_chany_out_196_[0]),
		.chany_out_197_(cby_0__1__1_chany_out_197_[0]),
		.chany_out_198_(cby_0__1__1_chany_out_198_[0]),
		.chany_out_199_(cby_0__1__1_chany_out_199_[0]),
		.left_grid_pin_0_(cby_0__1__1_left_grid_pin_0_[0]),
		.ccff_tail(cby_0__1__1_ccff_tail[0]));

	cby_1__1_ cby_1__1_ (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.chany_in_0_(sb_1__0__0_chany_top_out_0_[0]),
		.chany_in_1_(sb_1__1__0_chany_bottom_out_1_[0]),
		.chany_in_2_(sb_1__0__0_chany_top_out_2_[0]),
		.chany_in_3_(sb_1__1__0_chany_bottom_out_3_[0]),
		.chany_in_4_(sb_1__0__0_chany_top_out_4_[0]),
		.chany_in_5_(sb_1__1__0_chany_bottom_out_5_[0]),
		.chany_in_6_(sb_1__0__0_chany_top_out_6_[0]),
		.chany_in_7_(sb_1__1__0_chany_bottom_out_7_[0]),
		.chany_in_8_(sb_1__0__0_chany_top_out_8_[0]),
		.chany_in_9_(sb_1__1__0_chany_bottom_out_9_[0]),
		.chany_in_10_(sb_1__0__0_chany_top_out_10_[0]),
		.chany_in_11_(sb_1__1__0_chany_bottom_out_11_[0]),
		.chany_in_12_(sb_1__0__0_chany_top_out_12_[0]),
		.chany_in_13_(sb_1__1__0_chany_bottom_out_13_[0]),
		.chany_in_14_(sb_1__0__0_chany_top_out_14_[0]),
		.chany_in_15_(sb_1__1__0_chany_bottom_out_15_[0]),
		.chany_in_16_(sb_1__0__0_chany_top_out_16_[0]),
		.chany_in_17_(sb_1__1__0_chany_bottom_out_17_[0]),
		.chany_in_18_(sb_1__0__0_chany_top_out_18_[0]),
		.chany_in_19_(sb_1__1__0_chany_bottom_out_19_[0]),
		.chany_in_20_(sb_1__0__0_chany_top_out_20_[0]),
		.chany_in_21_(sb_1__1__0_chany_bottom_out_21_[0]),
		.chany_in_22_(sb_1__0__0_chany_top_out_22_[0]),
		.chany_in_23_(sb_1__1__0_chany_bottom_out_23_[0]),
		.chany_in_24_(sb_1__0__0_chany_top_out_24_[0]),
		.chany_in_25_(sb_1__1__0_chany_bottom_out_25_[0]),
		.chany_in_26_(sb_1__0__0_chany_top_out_26_[0]),
		.chany_in_27_(sb_1__1__0_chany_bottom_out_27_[0]),
		.chany_in_28_(sb_1__0__0_chany_top_out_28_[0]),
		.chany_in_29_(sb_1__1__0_chany_bottom_out_29_[0]),
		.chany_in_30_(sb_1__0__0_chany_top_out_30_[0]),
		.chany_in_31_(sb_1__1__0_chany_bottom_out_31_[0]),
		.chany_in_32_(sb_1__0__0_chany_top_out_32_[0]),
		.chany_in_33_(sb_1__1__0_chany_bottom_out_33_[0]),
		.chany_in_34_(sb_1__0__0_chany_top_out_34_[0]),
		.chany_in_35_(sb_1__1__0_chany_bottom_out_35_[0]),
		.chany_in_36_(sb_1__0__0_chany_top_out_36_[0]),
		.chany_in_37_(sb_1__1__0_chany_bottom_out_37_[0]),
		.chany_in_38_(sb_1__0__0_chany_top_out_38_[0]),
		.chany_in_39_(sb_1__1__0_chany_bottom_out_39_[0]),
		.chany_in_40_(sb_1__0__0_chany_top_out_40_[0]),
		.chany_in_41_(sb_1__1__0_chany_bottom_out_41_[0]),
		.chany_in_42_(sb_1__0__0_chany_top_out_42_[0]),
		.chany_in_43_(sb_1__1__0_chany_bottom_out_43_[0]),
		.chany_in_44_(sb_1__0__0_chany_top_out_44_[0]),
		.chany_in_45_(sb_1__1__0_chany_bottom_out_45_[0]),
		.chany_in_46_(sb_1__0__0_chany_top_out_46_[0]),
		.chany_in_47_(sb_1__1__0_chany_bottom_out_47_[0]),
		.chany_in_48_(sb_1__0__0_chany_top_out_48_[0]),
		.chany_in_49_(sb_1__1__0_chany_bottom_out_49_[0]),
		.chany_in_50_(sb_1__0__0_chany_top_out_50_[0]),
		.chany_in_51_(sb_1__1__0_chany_bottom_out_51_[0]),
		.chany_in_52_(sb_1__0__0_chany_top_out_52_[0]),
		.chany_in_53_(sb_1__1__0_chany_bottom_out_53_[0]),
		.chany_in_54_(sb_1__0__0_chany_top_out_54_[0]),
		.chany_in_55_(sb_1__1__0_chany_bottom_out_55_[0]),
		.chany_in_56_(sb_1__0__0_chany_top_out_56_[0]),
		.chany_in_57_(sb_1__1__0_chany_bottom_out_57_[0]),
		.chany_in_58_(sb_1__0__0_chany_top_out_58_[0]),
		.chany_in_59_(sb_1__1__0_chany_bottom_out_59_[0]),
		.chany_in_60_(sb_1__0__0_chany_top_out_60_[0]),
		.chany_in_61_(sb_1__1__0_chany_bottom_out_61_[0]),
		.chany_in_62_(sb_1__0__0_chany_top_out_62_[0]),
		.chany_in_63_(sb_1__1__0_chany_bottom_out_63_[0]),
		.chany_in_64_(sb_1__0__0_chany_top_out_64_[0]),
		.chany_in_65_(sb_1__1__0_chany_bottom_out_65_[0]),
		.chany_in_66_(sb_1__0__0_chany_top_out_66_[0]),
		.chany_in_67_(sb_1__1__0_chany_bottom_out_67_[0]),
		.chany_in_68_(sb_1__0__0_chany_top_out_68_[0]),
		.chany_in_69_(sb_1__1__0_chany_bottom_out_69_[0]),
		.chany_in_70_(sb_1__0__0_chany_top_out_70_[0]),
		.chany_in_71_(sb_1__1__0_chany_bottom_out_71_[0]),
		.chany_in_72_(sb_1__0__0_chany_top_out_72_[0]),
		.chany_in_73_(sb_1__1__0_chany_bottom_out_73_[0]),
		.chany_in_74_(sb_1__0__0_chany_top_out_74_[0]),
		.chany_in_75_(sb_1__1__0_chany_bottom_out_75_[0]),
		.chany_in_76_(sb_1__0__0_chany_top_out_76_[0]),
		.chany_in_77_(sb_1__1__0_chany_bottom_out_77_[0]),
		.chany_in_78_(sb_1__0__0_chany_top_out_78_[0]),
		.chany_in_79_(sb_1__1__0_chany_bottom_out_79_[0]),
		.chany_in_80_(sb_1__0__0_chany_top_out_80_[0]),
		.chany_in_81_(sb_1__1__0_chany_bottom_out_81_[0]),
		.chany_in_82_(sb_1__0__0_chany_top_out_82_[0]),
		.chany_in_83_(sb_1__1__0_chany_bottom_out_83_[0]),
		.chany_in_84_(sb_1__0__0_chany_top_out_84_[0]),
		.chany_in_85_(sb_1__1__0_chany_bottom_out_85_[0]),
		.chany_in_86_(sb_1__0__0_chany_top_out_86_[0]),
		.chany_in_87_(sb_1__1__0_chany_bottom_out_87_[0]),
		.chany_in_88_(sb_1__0__0_chany_top_out_88_[0]),
		.chany_in_89_(sb_1__1__0_chany_bottom_out_89_[0]),
		.chany_in_90_(sb_1__0__0_chany_top_out_90_[0]),
		.chany_in_91_(sb_1__1__0_chany_bottom_out_91_[0]),
		.chany_in_92_(sb_1__0__0_chany_top_out_92_[0]),
		.chany_in_93_(sb_1__1__0_chany_bottom_out_93_[0]),
		.chany_in_94_(sb_1__0__0_chany_top_out_94_[0]),
		.chany_in_95_(sb_1__1__0_chany_bottom_out_95_[0]),
		.chany_in_96_(sb_1__0__0_chany_top_out_96_[0]),
		.chany_in_97_(sb_1__1__0_chany_bottom_out_97_[0]),
		.chany_in_98_(sb_1__0__0_chany_top_out_98_[0]),
		.chany_in_99_(sb_1__1__0_chany_bottom_out_99_[0]),
		.chany_in_100_(sb_1__0__0_chany_top_out_100_[0]),
		.chany_in_101_(sb_1__1__0_chany_bottom_out_101_[0]),
		.chany_in_102_(sb_1__0__0_chany_top_out_102_[0]),
		.chany_in_103_(sb_1__1__0_chany_bottom_out_103_[0]),
		.chany_in_104_(sb_1__0__0_chany_top_out_104_[0]),
		.chany_in_105_(sb_1__1__0_chany_bottom_out_105_[0]),
		.chany_in_106_(sb_1__0__0_chany_top_out_106_[0]),
		.chany_in_107_(sb_1__1__0_chany_bottom_out_107_[0]),
		.chany_in_108_(sb_1__0__0_chany_top_out_108_[0]),
		.chany_in_109_(sb_1__1__0_chany_bottom_out_109_[0]),
		.chany_in_110_(sb_1__0__0_chany_top_out_110_[0]),
		.chany_in_111_(sb_1__1__0_chany_bottom_out_111_[0]),
		.chany_in_112_(sb_1__0__0_chany_top_out_112_[0]),
		.chany_in_113_(sb_1__1__0_chany_bottom_out_113_[0]),
		.chany_in_114_(sb_1__0__0_chany_top_out_114_[0]),
		.chany_in_115_(sb_1__1__0_chany_bottom_out_115_[0]),
		.chany_in_116_(sb_1__0__0_chany_top_out_116_[0]),
		.chany_in_117_(sb_1__1__0_chany_bottom_out_117_[0]),
		.chany_in_118_(sb_1__0__0_chany_top_out_118_[0]),
		.chany_in_119_(sb_1__1__0_chany_bottom_out_119_[0]),
		.chany_in_120_(sb_1__0__0_chany_top_out_120_[0]),
		.chany_in_121_(sb_1__1__0_chany_bottom_out_121_[0]),
		.chany_in_122_(sb_1__0__0_chany_top_out_122_[0]),
		.chany_in_123_(sb_1__1__0_chany_bottom_out_123_[0]),
		.chany_in_124_(sb_1__0__0_chany_top_out_124_[0]),
		.chany_in_125_(sb_1__1__0_chany_bottom_out_125_[0]),
		.chany_in_126_(sb_1__0__0_chany_top_out_126_[0]),
		.chany_in_127_(sb_1__1__0_chany_bottom_out_127_[0]),
		.chany_in_128_(sb_1__0__0_chany_top_out_128_[0]),
		.chany_in_129_(sb_1__1__0_chany_bottom_out_129_[0]),
		.chany_in_130_(sb_1__0__0_chany_top_out_130_[0]),
		.chany_in_131_(sb_1__1__0_chany_bottom_out_131_[0]),
		.chany_in_132_(sb_1__0__0_chany_top_out_132_[0]),
		.chany_in_133_(sb_1__1__0_chany_bottom_out_133_[0]),
		.chany_in_134_(sb_1__0__0_chany_top_out_134_[0]),
		.chany_in_135_(sb_1__1__0_chany_bottom_out_135_[0]),
		.chany_in_136_(sb_1__0__0_chany_top_out_136_[0]),
		.chany_in_137_(sb_1__1__0_chany_bottom_out_137_[0]),
		.chany_in_138_(sb_1__0__0_chany_top_out_138_[0]),
		.chany_in_139_(sb_1__1__0_chany_bottom_out_139_[0]),
		.chany_in_140_(sb_1__0__0_chany_top_out_140_[0]),
		.chany_in_141_(sb_1__1__0_chany_bottom_out_141_[0]),
		.chany_in_142_(sb_1__0__0_chany_top_out_142_[0]),
		.chany_in_143_(sb_1__1__0_chany_bottom_out_143_[0]),
		.chany_in_144_(sb_1__0__0_chany_top_out_144_[0]),
		.chany_in_145_(sb_1__1__0_chany_bottom_out_145_[0]),
		.chany_in_146_(sb_1__0__0_chany_top_out_146_[0]),
		.chany_in_147_(sb_1__1__0_chany_bottom_out_147_[0]),
		.chany_in_148_(sb_1__0__0_chany_top_out_148_[0]),
		.chany_in_149_(sb_1__1__0_chany_bottom_out_149_[0]),
		.chany_in_150_(sb_1__0__0_chany_top_out_150_[0]),
		.chany_in_151_(sb_1__1__0_chany_bottom_out_151_[0]),
		.chany_in_152_(sb_1__0__0_chany_top_out_152_[0]),
		.chany_in_153_(sb_1__1__0_chany_bottom_out_153_[0]),
		.chany_in_154_(sb_1__0__0_chany_top_out_154_[0]),
		.chany_in_155_(sb_1__1__0_chany_bottom_out_155_[0]),
		.chany_in_156_(sb_1__0__0_chany_top_out_156_[0]),
		.chany_in_157_(sb_1__1__0_chany_bottom_out_157_[0]),
		.chany_in_158_(sb_1__0__0_chany_top_out_158_[0]),
		.chany_in_159_(sb_1__1__0_chany_bottom_out_159_[0]),
		.chany_in_160_(sb_1__0__0_chany_top_out_160_[0]),
		.chany_in_161_(sb_1__1__0_chany_bottom_out_161_[0]),
		.chany_in_162_(sb_1__0__0_chany_top_out_162_[0]),
		.chany_in_163_(sb_1__1__0_chany_bottom_out_163_[0]),
		.chany_in_164_(sb_1__0__0_chany_top_out_164_[0]),
		.chany_in_165_(sb_1__1__0_chany_bottom_out_165_[0]),
		.chany_in_166_(sb_1__0__0_chany_top_out_166_[0]),
		.chany_in_167_(sb_1__1__0_chany_bottom_out_167_[0]),
		.chany_in_168_(sb_1__0__0_chany_top_out_168_[0]),
		.chany_in_169_(sb_1__1__0_chany_bottom_out_169_[0]),
		.chany_in_170_(sb_1__0__0_chany_top_out_170_[0]),
		.chany_in_171_(sb_1__1__0_chany_bottom_out_171_[0]),
		.chany_in_172_(sb_1__0__0_chany_top_out_172_[0]),
		.chany_in_173_(sb_1__1__0_chany_bottom_out_173_[0]),
		.chany_in_174_(sb_1__0__0_chany_top_out_174_[0]),
		.chany_in_175_(sb_1__1__0_chany_bottom_out_175_[0]),
		.chany_in_176_(sb_1__0__0_chany_top_out_176_[0]),
		.chany_in_177_(sb_1__1__0_chany_bottom_out_177_[0]),
		.chany_in_178_(sb_1__0__0_chany_top_out_178_[0]),
		.chany_in_179_(sb_1__1__0_chany_bottom_out_179_[0]),
		.chany_in_180_(sb_1__0__0_chany_top_out_180_[0]),
		.chany_in_181_(sb_1__1__0_chany_bottom_out_181_[0]),
		.chany_in_182_(sb_1__0__0_chany_top_out_182_[0]),
		.chany_in_183_(sb_1__1__0_chany_bottom_out_183_[0]),
		.chany_in_184_(sb_1__0__0_chany_top_out_184_[0]),
		.chany_in_185_(sb_1__1__0_chany_bottom_out_185_[0]),
		.chany_in_186_(sb_1__0__0_chany_top_out_186_[0]),
		.chany_in_187_(sb_1__1__0_chany_bottom_out_187_[0]),
		.chany_in_188_(sb_1__0__0_chany_top_out_188_[0]),
		.chany_in_189_(sb_1__1__0_chany_bottom_out_189_[0]),
		.chany_in_190_(sb_1__0__0_chany_top_out_190_[0]),
		.chany_in_191_(sb_1__1__0_chany_bottom_out_191_[0]),
		.chany_in_192_(sb_1__0__0_chany_top_out_192_[0]),
		.chany_in_193_(sb_1__1__0_chany_bottom_out_193_[0]),
		.chany_in_194_(sb_1__0__0_chany_top_out_194_[0]),
		.chany_in_195_(sb_1__1__0_chany_bottom_out_195_[0]),
		.chany_in_196_(sb_1__0__0_chany_top_out_196_[0]),
		.chany_in_197_(sb_1__1__0_chany_bottom_out_197_[0]),
		.chany_in_198_(sb_1__0__0_chany_top_out_198_[0]),
		.chany_in_199_(sb_1__1__0_chany_bottom_out_199_[0]),
		.ccff_head(cbx_1__0__0_ccff_tail[0]),
		.chany_out_0_(cby_1__1__0_chany_out_0_[0]),
		.chany_out_1_(cby_1__1__0_chany_out_1_[0]),
		.chany_out_2_(cby_1__1__0_chany_out_2_[0]),
		.chany_out_3_(cby_1__1__0_chany_out_3_[0]),
		.chany_out_4_(cby_1__1__0_chany_out_4_[0]),
		.chany_out_5_(cby_1__1__0_chany_out_5_[0]),
		.chany_out_6_(cby_1__1__0_chany_out_6_[0]),
		.chany_out_7_(cby_1__1__0_chany_out_7_[0]),
		.chany_out_8_(cby_1__1__0_chany_out_8_[0]),
		.chany_out_9_(cby_1__1__0_chany_out_9_[0]),
		.chany_out_10_(cby_1__1__0_chany_out_10_[0]),
		.chany_out_11_(cby_1__1__0_chany_out_11_[0]),
		.chany_out_12_(cby_1__1__0_chany_out_12_[0]),
		.chany_out_13_(cby_1__1__0_chany_out_13_[0]),
		.chany_out_14_(cby_1__1__0_chany_out_14_[0]),
		.chany_out_15_(cby_1__1__0_chany_out_15_[0]),
		.chany_out_16_(cby_1__1__0_chany_out_16_[0]),
		.chany_out_17_(cby_1__1__0_chany_out_17_[0]),
		.chany_out_18_(cby_1__1__0_chany_out_18_[0]),
		.chany_out_19_(cby_1__1__0_chany_out_19_[0]),
		.chany_out_20_(cby_1__1__0_chany_out_20_[0]),
		.chany_out_21_(cby_1__1__0_chany_out_21_[0]),
		.chany_out_22_(cby_1__1__0_chany_out_22_[0]),
		.chany_out_23_(cby_1__1__0_chany_out_23_[0]),
		.chany_out_24_(cby_1__1__0_chany_out_24_[0]),
		.chany_out_25_(cby_1__1__0_chany_out_25_[0]),
		.chany_out_26_(cby_1__1__0_chany_out_26_[0]),
		.chany_out_27_(cby_1__1__0_chany_out_27_[0]),
		.chany_out_28_(cby_1__1__0_chany_out_28_[0]),
		.chany_out_29_(cby_1__1__0_chany_out_29_[0]),
		.chany_out_30_(cby_1__1__0_chany_out_30_[0]),
		.chany_out_31_(cby_1__1__0_chany_out_31_[0]),
		.chany_out_32_(cby_1__1__0_chany_out_32_[0]),
		.chany_out_33_(cby_1__1__0_chany_out_33_[0]),
		.chany_out_34_(cby_1__1__0_chany_out_34_[0]),
		.chany_out_35_(cby_1__1__0_chany_out_35_[0]),
		.chany_out_36_(cby_1__1__0_chany_out_36_[0]),
		.chany_out_37_(cby_1__1__0_chany_out_37_[0]),
		.chany_out_38_(cby_1__1__0_chany_out_38_[0]),
		.chany_out_39_(cby_1__1__0_chany_out_39_[0]),
		.chany_out_40_(cby_1__1__0_chany_out_40_[0]),
		.chany_out_41_(cby_1__1__0_chany_out_41_[0]),
		.chany_out_42_(cby_1__1__0_chany_out_42_[0]),
		.chany_out_43_(cby_1__1__0_chany_out_43_[0]),
		.chany_out_44_(cby_1__1__0_chany_out_44_[0]),
		.chany_out_45_(cby_1__1__0_chany_out_45_[0]),
		.chany_out_46_(cby_1__1__0_chany_out_46_[0]),
		.chany_out_47_(cby_1__1__0_chany_out_47_[0]),
		.chany_out_48_(cby_1__1__0_chany_out_48_[0]),
		.chany_out_49_(cby_1__1__0_chany_out_49_[0]),
		.chany_out_50_(cby_1__1__0_chany_out_50_[0]),
		.chany_out_51_(cby_1__1__0_chany_out_51_[0]),
		.chany_out_52_(cby_1__1__0_chany_out_52_[0]),
		.chany_out_53_(cby_1__1__0_chany_out_53_[0]),
		.chany_out_54_(cby_1__1__0_chany_out_54_[0]),
		.chany_out_55_(cby_1__1__0_chany_out_55_[0]),
		.chany_out_56_(cby_1__1__0_chany_out_56_[0]),
		.chany_out_57_(cby_1__1__0_chany_out_57_[0]),
		.chany_out_58_(cby_1__1__0_chany_out_58_[0]),
		.chany_out_59_(cby_1__1__0_chany_out_59_[0]),
		.chany_out_60_(cby_1__1__0_chany_out_60_[0]),
		.chany_out_61_(cby_1__1__0_chany_out_61_[0]),
		.chany_out_62_(cby_1__1__0_chany_out_62_[0]),
		.chany_out_63_(cby_1__1__0_chany_out_63_[0]),
		.chany_out_64_(cby_1__1__0_chany_out_64_[0]),
		.chany_out_65_(cby_1__1__0_chany_out_65_[0]),
		.chany_out_66_(cby_1__1__0_chany_out_66_[0]),
		.chany_out_67_(cby_1__1__0_chany_out_67_[0]),
		.chany_out_68_(cby_1__1__0_chany_out_68_[0]),
		.chany_out_69_(cby_1__1__0_chany_out_69_[0]),
		.chany_out_70_(cby_1__1__0_chany_out_70_[0]),
		.chany_out_71_(cby_1__1__0_chany_out_71_[0]),
		.chany_out_72_(cby_1__1__0_chany_out_72_[0]),
		.chany_out_73_(cby_1__1__0_chany_out_73_[0]),
		.chany_out_74_(cby_1__1__0_chany_out_74_[0]),
		.chany_out_75_(cby_1__1__0_chany_out_75_[0]),
		.chany_out_76_(cby_1__1__0_chany_out_76_[0]),
		.chany_out_77_(cby_1__1__0_chany_out_77_[0]),
		.chany_out_78_(cby_1__1__0_chany_out_78_[0]),
		.chany_out_79_(cby_1__1__0_chany_out_79_[0]),
		.chany_out_80_(cby_1__1__0_chany_out_80_[0]),
		.chany_out_81_(cby_1__1__0_chany_out_81_[0]),
		.chany_out_82_(cby_1__1__0_chany_out_82_[0]),
		.chany_out_83_(cby_1__1__0_chany_out_83_[0]),
		.chany_out_84_(cby_1__1__0_chany_out_84_[0]),
		.chany_out_85_(cby_1__1__0_chany_out_85_[0]),
		.chany_out_86_(cby_1__1__0_chany_out_86_[0]),
		.chany_out_87_(cby_1__1__0_chany_out_87_[0]),
		.chany_out_88_(cby_1__1__0_chany_out_88_[0]),
		.chany_out_89_(cby_1__1__0_chany_out_89_[0]),
		.chany_out_90_(cby_1__1__0_chany_out_90_[0]),
		.chany_out_91_(cby_1__1__0_chany_out_91_[0]),
		.chany_out_92_(cby_1__1__0_chany_out_92_[0]),
		.chany_out_93_(cby_1__1__0_chany_out_93_[0]),
		.chany_out_94_(cby_1__1__0_chany_out_94_[0]),
		.chany_out_95_(cby_1__1__0_chany_out_95_[0]),
		.chany_out_96_(cby_1__1__0_chany_out_96_[0]),
		.chany_out_97_(cby_1__1__0_chany_out_97_[0]),
		.chany_out_98_(cby_1__1__0_chany_out_98_[0]),
		.chany_out_99_(cby_1__1__0_chany_out_99_[0]),
		.chany_out_100_(cby_1__1__0_chany_out_100_[0]),
		.chany_out_101_(cby_1__1__0_chany_out_101_[0]),
		.chany_out_102_(cby_1__1__0_chany_out_102_[0]),
		.chany_out_103_(cby_1__1__0_chany_out_103_[0]),
		.chany_out_104_(cby_1__1__0_chany_out_104_[0]),
		.chany_out_105_(cby_1__1__0_chany_out_105_[0]),
		.chany_out_106_(cby_1__1__0_chany_out_106_[0]),
		.chany_out_107_(cby_1__1__0_chany_out_107_[0]),
		.chany_out_108_(cby_1__1__0_chany_out_108_[0]),
		.chany_out_109_(cby_1__1__0_chany_out_109_[0]),
		.chany_out_110_(cby_1__1__0_chany_out_110_[0]),
		.chany_out_111_(cby_1__1__0_chany_out_111_[0]),
		.chany_out_112_(cby_1__1__0_chany_out_112_[0]),
		.chany_out_113_(cby_1__1__0_chany_out_113_[0]),
		.chany_out_114_(cby_1__1__0_chany_out_114_[0]),
		.chany_out_115_(cby_1__1__0_chany_out_115_[0]),
		.chany_out_116_(cby_1__1__0_chany_out_116_[0]),
		.chany_out_117_(cby_1__1__0_chany_out_117_[0]),
		.chany_out_118_(cby_1__1__0_chany_out_118_[0]),
		.chany_out_119_(cby_1__1__0_chany_out_119_[0]),
		.chany_out_120_(cby_1__1__0_chany_out_120_[0]),
		.chany_out_121_(cby_1__1__0_chany_out_121_[0]),
		.chany_out_122_(cby_1__1__0_chany_out_122_[0]),
		.chany_out_123_(cby_1__1__0_chany_out_123_[0]),
		.chany_out_124_(cby_1__1__0_chany_out_124_[0]),
		.chany_out_125_(cby_1__1__0_chany_out_125_[0]),
		.chany_out_126_(cby_1__1__0_chany_out_126_[0]),
		.chany_out_127_(cby_1__1__0_chany_out_127_[0]),
		.chany_out_128_(cby_1__1__0_chany_out_128_[0]),
		.chany_out_129_(cby_1__1__0_chany_out_129_[0]),
		.chany_out_130_(cby_1__1__0_chany_out_130_[0]),
		.chany_out_131_(cby_1__1__0_chany_out_131_[0]),
		.chany_out_132_(cby_1__1__0_chany_out_132_[0]),
		.chany_out_133_(cby_1__1__0_chany_out_133_[0]),
		.chany_out_134_(cby_1__1__0_chany_out_134_[0]),
		.chany_out_135_(cby_1__1__0_chany_out_135_[0]),
		.chany_out_136_(cby_1__1__0_chany_out_136_[0]),
		.chany_out_137_(cby_1__1__0_chany_out_137_[0]),
		.chany_out_138_(cby_1__1__0_chany_out_138_[0]),
		.chany_out_139_(cby_1__1__0_chany_out_139_[0]),
		.chany_out_140_(cby_1__1__0_chany_out_140_[0]),
		.chany_out_141_(cby_1__1__0_chany_out_141_[0]),
		.chany_out_142_(cby_1__1__0_chany_out_142_[0]),
		.chany_out_143_(cby_1__1__0_chany_out_143_[0]),
		.chany_out_144_(cby_1__1__0_chany_out_144_[0]),
		.chany_out_145_(cby_1__1__0_chany_out_145_[0]),
		.chany_out_146_(cby_1__1__0_chany_out_146_[0]),
		.chany_out_147_(cby_1__1__0_chany_out_147_[0]),
		.chany_out_148_(cby_1__1__0_chany_out_148_[0]),
		.chany_out_149_(cby_1__1__0_chany_out_149_[0]),
		.chany_out_150_(cby_1__1__0_chany_out_150_[0]),
		.chany_out_151_(cby_1__1__0_chany_out_151_[0]),
		.chany_out_152_(cby_1__1__0_chany_out_152_[0]),
		.chany_out_153_(cby_1__1__0_chany_out_153_[0]),
		.chany_out_154_(cby_1__1__0_chany_out_154_[0]),
		.chany_out_155_(cby_1__1__0_chany_out_155_[0]),
		.chany_out_156_(cby_1__1__0_chany_out_156_[0]),
		.chany_out_157_(cby_1__1__0_chany_out_157_[0]),
		.chany_out_158_(cby_1__1__0_chany_out_158_[0]),
		.chany_out_159_(cby_1__1__0_chany_out_159_[0]),
		.chany_out_160_(cby_1__1__0_chany_out_160_[0]),
		.chany_out_161_(cby_1__1__0_chany_out_161_[0]),
		.chany_out_162_(cby_1__1__0_chany_out_162_[0]),
		.chany_out_163_(cby_1__1__0_chany_out_163_[0]),
		.chany_out_164_(cby_1__1__0_chany_out_164_[0]),
		.chany_out_165_(cby_1__1__0_chany_out_165_[0]),
		.chany_out_166_(cby_1__1__0_chany_out_166_[0]),
		.chany_out_167_(cby_1__1__0_chany_out_167_[0]),
		.chany_out_168_(cby_1__1__0_chany_out_168_[0]),
		.chany_out_169_(cby_1__1__0_chany_out_169_[0]),
		.chany_out_170_(cby_1__1__0_chany_out_170_[0]),
		.chany_out_171_(cby_1__1__0_chany_out_171_[0]),
		.chany_out_172_(cby_1__1__0_chany_out_172_[0]),
		.chany_out_173_(cby_1__1__0_chany_out_173_[0]),
		.chany_out_174_(cby_1__1__0_chany_out_174_[0]),
		.chany_out_175_(cby_1__1__0_chany_out_175_[0]),
		.chany_out_176_(cby_1__1__0_chany_out_176_[0]),
		.chany_out_177_(cby_1__1__0_chany_out_177_[0]),
		.chany_out_178_(cby_1__1__0_chany_out_178_[0]),
		.chany_out_179_(cby_1__1__0_chany_out_179_[0]),
		.chany_out_180_(cby_1__1__0_chany_out_180_[0]),
		.chany_out_181_(cby_1__1__0_chany_out_181_[0]),
		.chany_out_182_(cby_1__1__0_chany_out_182_[0]),
		.chany_out_183_(cby_1__1__0_chany_out_183_[0]),
		.chany_out_184_(cby_1__1__0_chany_out_184_[0]),
		.chany_out_185_(cby_1__1__0_chany_out_185_[0]),
		.chany_out_186_(cby_1__1__0_chany_out_186_[0]),
		.chany_out_187_(cby_1__1__0_chany_out_187_[0]),
		.chany_out_188_(cby_1__1__0_chany_out_188_[0]),
		.chany_out_189_(cby_1__1__0_chany_out_189_[0]),
		.chany_out_190_(cby_1__1__0_chany_out_190_[0]),
		.chany_out_191_(cby_1__1__0_chany_out_191_[0]),
		.chany_out_192_(cby_1__1__0_chany_out_192_[0]),
		.chany_out_193_(cby_1__1__0_chany_out_193_[0]),
		.chany_out_194_(cby_1__1__0_chany_out_194_[0]),
		.chany_out_195_(cby_1__1__0_chany_out_195_[0]),
		.chany_out_196_(cby_1__1__0_chany_out_196_[0]),
		.chany_out_197_(cby_1__1__0_chany_out_197_[0]),
		.chany_out_198_(cby_1__1__0_chany_out_198_[0]),
		.chany_out_199_(cby_1__1__0_chany_out_199_[0]),
		.left_grid_pin_0_(cby_1__1__0_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__0_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__0_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__0_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__0_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__0_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__0_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__0_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__0_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__0_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__0_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__0_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__0_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__0_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__0_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__0_left_grid_pin_15_[0]),
		.left_grid_pin_16_(cby_1__1__0_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__0_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__0_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__0_left_grid_pin_19_[0]),
		.ccff_tail(cby_1__1__0_ccff_tail[0]));

	cby_1__1_ cby_1__2_ (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.chany_in_0_(sb_1__1__0_chany_top_out_0_[0]),
		.chany_in_1_(sb_1__2__0_chany_bottom_out_1_[0]),
		.chany_in_2_(sb_1__1__0_chany_top_out_2_[0]),
		.chany_in_3_(sb_1__2__0_chany_bottom_out_3_[0]),
		.chany_in_4_(sb_1__1__0_chany_top_out_4_[0]),
		.chany_in_5_(sb_1__2__0_chany_bottom_out_5_[0]),
		.chany_in_6_(sb_1__1__0_chany_top_out_6_[0]),
		.chany_in_7_(sb_1__2__0_chany_bottom_out_7_[0]),
		.chany_in_8_(sb_1__1__0_chany_top_out_8_[0]),
		.chany_in_9_(sb_1__2__0_chany_bottom_out_9_[0]),
		.chany_in_10_(sb_1__1__0_chany_top_out_10_[0]),
		.chany_in_11_(sb_1__2__0_chany_bottom_out_11_[0]),
		.chany_in_12_(sb_1__1__0_chany_top_out_12_[0]),
		.chany_in_13_(sb_1__2__0_chany_bottom_out_13_[0]),
		.chany_in_14_(sb_1__1__0_chany_top_out_14_[0]),
		.chany_in_15_(sb_1__2__0_chany_bottom_out_15_[0]),
		.chany_in_16_(sb_1__1__0_chany_top_out_16_[0]),
		.chany_in_17_(sb_1__2__0_chany_bottom_out_17_[0]),
		.chany_in_18_(sb_1__1__0_chany_top_out_18_[0]),
		.chany_in_19_(sb_1__2__0_chany_bottom_out_19_[0]),
		.chany_in_20_(sb_1__1__0_chany_top_out_20_[0]),
		.chany_in_21_(sb_1__2__0_chany_bottom_out_21_[0]),
		.chany_in_22_(sb_1__1__0_chany_top_out_22_[0]),
		.chany_in_23_(sb_1__2__0_chany_bottom_out_23_[0]),
		.chany_in_24_(sb_1__1__0_chany_top_out_24_[0]),
		.chany_in_25_(sb_1__2__0_chany_bottom_out_25_[0]),
		.chany_in_26_(sb_1__1__0_chany_top_out_26_[0]),
		.chany_in_27_(sb_1__2__0_chany_bottom_out_27_[0]),
		.chany_in_28_(sb_1__1__0_chany_top_out_28_[0]),
		.chany_in_29_(sb_1__2__0_chany_bottom_out_29_[0]),
		.chany_in_30_(sb_1__1__0_chany_top_out_30_[0]),
		.chany_in_31_(sb_1__2__0_chany_bottom_out_31_[0]),
		.chany_in_32_(sb_1__1__0_chany_top_out_32_[0]),
		.chany_in_33_(sb_1__2__0_chany_bottom_out_33_[0]),
		.chany_in_34_(sb_1__1__0_chany_top_out_34_[0]),
		.chany_in_35_(sb_1__2__0_chany_bottom_out_35_[0]),
		.chany_in_36_(sb_1__1__0_chany_top_out_36_[0]),
		.chany_in_37_(sb_1__2__0_chany_bottom_out_37_[0]),
		.chany_in_38_(sb_1__1__0_chany_top_out_38_[0]),
		.chany_in_39_(sb_1__2__0_chany_bottom_out_39_[0]),
		.chany_in_40_(sb_1__1__0_chany_top_out_40_[0]),
		.chany_in_41_(sb_1__2__0_chany_bottom_out_41_[0]),
		.chany_in_42_(sb_1__1__0_chany_top_out_42_[0]),
		.chany_in_43_(sb_1__2__0_chany_bottom_out_43_[0]),
		.chany_in_44_(sb_1__1__0_chany_top_out_44_[0]),
		.chany_in_45_(sb_1__2__0_chany_bottom_out_45_[0]),
		.chany_in_46_(sb_1__1__0_chany_top_out_46_[0]),
		.chany_in_47_(sb_1__2__0_chany_bottom_out_47_[0]),
		.chany_in_48_(sb_1__1__0_chany_top_out_48_[0]),
		.chany_in_49_(sb_1__2__0_chany_bottom_out_49_[0]),
		.chany_in_50_(sb_1__1__0_chany_top_out_50_[0]),
		.chany_in_51_(sb_1__2__0_chany_bottom_out_51_[0]),
		.chany_in_52_(sb_1__1__0_chany_top_out_52_[0]),
		.chany_in_53_(sb_1__2__0_chany_bottom_out_53_[0]),
		.chany_in_54_(sb_1__1__0_chany_top_out_54_[0]),
		.chany_in_55_(sb_1__2__0_chany_bottom_out_55_[0]),
		.chany_in_56_(sb_1__1__0_chany_top_out_56_[0]),
		.chany_in_57_(sb_1__2__0_chany_bottom_out_57_[0]),
		.chany_in_58_(sb_1__1__0_chany_top_out_58_[0]),
		.chany_in_59_(sb_1__2__0_chany_bottom_out_59_[0]),
		.chany_in_60_(sb_1__1__0_chany_top_out_60_[0]),
		.chany_in_61_(sb_1__2__0_chany_bottom_out_61_[0]),
		.chany_in_62_(sb_1__1__0_chany_top_out_62_[0]),
		.chany_in_63_(sb_1__2__0_chany_bottom_out_63_[0]),
		.chany_in_64_(sb_1__1__0_chany_top_out_64_[0]),
		.chany_in_65_(sb_1__2__0_chany_bottom_out_65_[0]),
		.chany_in_66_(sb_1__1__0_chany_top_out_66_[0]),
		.chany_in_67_(sb_1__2__0_chany_bottom_out_67_[0]),
		.chany_in_68_(sb_1__1__0_chany_top_out_68_[0]),
		.chany_in_69_(sb_1__2__0_chany_bottom_out_69_[0]),
		.chany_in_70_(sb_1__1__0_chany_top_out_70_[0]),
		.chany_in_71_(sb_1__2__0_chany_bottom_out_71_[0]),
		.chany_in_72_(sb_1__1__0_chany_top_out_72_[0]),
		.chany_in_73_(sb_1__2__0_chany_bottom_out_73_[0]),
		.chany_in_74_(sb_1__1__0_chany_top_out_74_[0]),
		.chany_in_75_(sb_1__2__0_chany_bottom_out_75_[0]),
		.chany_in_76_(sb_1__1__0_chany_top_out_76_[0]),
		.chany_in_77_(sb_1__2__0_chany_bottom_out_77_[0]),
		.chany_in_78_(sb_1__1__0_chany_top_out_78_[0]),
		.chany_in_79_(sb_1__2__0_chany_bottom_out_79_[0]),
		.chany_in_80_(sb_1__1__0_chany_top_out_80_[0]),
		.chany_in_81_(sb_1__2__0_chany_bottom_out_81_[0]),
		.chany_in_82_(sb_1__1__0_chany_top_out_82_[0]),
		.chany_in_83_(sb_1__2__0_chany_bottom_out_83_[0]),
		.chany_in_84_(sb_1__1__0_chany_top_out_84_[0]),
		.chany_in_85_(sb_1__2__0_chany_bottom_out_85_[0]),
		.chany_in_86_(sb_1__1__0_chany_top_out_86_[0]),
		.chany_in_87_(sb_1__2__0_chany_bottom_out_87_[0]),
		.chany_in_88_(sb_1__1__0_chany_top_out_88_[0]),
		.chany_in_89_(sb_1__2__0_chany_bottom_out_89_[0]),
		.chany_in_90_(sb_1__1__0_chany_top_out_90_[0]),
		.chany_in_91_(sb_1__2__0_chany_bottom_out_91_[0]),
		.chany_in_92_(sb_1__1__0_chany_top_out_92_[0]),
		.chany_in_93_(sb_1__2__0_chany_bottom_out_93_[0]),
		.chany_in_94_(sb_1__1__0_chany_top_out_94_[0]),
		.chany_in_95_(sb_1__2__0_chany_bottom_out_95_[0]),
		.chany_in_96_(sb_1__1__0_chany_top_out_96_[0]),
		.chany_in_97_(sb_1__2__0_chany_bottom_out_97_[0]),
		.chany_in_98_(sb_1__1__0_chany_top_out_98_[0]),
		.chany_in_99_(sb_1__2__0_chany_bottom_out_99_[0]),
		.chany_in_100_(sb_1__1__0_chany_top_out_100_[0]),
		.chany_in_101_(sb_1__2__0_chany_bottom_out_101_[0]),
		.chany_in_102_(sb_1__1__0_chany_top_out_102_[0]),
		.chany_in_103_(sb_1__2__0_chany_bottom_out_103_[0]),
		.chany_in_104_(sb_1__1__0_chany_top_out_104_[0]),
		.chany_in_105_(sb_1__2__0_chany_bottom_out_105_[0]),
		.chany_in_106_(sb_1__1__0_chany_top_out_106_[0]),
		.chany_in_107_(sb_1__2__0_chany_bottom_out_107_[0]),
		.chany_in_108_(sb_1__1__0_chany_top_out_108_[0]),
		.chany_in_109_(sb_1__2__0_chany_bottom_out_109_[0]),
		.chany_in_110_(sb_1__1__0_chany_top_out_110_[0]),
		.chany_in_111_(sb_1__2__0_chany_bottom_out_111_[0]),
		.chany_in_112_(sb_1__1__0_chany_top_out_112_[0]),
		.chany_in_113_(sb_1__2__0_chany_bottom_out_113_[0]),
		.chany_in_114_(sb_1__1__0_chany_top_out_114_[0]),
		.chany_in_115_(sb_1__2__0_chany_bottom_out_115_[0]),
		.chany_in_116_(sb_1__1__0_chany_top_out_116_[0]),
		.chany_in_117_(sb_1__2__0_chany_bottom_out_117_[0]),
		.chany_in_118_(sb_1__1__0_chany_top_out_118_[0]),
		.chany_in_119_(sb_1__2__0_chany_bottom_out_119_[0]),
		.chany_in_120_(sb_1__1__0_chany_top_out_120_[0]),
		.chany_in_121_(sb_1__2__0_chany_bottom_out_121_[0]),
		.chany_in_122_(sb_1__1__0_chany_top_out_122_[0]),
		.chany_in_123_(sb_1__2__0_chany_bottom_out_123_[0]),
		.chany_in_124_(sb_1__1__0_chany_top_out_124_[0]),
		.chany_in_125_(sb_1__2__0_chany_bottom_out_125_[0]),
		.chany_in_126_(sb_1__1__0_chany_top_out_126_[0]),
		.chany_in_127_(sb_1__2__0_chany_bottom_out_127_[0]),
		.chany_in_128_(sb_1__1__0_chany_top_out_128_[0]),
		.chany_in_129_(sb_1__2__0_chany_bottom_out_129_[0]),
		.chany_in_130_(sb_1__1__0_chany_top_out_130_[0]),
		.chany_in_131_(sb_1__2__0_chany_bottom_out_131_[0]),
		.chany_in_132_(sb_1__1__0_chany_top_out_132_[0]),
		.chany_in_133_(sb_1__2__0_chany_bottom_out_133_[0]),
		.chany_in_134_(sb_1__1__0_chany_top_out_134_[0]),
		.chany_in_135_(sb_1__2__0_chany_bottom_out_135_[0]),
		.chany_in_136_(sb_1__1__0_chany_top_out_136_[0]),
		.chany_in_137_(sb_1__2__0_chany_bottom_out_137_[0]),
		.chany_in_138_(sb_1__1__0_chany_top_out_138_[0]),
		.chany_in_139_(sb_1__2__0_chany_bottom_out_139_[0]),
		.chany_in_140_(sb_1__1__0_chany_top_out_140_[0]),
		.chany_in_141_(sb_1__2__0_chany_bottom_out_141_[0]),
		.chany_in_142_(sb_1__1__0_chany_top_out_142_[0]),
		.chany_in_143_(sb_1__2__0_chany_bottom_out_143_[0]),
		.chany_in_144_(sb_1__1__0_chany_top_out_144_[0]),
		.chany_in_145_(sb_1__2__0_chany_bottom_out_145_[0]),
		.chany_in_146_(sb_1__1__0_chany_top_out_146_[0]),
		.chany_in_147_(sb_1__2__0_chany_bottom_out_147_[0]),
		.chany_in_148_(sb_1__1__0_chany_top_out_148_[0]),
		.chany_in_149_(sb_1__2__0_chany_bottom_out_149_[0]),
		.chany_in_150_(sb_1__1__0_chany_top_out_150_[0]),
		.chany_in_151_(sb_1__2__0_chany_bottom_out_151_[0]),
		.chany_in_152_(sb_1__1__0_chany_top_out_152_[0]),
		.chany_in_153_(sb_1__2__0_chany_bottom_out_153_[0]),
		.chany_in_154_(sb_1__1__0_chany_top_out_154_[0]),
		.chany_in_155_(sb_1__2__0_chany_bottom_out_155_[0]),
		.chany_in_156_(sb_1__1__0_chany_top_out_156_[0]),
		.chany_in_157_(sb_1__2__0_chany_bottom_out_157_[0]),
		.chany_in_158_(sb_1__1__0_chany_top_out_158_[0]),
		.chany_in_159_(sb_1__2__0_chany_bottom_out_159_[0]),
		.chany_in_160_(sb_1__1__0_chany_top_out_160_[0]),
		.chany_in_161_(sb_1__2__0_chany_bottom_out_161_[0]),
		.chany_in_162_(sb_1__1__0_chany_top_out_162_[0]),
		.chany_in_163_(sb_1__2__0_chany_bottom_out_163_[0]),
		.chany_in_164_(sb_1__1__0_chany_top_out_164_[0]),
		.chany_in_165_(sb_1__2__0_chany_bottom_out_165_[0]),
		.chany_in_166_(sb_1__1__0_chany_top_out_166_[0]),
		.chany_in_167_(sb_1__2__0_chany_bottom_out_167_[0]),
		.chany_in_168_(sb_1__1__0_chany_top_out_168_[0]),
		.chany_in_169_(sb_1__2__0_chany_bottom_out_169_[0]),
		.chany_in_170_(sb_1__1__0_chany_top_out_170_[0]),
		.chany_in_171_(sb_1__2__0_chany_bottom_out_171_[0]),
		.chany_in_172_(sb_1__1__0_chany_top_out_172_[0]),
		.chany_in_173_(sb_1__2__0_chany_bottom_out_173_[0]),
		.chany_in_174_(sb_1__1__0_chany_top_out_174_[0]),
		.chany_in_175_(sb_1__2__0_chany_bottom_out_175_[0]),
		.chany_in_176_(sb_1__1__0_chany_top_out_176_[0]),
		.chany_in_177_(sb_1__2__0_chany_bottom_out_177_[0]),
		.chany_in_178_(sb_1__1__0_chany_top_out_178_[0]),
		.chany_in_179_(sb_1__2__0_chany_bottom_out_179_[0]),
		.chany_in_180_(sb_1__1__0_chany_top_out_180_[0]),
		.chany_in_181_(sb_1__2__0_chany_bottom_out_181_[0]),
		.chany_in_182_(sb_1__1__0_chany_top_out_182_[0]),
		.chany_in_183_(sb_1__2__0_chany_bottom_out_183_[0]),
		.chany_in_184_(sb_1__1__0_chany_top_out_184_[0]),
		.chany_in_185_(sb_1__2__0_chany_bottom_out_185_[0]),
		.chany_in_186_(sb_1__1__0_chany_top_out_186_[0]),
		.chany_in_187_(sb_1__2__0_chany_bottom_out_187_[0]),
		.chany_in_188_(sb_1__1__0_chany_top_out_188_[0]),
		.chany_in_189_(sb_1__2__0_chany_bottom_out_189_[0]),
		.chany_in_190_(sb_1__1__0_chany_top_out_190_[0]),
		.chany_in_191_(sb_1__2__0_chany_bottom_out_191_[0]),
		.chany_in_192_(sb_1__1__0_chany_top_out_192_[0]),
		.chany_in_193_(sb_1__2__0_chany_bottom_out_193_[0]),
		.chany_in_194_(sb_1__1__0_chany_top_out_194_[0]),
		.chany_in_195_(sb_1__2__0_chany_bottom_out_195_[0]),
		.chany_in_196_(sb_1__1__0_chany_top_out_196_[0]),
		.chany_in_197_(sb_1__2__0_chany_bottom_out_197_[0]),
		.chany_in_198_(sb_1__1__0_chany_top_out_198_[0]),
		.chany_in_199_(sb_1__2__0_chany_bottom_out_199_[0]),
		.ccff_head(cbx_1__1__0_ccff_tail[0]),
		.chany_out_0_(cby_1__1__1_chany_out_0_[0]),
		.chany_out_1_(cby_1__1__1_chany_out_1_[0]),
		.chany_out_2_(cby_1__1__1_chany_out_2_[0]),
		.chany_out_3_(cby_1__1__1_chany_out_3_[0]),
		.chany_out_4_(cby_1__1__1_chany_out_4_[0]),
		.chany_out_5_(cby_1__1__1_chany_out_5_[0]),
		.chany_out_6_(cby_1__1__1_chany_out_6_[0]),
		.chany_out_7_(cby_1__1__1_chany_out_7_[0]),
		.chany_out_8_(cby_1__1__1_chany_out_8_[0]),
		.chany_out_9_(cby_1__1__1_chany_out_9_[0]),
		.chany_out_10_(cby_1__1__1_chany_out_10_[0]),
		.chany_out_11_(cby_1__1__1_chany_out_11_[0]),
		.chany_out_12_(cby_1__1__1_chany_out_12_[0]),
		.chany_out_13_(cby_1__1__1_chany_out_13_[0]),
		.chany_out_14_(cby_1__1__1_chany_out_14_[0]),
		.chany_out_15_(cby_1__1__1_chany_out_15_[0]),
		.chany_out_16_(cby_1__1__1_chany_out_16_[0]),
		.chany_out_17_(cby_1__1__1_chany_out_17_[0]),
		.chany_out_18_(cby_1__1__1_chany_out_18_[0]),
		.chany_out_19_(cby_1__1__1_chany_out_19_[0]),
		.chany_out_20_(cby_1__1__1_chany_out_20_[0]),
		.chany_out_21_(cby_1__1__1_chany_out_21_[0]),
		.chany_out_22_(cby_1__1__1_chany_out_22_[0]),
		.chany_out_23_(cby_1__1__1_chany_out_23_[0]),
		.chany_out_24_(cby_1__1__1_chany_out_24_[0]),
		.chany_out_25_(cby_1__1__1_chany_out_25_[0]),
		.chany_out_26_(cby_1__1__1_chany_out_26_[0]),
		.chany_out_27_(cby_1__1__1_chany_out_27_[0]),
		.chany_out_28_(cby_1__1__1_chany_out_28_[0]),
		.chany_out_29_(cby_1__1__1_chany_out_29_[0]),
		.chany_out_30_(cby_1__1__1_chany_out_30_[0]),
		.chany_out_31_(cby_1__1__1_chany_out_31_[0]),
		.chany_out_32_(cby_1__1__1_chany_out_32_[0]),
		.chany_out_33_(cby_1__1__1_chany_out_33_[0]),
		.chany_out_34_(cby_1__1__1_chany_out_34_[0]),
		.chany_out_35_(cby_1__1__1_chany_out_35_[0]),
		.chany_out_36_(cby_1__1__1_chany_out_36_[0]),
		.chany_out_37_(cby_1__1__1_chany_out_37_[0]),
		.chany_out_38_(cby_1__1__1_chany_out_38_[0]),
		.chany_out_39_(cby_1__1__1_chany_out_39_[0]),
		.chany_out_40_(cby_1__1__1_chany_out_40_[0]),
		.chany_out_41_(cby_1__1__1_chany_out_41_[0]),
		.chany_out_42_(cby_1__1__1_chany_out_42_[0]),
		.chany_out_43_(cby_1__1__1_chany_out_43_[0]),
		.chany_out_44_(cby_1__1__1_chany_out_44_[0]),
		.chany_out_45_(cby_1__1__1_chany_out_45_[0]),
		.chany_out_46_(cby_1__1__1_chany_out_46_[0]),
		.chany_out_47_(cby_1__1__1_chany_out_47_[0]),
		.chany_out_48_(cby_1__1__1_chany_out_48_[0]),
		.chany_out_49_(cby_1__1__1_chany_out_49_[0]),
		.chany_out_50_(cby_1__1__1_chany_out_50_[0]),
		.chany_out_51_(cby_1__1__1_chany_out_51_[0]),
		.chany_out_52_(cby_1__1__1_chany_out_52_[0]),
		.chany_out_53_(cby_1__1__1_chany_out_53_[0]),
		.chany_out_54_(cby_1__1__1_chany_out_54_[0]),
		.chany_out_55_(cby_1__1__1_chany_out_55_[0]),
		.chany_out_56_(cby_1__1__1_chany_out_56_[0]),
		.chany_out_57_(cby_1__1__1_chany_out_57_[0]),
		.chany_out_58_(cby_1__1__1_chany_out_58_[0]),
		.chany_out_59_(cby_1__1__1_chany_out_59_[0]),
		.chany_out_60_(cby_1__1__1_chany_out_60_[0]),
		.chany_out_61_(cby_1__1__1_chany_out_61_[0]),
		.chany_out_62_(cby_1__1__1_chany_out_62_[0]),
		.chany_out_63_(cby_1__1__1_chany_out_63_[0]),
		.chany_out_64_(cby_1__1__1_chany_out_64_[0]),
		.chany_out_65_(cby_1__1__1_chany_out_65_[0]),
		.chany_out_66_(cby_1__1__1_chany_out_66_[0]),
		.chany_out_67_(cby_1__1__1_chany_out_67_[0]),
		.chany_out_68_(cby_1__1__1_chany_out_68_[0]),
		.chany_out_69_(cby_1__1__1_chany_out_69_[0]),
		.chany_out_70_(cby_1__1__1_chany_out_70_[0]),
		.chany_out_71_(cby_1__1__1_chany_out_71_[0]),
		.chany_out_72_(cby_1__1__1_chany_out_72_[0]),
		.chany_out_73_(cby_1__1__1_chany_out_73_[0]),
		.chany_out_74_(cby_1__1__1_chany_out_74_[0]),
		.chany_out_75_(cby_1__1__1_chany_out_75_[0]),
		.chany_out_76_(cby_1__1__1_chany_out_76_[0]),
		.chany_out_77_(cby_1__1__1_chany_out_77_[0]),
		.chany_out_78_(cby_1__1__1_chany_out_78_[0]),
		.chany_out_79_(cby_1__1__1_chany_out_79_[0]),
		.chany_out_80_(cby_1__1__1_chany_out_80_[0]),
		.chany_out_81_(cby_1__1__1_chany_out_81_[0]),
		.chany_out_82_(cby_1__1__1_chany_out_82_[0]),
		.chany_out_83_(cby_1__1__1_chany_out_83_[0]),
		.chany_out_84_(cby_1__1__1_chany_out_84_[0]),
		.chany_out_85_(cby_1__1__1_chany_out_85_[0]),
		.chany_out_86_(cby_1__1__1_chany_out_86_[0]),
		.chany_out_87_(cby_1__1__1_chany_out_87_[0]),
		.chany_out_88_(cby_1__1__1_chany_out_88_[0]),
		.chany_out_89_(cby_1__1__1_chany_out_89_[0]),
		.chany_out_90_(cby_1__1__1_chany_out_90_[0]),
		.chany_out_91_(cby_1__1__1_chany_out_91_[0]),
		.chany_out_92_(cby_1__1__1_chany_out_92_[0]),
		.chany_out_93_(cby_1__1__1_chany_out_93_[0]),
		.chany_out_94_(cby_1__1__1_chany_out_94_[0]),
		.chany_out_95_(cby_1__1__1_chany_out_95_[0]),
		.chany_out_96_(cby_1__1__1_chany_out_96_[0]),
		.chany_out_97_(cby_1__1__1_chany_out_97_[0]),
		.chany_out_98_(cby_1__1__1_chany_out_98_[0]),
		.chany_out_99_(cby_1__1__1_chany_out_99_[0]),
		.chany_out_100_(cby_1__1__1_chany_out_100_[0]),
		.chany_out_101_(cby_1__1__1_chany_out_101_[0]),
		.chany_out_102_(cby_1__1__1_chany_out_102_[0]),
		.chany_out_103_(cby_1__1__1_chany_out_103_[0]),
		.chany_out_104_(cby_1__1__1_chany_out_104_[0]),
		.chany_out_105_(cby_1__1__1_chany_out_105_[0]),
		.chany_out_106_(cby_1__1__1_chany_out_106_[0]),
		.chany_out_107_(cby_1__1__1_chany_out_107_[0]),
		.chany_out_108_(cby_1__1__1_chany_out_108_[0]),
		.chany_out_109_(cby_1__1__1_chany_out_109_[0]),
		.chany_out_110_(cby_1__1__1_chany_out_110_[0]),
		.chany_out_111_(cby_1__1__1_chany_out_111_[0]),
		.chany_out_112_(cby_1__1__1_chany_out_112_[0]),
		.chany_out_113_(cby_1__1__1_chany_out_113_[0]),
		.chany_out_114_(cby_1__1__1_chany_out_114_[0]),
		.chany_out_115_(cby_1__1__1_chany_out_115_[0]),
		.chany_out_116_(cby_1__1__1_chany_out_116_[0]),
		.chany_out_117_(cby_1__1__1_chany_out_117_[0]),
		.chany_out_118_(cby_1__1__1_chany_out_118_[0]),
		.chany_out_119_(cby_1__1__1_chany_out_119_[0]),
		.chany_out_120_(cby_1__1__1_chany_out_120_[0]),
		.chany_out_121_(cby_1__1__1_chany_out_121_[0]),
		.chany_out_122_(cby_1__1__1_chany_out_122_[0]),
		.chany_out_123_(cby_1__1__1_chany_out_123_[0]),
		.chany_out_124_(cby_1__1__1_chany_out_124_[0]),
		.chany_out_125_(cby_1__1__1_chany_out_125_[0]),
		.chany_out_126_(cby_1__1__1_chany_out_126_[0]),
		.chany_out_127_(cby_1__1__1_chany_out_127_[0]),
		.chany_out_128_(cby_1__1__1_chany_out_128_[0]),
		.chany_out_129_(cby_1__1__1_chany_out_129_[0]),
		.chany_out_130_(cby_1__1__1_chany_out_130_[0]),
		.chany_out_131_(cby_1__1__1_chany_out_131_[0]),
		.chany_out_132_(cby_1__1__1_chany_out_132_[0]),
		.chany_out_133_(cby_1__1__1_chany_out_133_[0]),
		.chany_out_134_(cby_1__1__1_chany_out_134_[0]),
		.chany_out_135_(cby_1__1__1_chany_out_135_[0]),
		.chany_out_136_(cby_1__1__1_chany_out_136_[0]),
		.chany_out_137_(cby_1__1__1_chany_out_137_[0]),
		.chany_out_138_(cby_1__1__1_chany_out_138_[0]),
		.chany_out_139_(cby_1__1__1_chany_out_139_[0]),
		.chany_out_140_(cby_1__1__1_chany_out_140_[0]),
		.chany_out_141_(cby_1__1__1_chany_out_141_[0]),
		.chany_out_142_(cby_1__1__1_chany_out_142_[0]),
		.chany_out_143_(cby_1__1__1_chany_out_143_[0]),
		.chany_out_144_(cby_1__1__1_chany_out_144_[0]),
		.chany_out_145_(cby_1__1__1_chany_out_145_[0]),
		.chany_out_146_(cby_1__1__1_chany_out_146_[0]),
		.chany_out_147_(cby_1__1__1_chany_out_147_[0]),
		.chany_out_148_(cby_1__1__1_chany_out_148_[0]),
		.chany_out_149_(cby_1__1__1_chany_out_149_[0]),
		.chany_out_150_(cby_1__1__1_chany_out_150_[0]),
		.chany_out_151_(cby_1__1__1_chany_out_151_[0]),
		.chany_out_152_(cby_1__1__1_chany_out_152_[0]),
		.chany_out_153_(cby_1__1__1_chany_out_153_[0]),
		.chany_out_154_(cby_1__1__1_chany_out_154_[0]),
		.chany_out_155_(cby_1__1__1_chany_out_155_[0]),
		.chany_out_156_(cby_1__1__1_chany_out_156_[0]),
		.chany_out_157_(cby_1__1__1_chany_out_157_[0]),
		.chany_out_158_(cby_1__1__1_chany_out_158_[0]),
		.chany_out_159_(cby_1__1__1_chany_out_159_[0]),
		.chany_out_160_(cby_1__1__1_chany_out_160_[0]),
		.chany_out_161_(cby_1__1__1_chany_out_161_[0]),
		.chany_out_162_(cby_1__1__1_chany_out_162_[0]),
		.chany_out_163_(cby_1__1__1_chany_out_163_[0]),
		.chany_out_164_(cby_1__1__1_chany_out_164_[0]),
		.chany_out_165_(cby_1__1__1_chany_out_165_[0]),
		.chany_out_166_(cby_1__1__1_chany_out_166_[0]),
		.chany_out_167_(cby_1__1__1_chany_out_167_[0]),
		.chany_out_168_(cby_1__1__1_chany_out_168_[0]),
		.chany_out_169_(cby_1__1__1_chany_out_169_[0]),
		.chany_out_170_(cby_1__1__1_chany_out_170_[0]),
		.chany_out_171_(cby_1__1__1_chany_out_171_[0]),
		.chany_out_172_(cby_1__1__1_chany_out_172_[0]),
		.chany_out_173_(cby_1__1__1_chany_out_173_[0]),
		.chany_out_174_(cby_1__1__1_chany_out_174_[0]),
		.chany_out_175_(cby_1__1__1_chany_out_175_[0]),
		.chany_out_176_(cby_1__1__1_chany_out_176_[0]),
		.chany_out_177_(cby_1__1__1_chany_out_177_[0]),
		.chany_out_178_(cby_1__1__1_chany_out_178_[0]),
		.chany_out_179_(cby_1__1__1_chany_out_179_[0]),
		.chany_out_180_(cby_1__1__1_chany_out_180_[0]),
		.chany_out_181_(cby_1__1__1_chany_out_181_[0]),
		.chany_out_182_(cby_1__1__1_chany_out_182_[0]),
		.chany_out_183_(cby_1__1__1_chany_out_183_[0]),
		.chany_out_184_(cby_1__1__1_chany_out_184_[0]),
		.chany_out_185_(cby_1__1__1_chany_out_185_[0]),
		.chany_out_186_(cby_1__1__1_chany_out_186_[0]),
		.chany_out_187_(cby_1__1__1_chany_out_187_[0]),
		.chany_out_188_(cby_1__1__1_chany_out_188_[0]),
		.chany_out_189_(cby_1__1__1_chany_out_189_[0]),
		.chany_out_190_(cby_1__1__1_chany_out_190_[0]),
		.chany_out_191_(cby_1__1__1_chany_out_191_[0]),
		.chany_out_192_(cby_1__1__1_chany_out_192_[0]),
		.chany_out_193_(cby_1__1__1_chany_out_193_[0]),
		.chany_out_194_(cby_1__1__1_chany_out_194_[0]),
		.chany_out_195_(cby_1__1__1_chany_out_195_[0]),
		.chany_out_196_(cby_1__1__1_chany_out_196_[0]),
		.chany_out_197_(cby_1__1__1_chany_out_197_[0]),
		.chany_out_198_(cby_1__1__1_chany_out_198_[0]),
		.chany_out_199_(cby_1__1__1_chany_out_199_[0]),
		.left_grid_pin_0_(cby_1__1__1_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__1_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__1_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__1_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__1_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__1_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__1_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__1_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__1_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__1_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__1_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__1_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__1_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__1_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__1_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__1_left_grid_pin_15_[0]),
		.left_grid_pin_16_(cby_1__1__1_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__1_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__1_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__1_left_grid_pin_19_[0]),
		.ccff_tail(cby_1__1__1_ccff_tail[0]));

	cby_2__1_ cby_2__1_ (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.chany_in_0_(sb_2__0__0_chany_top_out_0_[0]),
		.chany_in_1_(sb_2__1__0_chany_bottom_out_1_[0]),
		.chany_in_2_(sb_2__0__0_chany_top_out_2_[0]),
		.chany_in_3_(sb_2__1__0_chany_bottom_out_3_[0]),
		.chany_in_4_(sb_2__0__0_chany_top_out_4_[0]),
		.chany_in_5_(sb_2__1__0_chany_bottom_out_5_[0]),
		.chany_in_6_(sb_2__0__0_chany_top_out_6_[0]),
		.chany_in_7_(sb_2__1__0_chany_bottom_out_7_[0]),
		.chany_in_8_(sb_2__0__0_chany_top_out_8_[0]),
		.chany_in_9_(sb_2__1__0_chany_bottom_out_9_[0]),
		.chany_in_10_(sb_2__0__0_chany_top_out_10_[0]),
		.chany_in_11_(sb_2__1__0_chany_bottom_out_11_[0]),
		.chany_in_12_(sb_2__0__0_chany_top_out_12_[0]),
		.chany_in_13_(sb_2__1__0_chany_bottom_out_13_[0]),
		.chany_in_14_(sb_2__0__0_chany_top_out_14_[0]),
		.chany_in_15_(sb_2__1__0_chany_bottom_out_15_[0]),
		.chany_in_16_(sb_2__0__0_chany_top_out_16_[0]),
		.chany_in_17_(sb_2__1__0_chany_bottom_out_17_[0]),
		.chany_in_18_(sb_2__0__0_chany_top_out_18_[0]),
		.chany_in_19_(sb_2__1__0_chany_bottom_out_19_[0]),
		.chany_in_20_(sb_2__0__0_chany_top_out_20_[0]),
		.chany_in_21_(sb_2__1__0_chany_bottom_out_21_[0]),
		.chany_in_22_(sb_2__0__0_chany_top_out_22_[0]),
		.chany_in_23_(sb_2__1__0_chany_bottom_out_23_[0]),
		.chany_in_24_(sb_2__0__0_chany_top_out_24_[0]),
		.chany_in_25_(sb_2__1__0_chany_bottom_out_25_[0]),
		.chany_in_26_(sb_2__0__0_chany_top_out_26_[0]),
		.chany_in_27_(sb_2__1__0_chany_bottom_out_27_[0]),
		.chany_in_28_(sb_2__0__0_chany_top_out_28_[0]),
		.chany_in_29_(sb_2__1__0_chany_bottom_out_29_[0]),
		.chany_in_30_(sb_2__0__0_chany_top_out_30_[0]),
		.chany_in_31_(sb_2__1__0_chany_bottom_out_31_[0]),
		.chany_in_32_(sb_2__0__0_chany_top_out_32_[0]),
		.chany_in_33_(sb_2__1__0_chany_bottom_out_33_[0]),
		.chany_in_34_(sb_2__0__0_chany_top_out_34_[0]),
		.chany_in_35_(sb_2__1__0_chany_bottom_out_35_[0]),
		.chany_in_36_(sb_2__0__0_chany_top_out_36_[0]),
		.chany_in_37_(sb_2__1__0_chany_bottom_out_37_[0]),
		.chany_in_38_(sb_2__0__0_chany_top_out_38_[0]),
		.chany_in_39_(sb_2__1__0_chany_bottom_out_39_[0]),
		.chany_in_40_(sb_2__0__0_chany_top_out_40_[0]),
		.chany_in_41_(sb_2__1__0_chany_bottom_out_41_[0]),
		.chany_in_42_(sb_2__0__0_chany_top_out_42_[0]),
		.chany_in_43_(sb_2__1__0_chany_bottom_out_43_[0]),
		.chany_in_44_(sb_2__0__0_chany_top_out_44_[0]),
		.chany_in_45_(sb_2__1__0_chany_bottom_out_45_[0]),
		.chany_in_46_(sb_2__0__0_chany_top_out_46_[0]),
		.chany_in_47_(sb_2__1__0_chany_bottom_out_47_[0]),
		.chany_in_48_(sb_2__0__0_chany_top_out_48_[0]),
		.chany_in_49_(sb_2__1__0_chany_bottom_out_49_[0]),
		.chany_in_50_(sb_2__0__0_chany_top_out_50_[0]),
		.chany_in_51_(sb_2__1__0_chany_bottom_out_51_[0]),
		.chany_in_52_(sb_2__0__0_chany_top_out_52_[0]),
		.chany_in_53_(sb_2__1__0_chany_bottom_out_53_[0]),
		.chany_in_54_(sb_2__0__0_chany_top_out_54_[0]),
		.chany_in_55_(sb_2__1__0_chany_bottom_out_55_[0]),
		.chany_in_56_(sb_2__0__0_chany_top_out_56_[0]),
		.chany_in_57_(sb_2__1__0_chany_bottom_out_57_[0]),
		.chany_in_58_(sb_2__0__0_chany_top_out_58_[0]),
		.chany_in_59_(sb_2__1__0_chany_bottom_out_59_[0]),
		.chany_in_60_(sb_2__0__0_chany_top_out_60_[0]),
		.chany_in_61_(sb_2__1__0_chany_bottom_out_61_[0]),
		.chany_in_62_(sb_2__0__0_chany_top_out_62_[0]),
		.chany_in_63_(sb_2__1__0_chany_bottom_out_63_[0]),
		.chany_in_64_(sb_2__0__0_chany_top_out_64_[0]),
		.chany_in_65_(sb_2__1__0_chany_bottom_out_65_[0]),
		.chany_in_66_(sb_2__0__0_chany_top_out_66_[0]),
		.chany_in_67_(sb_2__1__0_chany_bottom_out_67_[0]),
		.chany_in_68_(sb_2__0__0_chany_top_out_68_[0]),
		.chany_in_69_(sb_2__1__0_chany_bottom_out_69_[0]),
		.chany_in_70_(sb_2__0__0_chany_top_out_70_[0]),
		.chany_in_71_(sb_2__1__0_chany_bottom_out_71_[0]),
		.chany_in_72_(sb_2__0__0_chany_top_out_72_[0]),
		.chany_in_73_(sb_2__1__0_chany_bottom_out_73_[0]),
		.chany_in_74_(sb_2__0__0_chany_top_out_74_[0]),
		.chany_in_75_(sb_2__1__0_chany_bottom_out_75_[0]),
		.chany_in_76_(sb_2__0__0_chany_top_out_76_[0]),
		.chany_in_77_(sb_2__1__0_chany_bottom_out_77_[0]),
		.chany_in_78_(sb_2__0__0_chany_top_out_78_[0]),
		.chany_in_79_(sb_2__1__0_chany_bottom_out_79_[0]),
		.chany_in_80_(sb_2__0__0_chany_top_out_80_[0]),
		.chany_in_81_(sb_2__1__0_chany_bottom_out_81_[0]),
		.chany_in_82_(sb_2__0__0_chany_top_out_82_[0]),
		.chany_in_83_(sb_2__1__0_chany_bottom_out_83_[0]),
		.chany_in_84_(sb_2__0__0_chany_top_out_84_[0]),
		.chany_in_85_(sb_2__1__0_chany_bottom_out_85_[0]),
		.chany_in_86_(sb_2__0__0_chany_top_out_86_[0]),
		.chany_in_87_(sb_2__1__0_chany_bottom_out_87_[0]),
		.chany_in_88_(sb_2__0__0_chany_top_out_88_[0]),
		.chany_in_89_(sb_2__1__0_chany_bottom_out_89_[0]),
		.chany_in_90_(sb_2__0__0_chany_top_out_90_[0]),
		.chany_in_91_(sb_2__1__0_chany_bottom_out_91_[0]),
		.chany_in_92_(sb_2__0__0_chany_top_out_92_[0]),
		.chany_in_93_(sb_2__1__0_chany_bottom_out_93_[0]),
		.chany_in_94_(sb_2__0__0_chany_top_out_94_[0]),
		.chany_in_95_(sb_2__1__0_chany_bottom_out_95_[0]),
		.chany_in_96_(sb_2__0__0_chany_top_out_96_[0]),
		.chany_in_97_(sb_2__1__0_chany_bottom_out_97_[0]),
		.chany_in_98_(sb_2__0__0_chany_top_out_98_[0]),
		.chany_in_99_(sb_2__1__0_chany_bottom_out_99_[0]),
		.chany_in_100_(sb_2__0__0_chany_top_out_100_[0]),
		.chany_in_101_(sb_2__1__0_chany_bottom_out_101_[0]),
		.chany_in_102_(sb_2__0__0_chany_top_out_102_[0]),
		.chany_in_103_(sb_2__1__0_chany_bottom_out_103_[0]),
		.chany_in_104_(sb_2__0__0_chany_top_out_104_[0]),
		.chany_in_105_(sb_2__1__0_chany_bottom_out_105_[0]),
		.chany_in_106_(sb_2__0__0_chany_top_out_106_[0]),
		.chany_in_107_(sb_2__1__0_chany_bottom_out_107_[0]),
		.chany_in_108_(sb_2__0__0_chany_top_out_108_[0]),
		.chany_in_109_(sb_2__1__0_chany_bottom_out_109_[0]),
		.chany_in_110_(sb_2__0__0_chany_top_out_110_[0]),
		.chany_in_111_(sb_2__1__0_chany_bottom_out_111_[0]),
		.chany_in_112_(sb_2__0__0_chany_top_out_112_[0]),
		.chany_in_113_(sb_2__1__0_chany_bottom_out_113_[0]),
		.chany_in_114_(sb_2__0__0_chany_top_out_114_[0]),
		.chany_in_115_(sb_2__1__0_chany_bottom_out_115_[0]),
		.chany_in_116_(sb_2__0__0_chany_top_out_116_[0]),
		.chany_in_117_(sb_2__1__0_chany_bottom_out_117_[0]),
		.chany_in_118_(sb_2__0__0_chany_top_out_118_[0]),
		.chany_in_119_(sb_2__1__0_chany_bottom_out_119_[0]),
		.chany_in_120_(sb_2__0__0_chany_top_out_120_[0]),
		.chany_in_121_(sb_2__1__0_chany_bottom_out_121_[0]),
		.chany_in_122_(sb_2__0__0_chany_top_out_122_[0]),
		.chany_in_123_(sb_2__1__0_chany_bottom_out_123_[0]),
		.chany_in_124_(sb_2__0__0_chany_top_out_124_[0]),
		.chany_in_125_(sb_2__1__0_chany_bottom_out_125_[0]),
		.chany_in_126_(sb_2__0__0_chany_top_out_126_[0]),
		.chany_in_127_(sb_2__1__0_chany_bottom_out_127_[0]),
		.chany_in_128_(sb_2__0__0_chany_top_out_128_[0]),
		.chany_in_129_(sb_2__1__0_chany_bottom_out_129_[0]),
		.chany_in_130_(sb_2__0__0_chany_top_out_130_[0]),
		.chany_in_131_(sb_2__1__0_chany_bottom_out_131_[0]),
		.chany_in_132_(sb_2__0__0_chany_top_out_132_[0]),
		.chany_in_133_(sb_2__1__0_chany_bottom_out_133_[0]),
		.chany_in_134_(sb_2__0__0_chany_top_out_134_[0]),
		.chany_in_135_(sb_2__1__0_chany_bottom_out_135_[0]),
		.chany_in_136_(sb_2__0__0_chany_top_out_136_[0]),
		.chany_in_137_(sb_2__1__0_chany_bottom_out_137_[0]),
		.chany_in_138_(sb_2__0__0_chany_top_out_138_[0]),
		.chany_in_139_(sb_2__1__0_chany_bottom_out_139_[0]),
		.chany_in_140_(sb_2__0__0_chany_top_out_140_[0]),
		.chany_in_141_(sb_2__1__0_chany_bottom_out_141_[0]),
		.chany_in_142_(sb_2__0__0_chany_top_out_142_[0]),
		.chany_in_143_(sb_2__1__0_chany_bottom_out_143_[0]),
		.chany_in_144_(sb_2__0__0_chany_top_out_144_[0]),
		.chany_in_145_(sb_2__1__0_chany_bottom_out_145_[0]),
		.chany_in_146_(sb_2__0__0_chany_top_out_146_[0]),
		.chany_in_147_(sb_2__1__0_chany_bottom_out_147_[0]),
		.chany_in_148_(sb_2__0__0_chany_top_out_148_[0]),
		.chany_in_149_(sb_2__1__0_chany_bottom_out_149_[0]),
		.chany_in_150_(sb_2__0__0_chany_top_out_150_[0]),
		.chany_in_151_(sb_2__1__0_chany_bottom_out_151_[0]),
		.chany_in_152_(sb_2__0__0_chany_top_out_152_[0]),
		.chany_in_153_(sb_2__1__0_chany_bottom_out_153_[0]),
		.chany_in_154_(sb_2__0__0_chany_top_out_154_[0]),
		.chany_in_155_(sb_2__1__0_chany_bottom_out_155_[0]),
		.chany_in_156_(sb_2__0__0_chany_top_out_156_[0]),
		.chany_in_157_(sb_2__1__0_chany_bottom_out_157_[0]),
		.chany_in_158_(sb_2__0__0_chany_top_out_158_[0]),
		.chany_in_159_(sb_2__1__0_chany_bottom_out_159_[0]),
		.chany_in_160_(sb_2__0__0_chany_top_out_160_[0]),
		.chany_in_161_(sb_2__1__0_chany_bottom_out_161_[0]),
		.chany_in_162_(sb_2__0__0_chany_top_out_162_[0]),
		.chany_in_163_(sb_2__1__0_chany_bottom_out_163_[0]),
		.chany_in_164_(sb_2__0__0_chany_top_out_164_[0]),
		.chany_in_165_(sb_2__1__0_chany_bottom_out_165_[0]),
		.chany_in_166_(sb_2__0__0_chany_top_out_166_[0]),
		.chany_in_167_(sb_2__1__0_chany_bottom_out_167_[0]),
		.chany_in_168_(sb_2__0__0_chany_top_out_168_[0]),
		.chany_in_169_(sb_2__1__0_chany_bottom_out_169_[0]),
		.chany_in_170_(sb_2__0__0_chany_top_out_170_[0]),
		.chany_in_171_(sb_2__1__0_chany_bottom_out_171_[0]),
		.chany_in_172_(sb_2__0__0_chany_top_out_172_[0]),
		.chany_in_173_(sb_2__1__0_chany_bottom_out_173_[0]),
		.chany_in_174_(sb_2__0__0_chany_top_out_174_[0]),
		.chany_in_175_(sb_2__1__0_chany_bottom_out_175_[0]),
		.chany_in_176_(sb_2__0__0_chany_top_out_176_[0]),
		.chany_in_177_(sb_2__1__0_chany_bottom_out_177_[0]),
		.chany_in_178_(sb_2__0__0_chany_top_out_178_[0]),
		.chany_in_179_(sb_2__1__0_chany_bottom_out_179_[0]),
		.chany_in_180_(sb_2__0__0_chany_top_out_180_[0]),
		.chany_in_181_(sb_2__1__0_chany_bottom_out_181_[0]),
		.chany_in_182_(sb_2__0__0_chany_top_out_182_[0]),
		.chany_in_183_(sb_2__1__0_chany_bottom_out_183_[0]),
		.chany_in_184_(sb_2__0__0_chany_top_out_184_[0]),
		.chany_in_185_(sb_2__1__0_chany_bottom_out_185_[0]),
		.chany_in_186_(sb_2__0__0_chany_top_out_186_[0]),
		.chany_in_187_(sb_2__1__0_chany_bottom_out_187_[0]),
		.chany_in_188_(sb_2__0__0_chany_top_out_188_[0]),
		.chany_in_189_(sb_2__1__0_chany_bottom_out_189_[0]),
		.chany_in_190_(sb_2__0__0_chany_top_out_190_[0]),
		.chany_in_191_(sb_2__1__0_chany_bottom_out_191_[0]),
		.chany_in_192_(sb_2__0__0_chany_top_out_192_[0]),
		.chany_in_193_(sb_2__1__0_chany_bottom_out_193_[0]),
		.chany_in_194_(sb_2__0__0_chany_top_out_194_[0]),
		.chany_in_195_(sb_2__1__0_chany_bottom_out_195_[0]),
		.chany_in_196_(sb_2__0__0_chany_top_out_196_[0]),
		.chany_in_197_(sb_2__1__0_chany_bottom_out_197_[0]),
		.chany_in_198_(sb_2__0__0_chany_top_out_198_[0]),
		.chany_in_199_(sb_2__1__0_chany_bottom_out_199_[0]),
		.ccff_head(cbx_1__0__1_ccff_tail[0]),
		.chany_out_0_(cby_2__1__0_chany_out_0_[0]),
		.chany_out_1_(cby_2__1__0_chany_out_1_[0]),
		.chany_out_2_(cby_2__1__0_chany_out_2_[0]),
		.chany_out_3_(cby_2__1__0_chany_out_3_[0]),
		.chany_out_4_(cby_2__1__0_chany_out_4_[0]),
		.chany_out_5_(cby_2__1__0_chany_out_5_[0]),
		.chany_out_6_(cby_2__1__0_chany_out_6_[0]),
		.chany_out_7_(cby_2__1__0_chany_out_7_[0]),
		.chany_out_8_(cby_2__1__0_chany_out_8_[0]),
		.chany_out_9_(cby_2__1__0_chany_out_9_[0]),
		.chany_out_10_(cby_2__1__0_chany_out_10_[0]),
		.chany_out_11_(cby_2__1__0_chany_out_11_[0]),
		.chany_out_12_(cby_2__1__0_chany_out_12_[0]),
		.chany_out_13_(cby_2__1__0_chany_out_13_[0]),
		.chany_out_14_(cby_2__1__0_chany_out_14_[0]),
		.chany_out_15_(cby_2__1__0_chany_out_15_[0]),
		.chany_out_16_(cby_2__1__0_chany_out_16_[0]),
		.chany_out_17_(cby_2__1__0_chany_out_17_[0]),
		.chany_out_18_(cby_2__1__0_chany_out_18_[0]),
		.chany_out_19_(cby_2__1__0_chany_out_19_[0]),
		.chany_out_20_(cby_2__1__0_chany_out_20_[0]),
		.chany_out_21_(cby_2__1__0_chany_out_21_[0]),
		.chany_out_22_(cby_2__1__0_chany_out_22_[0]),
		.chany_out_23_(cby_2__1__0_chany_out_23_[0]),
		.chany_out_24_(cby_2__1__0_chany_out_24_[0]),
		.chany_out_25_(cby_2__1__0_chany_out_25_[0]),
		.chany_out_26_(cby_2__1__0_chany_out_26_[0]),
		.chany_out_27_(cby_2__1__0_chany_out_27_[0]),
		.chany_out_28_(cby_2__1__0_chany_out_28_[0]),
		.chany_out_29_(cby_2__1__0_chany_out_29_[0]),
		.chany_out_30_(cby_2__1__0_chany_out_30_[0]),
		.chany_out_31_(cby_2__1__0_chany_out_31_[0]),
		.chany_out_32_(cby_2__1__0_chany_out_32_[0]),
		.chany_out_33_(cby_2__1__0_chany_out_33_[0]),
		.chany_out_34_(cby_2__1__0_chany_out_34_[0]),
		.chany_out_35_(cby_2__1__0_chany_out_35_[0]),
		.chany_out_36_(cby_2__1__0_chany_out_36_[0]),
		.chany_out_37_(cby_2__1__0_chany_out_37_[0]),
		.chany_out_38_(cby_2__1__0_chany_out_38_[0]),
		.chany_out_39_(cby_2__1__0_chany_out_39_[0]),
		.chany_out_40_(cby_2__1__0_chany_out_40_[0]),
		.chany_out_41_(cby_2__1__0_chany_out_41_[0]),
		.chany_out_42_(cby_2__1__0_chany_out_42_[0]),
		.chany_out_43_(cby_2__1__0_chany_out_43_[0]),
		.chany_out_44_(cby_2__1__0_chany_out_44_[0]),
		.chany_out_45_(cby_2__1__0_chany_out_45_[0]),
		.chany_out_46_(cby_2__1__0_chany_out_46_[0]),
		.chany_out_47_(cby_2__1__0_chany_out_47_[0]),
		.chany_out_48_(cby_2__1__0_chany_out_48_[0]),
		.chany_out_49_(cby_2__1__0_chany_out_49_[0]),
		.chany_out_50_(cby_2__1__0_chany_out_50_[0]),
		.chany_out_51_(cby_2__1__0_chany_out_51_[0]),
		.chany_out_52_(cby_2__1__0_chany_out_52_[0]),
		.chany_out_53_(cby_2__1__0_chany_out_53_[0]),
		.chany_out_54_(cby_2__1__0_chany_out_54_[0]),
		.chany_out_55_(cby_2__1__0_chany_out_55_[0]),
		.chany_out_56_(cby_2__1__0_chany_out_56_[0]),
		.chany_out_57_(cby_2__1__0_chany_out_57_[0]),
		.chany_out_58_(cby_2__1__0_chany_out_58_[0]),
		.chany_out_59_(cby_2__1__0_chany_out_59_[0]),
		.chany_out_60_(cby_2__1__0_chany_out_60_[0]),
		.chany_out_61_(cby_2__1__0_chany_out_61_[0]),
		.chany_out_62_(cby_2__1__0_chany_out_62_[0]),
		.chany_out_63_(cby_2__1__0_chany_out_63_[0]),
		.chany_out_64_(cby_2__1__0_chany_out_64_[0]),
		.chany_out_65_(cby_2__1__0_chany_out_65_[0]),
		.chany_out_66_(cby_2__1__0_chany_out_66_[0]),
		.chany_out_67_(cby_2__1__0_chany_out_67_[0]),
		.chany_out_68_(cby_2__1__0_chany_out_68_[0]),
		.chany_out_69_(cby_2__1__0_chany_out_69_[0]),
		.chany_out_70_(cby_2__1__0_chany_out_70_[0]),
		.chany_out_71_(cby_2__1__0_chany_out_71_[0]),
		.chany_out_72_(cby_2__1__0_chany_out_72_[0]),
		.chany_out_73_(cby_2__1__0_chany_out_73_[0]),
		.chany_out_74_(cby_2__1__0_chany_out_74_[0]),
		.chany_out_75_(cby_2__1__0_chany_out_75_[0]),
		.chany_out_76_(cby_2__1__0_chany_out_76_[0]),
		.chany_out_77_(cby_2__1__0_chany_out_77_[0]),
		.chany_out_78_(cby_2__1__0_chany_out_78_[0]),
		.chany_out_79_(cby_2__1__0_chany_out_79_[0]),
		.chany_out_80_(cby_2__1__0_chany_out_80_[0]),
		.chany_out_81_(cby_2__1__0_chany_out_81_[0]),
		.chany_out_82_(cby_2__1__0_chany_out_82_[0]),
		.chany_out_83_(cby_2__1__0_chany_out_83_[0]),
		.chany_out_84_(cby_2__1__0_chany_out_84_[0]),
		.chany_out_85_(cby_2__1__0_chany_out_85_[0]),
		.chany_out_86_(cby_2__1__0_chany_out_86_[0]),
		.chany_out_87_(cby_2__1__0_chany_out_87_[0]),
		.chany_out_88_(cby_2__1__0_chany_out_88_[0]),
		.chany_out_89_(cby_2__1__0_chany_out_89_[0]),
		.chany_out_90_(cby_2__1__0_chany_out_90_[0]),
		.chany_out_91_(cby_2__1__0_chany_out_91_[0]),
		.chany_out_92_(cby_2__1__0_chany_out_92_[0]),
		.chany_out_93_(cby_2__1__0_chany_out_93_[0]),
		.chany_out_94_(cby_2__1__0_chany_out_94_[0]),
		.chany_out_95_(cby_2__1__0_chany_out_95_[0]),
		.chany_out_96_(cby_2__1__0_chany_out_96_[0]),
		.chany_out_97_(cby_2__1__0_chany_out_97_[0]),
		.chany_out_98_(cby_2__1__0_chany_out_98_[0]),
		.chany_out_99_(cby_2__1__0_chany_out_99_[0]),
		.chany_out_100_(cby_2__1__0_chany_out_100_[0]),
		.chany_out_101_(cby_2__1__0_chany_out_101_[0]),
		.chany_out_102_(cby_2__1__0_chany_out_102_[0]),
		.chany_out_103_(cby_2__1__0_chany_out_103_[0]),
		.chany_out_104_(cby_2__1__0_chany_out_104_[0]),
		.chany_out_105_(cby_2__1__0_chany_out_105_[0]),
		.chany_out_106_(cby_2__1__0_chany_out_106_[0]),
		.chany_out_107_(cby_2__1__0_chany_out_107_[0]),
		.chany_out_108_(cby_2__1__0_chany_out_108_[0]),
		.chany_out_109_(cby_2__1__0_chany_out_109_[0]),
		.chany_out_110_(cby_2__1__0_chany_out_110_[0]),
		.chany_out_111_(cby_2__1__0_chany_out_111_[0]),
		.chany_out_112_(cby_2__1__0_chany_out_112_[0]),
		.chany_out_113_(cby_2__1__0_chany_out_113_[0]),
		.chany_out_114_(cby_2__1__0_chany_out_114_[0]),
		.chany_out_115_(cby_2__1__0_chany_out_115_[0]),
		.chany_out_116_(cby_2__1__0_chany_out_116_[0]),
		.chany_out_117_(cby_2__1__0_chany_out_117_[0]),
		.chany_out_118_(cby_2__1__0_chany_out_118_[0]),
		.chany_out_119_(cby_2__1__0_chany_out_119_[0]),
		.chany_out_120_(cby_2__1__0_chany_out_120_[0]),
		.chany_out_121_(cby_2__1__0_chany_out_121_[0]),
		.chany_out_122_(cby_2__1__0_chany_out_122_[0]),
		.chany_out_123_(cby_2__1__0_chany_out_123_[0]),
		.chany_out_124_(cby_2__1__0_chany_out_124_[0]),
		.chany_out_125_(cby_2__1__0_chany_out_125_[0]),
		.chany_out_126_(cby_2__1__0_chany_out_126_[0]),
		.chany_out_127_(cby_2__1__0_chany_out_127_[0]),
		.chany_out_128_(cby_2__1__0_chany_out_128_[0]),
		.chany_out_129_(cby_2__1__0_chany_out_129_[0]),
		.chany_out_130_(cby_2__1__0_chany_out_130_[0]),
		.chany_out_131_(cby_2__1__0_chany_out_131_[0]),
		.chany_out_132_(cby_2__1__0_chany_out_132_[0]),
		.chany_out_133_(cby_2__1__0_chany_out_133_[0]),
		.chany_out_134_(cby_2__1__0_chany_out_134_[0]),
		.chany_out_135_(cby_2__1__0_chany_out_135_[0]),
		.chany_out_136_(cby_2__1__0_chany_out_136_[0]),
		.chany_out_137_(cby_2__1__0_chany_out_137_[0]),
		.chany_out_138_(cby_2__1__0_chany_out_138_[0]),
		.chany_out_139_(cby_2__1__0_chany_out_139_[0]),
		.chany_out_140_(cby_2__1__0_chany_out_140_[0]),
		.chany_out_141_(cby_2__1__0_chany_out_141_[0]),
		.chany_out_142_(cby_2__1__0_chany_out_142_[0]),
		.chany_out_143_(cby_2__1__0_chany_out_143_[0]),
		.chany_out_144_(cby_2__1__0_chany_out_144_[0]),
		.chany_out_145_(cby_2__1__0_chany_out_145_[0]),
		.chany_out_146_(cby_2__1__0_chany_out_146_[0]),
		.chany_out_147_(cby_2__1__0_chany_out_147_[0]),
		.chany_out_148_(cby_2__1__0_chany_out_148_[0]),
		.chany_out_149_(cby_2__1__0_chany_out_149_[0]),
		.chany_out_150_(cby_2__1__0_chany_out_150_[0]),
		.chany_out_151_(cby_2__1__0_chany_out_151_[0]),
		.chany_out_152_(cby_2__1__0_chany_out_152_[0]),
		.chany_out_153_(cby_2__1__0_chany_out_153_[0]),
		.chany_out_154_(cby_2__1__0_chany_out_154_[0]),
		.chany_out_155_(cby_2__1__0_chany_out_155_[0]),
		.chany_out_156_(cby_2__1__0_chany_out_156_[0]),
		.chany_out_157_(cby_2__1__0_chany_out_157_[0]),
		.chany_out_158_(cby_2__1__0_chany_out_158_[0]),
		.chany_out_159_(cby_2__1__0_chany_out_159_[0]),
		.chany_out_160_(cby_2__1__0_chany_out_160_[0]),
		.chany_out_161_(cby_2__1__0_chany_out_161_[0]),
		.chany_out_162_(cby_2__1__0_chany_out_162_[0]),
		.chany_out_163_(cby_2__1__0_chany_out_163_[0]),
		.chany_out_164_(cby_2__1__0_chany_out_164_[0]),
		.chany_out_165_(cby_2__1__0_chany_out_165_[0]),
		.chany_out_166_(cby_2__1__0_chany_out_166_[0]),
		.chany_out_167_(cby_2__1__0_chany_out_167_[0]),
		.chany_out_168_(cby_2__1__0_chany_out_168_[0]),
		.chany_out_169_(cby_2__1__0_chany_out_169_[0]),
		.chany_out_170_(cby_2__1__0_chany_out_170_[0]),
		.chany_out_171_(cby_2__1__0_chany_out_171_[0]),
		.chany_out_172_(cby_2__1__0_chany_out_172_[0]),
		.chany_out_173_(cby_2__1__0_chany_out_173_[0]),
		.chany_out_174_(cby_2__1__0_chany_out_174_[0]),
		.chany_out_175_(cby_2__1__0_chany_out_175_[0]),
		.chany_out_176_(cby_2__1__0_chany_out_176_[0]),
		.chany_out_177_(cby_2__1__0_chany_out_177_[0]),
		.chany_out_178_(cby_2__1__0_chany_out_178_[0]),
		.chany_out_179_(cby_2__1__0_chany_out_179_[0]),
		.chany_out_180_(cby_2__1__0_chany_out_180_[0]),
		.chany_out_181_(cby_2__1__0_chany_out_181_[0]),
		.chany_out_182_(cby_2__1__0_chany_out_182_[0]),
		.chany_out_183_(cby_2__1__0_chany_out_183_[0]),
		.chany_out_184_(cby_2__1__0_chany_out_184_[0]),
		.chany_out_185_(cby_2__1__0_chany_out_185_[0]),
		.chany_out_186_(cby_2__1__0_chany_out_186_[0]),
		.chany_out_187_(cby_2__1__0_chany_out_187_[0]),
		.chany_out_188_(cby_2__1__0_chany_out_188_[0]),
		.chany_out_189_(cby_2__1__0_chany_out_189_[0]),
		.chany_out_190_(cby_2__1__0_chany_out_190_[0]),
		.chany_out_191_(cby_2__1__0_chany_out_191_[0]),
		.chany_out_192_(cby_2__1__0_chany_out_192_[0]),
		.chany_out_193_(cby_2__1__0_chany_out_193_[0]),
		.chany_out_194_(cby_2__1__0_chany_out_194_[0]),
		.chany_out_195_(cby_2__1__0_chany_out_195_[0]),
		.chany_out_196_(cby_2__1__0_chany_out_196_[0]),
		.chany_out_197_(cby_2__1__0_chany_out_197_[0]),
		.chany_out_198_(cby_2__1__0_chany_out_198_[0]),
		.chany_out_199_(cby_2__1__0_chany_out_199_[0]),
		.right_grid_pin_0_(cby_2__1__0_right_grid_pin_0_[0]),
		.left_grid_pin_0_(cby_2__1__0_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_2__1__0_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_2__1__0_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_2__1__0_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_2__1__0_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_2__1__0_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_2__1__0_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_2__1__0_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_2__1__0_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_2__1__0_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_2__1__0_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_2__1__0_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_2__1__0_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_2__1__0_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_2__1__0_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_2__1__0_left_grid_pin_15_[0]),
		.left_grid_pin_16_(cby_2__1__0_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_2__1__0_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_2__1__0_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_2__1__0_left_grid_pin_19_[0]),
		.ccff_tail(cby_2__1__0_ccff_tail[0]));

	cby_2__1_ cby_2__2_ (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.chany_in_0_(sb_2__1__0_chany_top_out_0_[0]),
		.chany_in_1_(sb_2__2__0_chany_bottom_out_1_[0]),
		.chany_in_2_(sb_2__1__0_chany_top_out_2_[0]),
		.chany_in_3_(sb_2__2__0_chany_bottom_out_3_[0]),
		.chany_in_4_(sb_2__1__0_chany_top_out_4_[0]),
		.chany_in_5_(sb_2__2__0_chany_bottom_out_5_[0]),
		.chany_in_6_(sb_2__1__0_chany_top_out_6_[0]),
		.chany_in_7_(sb_2__2__0_chany_bottom_out_7_[0]),
		.chany_in_8_(sb_2__1__0_chany_top_out_8_[0]),
		.chany_in_9_(sb_2__2__0_chany_bottom_out_9_[0]),
		.chany_in_10_(sb_2__1__0_chany_top_out_10_[0]),
		.chany_in_11_(sb_2__2__0_chany_bottom_out_11_[0]),
		.chany_in_12_(sb_2__1__0_chany_top_out_12_[0]),
		.chany_in_13_(sb_2__2__0_chany_bottom_out_13_[0]),
		.chany_in_14_(sb_2__1__0_chany_top_out_14_[0]),
		.chany_in_15_(sb_2__2__0_chany_bottom_out_15_[0]),
		.chany_in_16_(sb_2__1__0_chany_top_out_16_[0]),
		.chany_in_17_(sb_2__2__0_chany_bottom_out_17_[0]),
		.chany_in_18_(sb_2__1__0_chany_top_out_18_[0]),
		.chany_in_19_(sb_2__2__0_chany_bottom_out_19_[0]),
		.chany_in_20_(sb_2__1__0_chany_top_out_20_[0]),
		.chany_in_21_(sb_2__2__0_chany_bottom_out_21_[0]),
		.chany_in_22_(sb_2__1__0_chany_top_out_22_[0]),
		.chany_in_23_(sb_2__2__0_chany_bottom_out_23_[0]),
		.chany_in_24_(sb_2__1__0_chany_top_out_24_[0]),
		.chany_in_25_(sb_2__2__0_chany_bottom_out_25_[0]),
		.chany_in_26_(sb_2__1__0_chany_top_out_26_[0]),
		.chany_in_27_(sb_2__2__0_chany_bottom_out_27_[0]),
		.chany_in_28_(sb_2__1__0_chany_top_out_28_[0]),
		.chany_in_29_(sb_2__2__0_chany_bottom_out_29_[0]),
		.chany_in_30_(sb_2__1__0_chany_top_out_30_[0]),
		.chany_in_31_(sb_2__2__0_chany_bottom_out_31_[0]),
		.chany_in_32_(sb_2__1__0_chany_top_out_32_[0]),
		.chany_in_33_(sb_2__2__0_chany_bottom_out_33_[0]),
		.chany_in_34_(sb_2__1__0_chany_top_out_34_[0]),
		.chany_in_35_(sb_2__2__0_chany_bottom_out_35_[0]),
		.chany_in_36_(sb_2__1__0_chany_top_out_36_[0]),
		.chany_in_37_(sb_2__2__0_chany_bottom_out_37_[0]),
		.chany_in_38_(sb_2__1__0_chany_top_out_38_[0]),
		.chany_in_39_(sb_2__2__0_chany_bottom_out_39_[0]),
		.chany_in_40_(sb_2__1__0_chany_top_out_40_[0]),
		.chany_in_41_(sb_2__2__0_chany_bottom_out_41_[0]),
		.chany_in_42_(sb_2__1__0_chany_top_out_42_[0]),
		.chany_in_43_(sb_2__2__0_chany_bottom_out_43_[0]),
		.chany_in_44_(sb_2__1__0_chany_top_out_44_[0]),
		.chany_in_45_(sb_2__2__0_chany_bottom_out_45_[0]),
		.chany_in_46_(sb_2__1__0_chany_top_out_46_[0]),
		.chany_in_47_(sb_2__2__0_chany_bottom_out_47_[0]),
		.chany_in_48_(sb_2__1__0_chany_top_out_48_[0]),
		.chany_in_49_(sb_2__2__0_chany_bottom_out_49_[0]),
		.chany_in_50_(sb_2__1__0_chany_top_out_50_[0]),
		.chany_in_51_(sb_2__2__0_chany_bottom_out_51_[0]),
		.chany_in_52_(sb_2__1__0_chany_top_out_52_[0]),
		.chany_in_53_(sb_2__2__0_chany_bottom_out_53_[0]),
		.chany_in_54_(sb_2__1__0_chany_top_out_54_[0]),
		.chany_in_55_(sb_2__2__0_chany_bottom_out_55_[0]),
		.chany_in_56_(sb_2__1__0_chany_top_out_56_[0]),
		.chany_in_57_(sb_2__2__0_chany_bottom_out_57_[0]),
		.chany_in_58_(sb_2__1__0_chany_top_out_58_[0]),
		.chany_in_59_(sb_2__2__0_chany_bottom_out_59_[0]),
		.chany_in_60_(sb_2__1__0_chany_top_out_60_[0]),
		.chany_in_61_(sb_2__2__0_chany_bottom_out_61_[0]),
		.chany_in_62_(sb_2__1__0_chany_top_out_62_[0]),
		.chany_in_63_(sb_2__2__0_chany_bottom_out_63_[0]),
		.chany_in_64_(sb_2__1__0_chany_top_out_64_[0]),
		.chany_in_65_(sb_2__2__0_chany_bottom_out_65_[0]),
		.chany_in_66_(sb_2__1__0_chany_top_out_66_[0]),
		.chany_in_67_(sb_2__2__0_chany_bottom_out_67_[0]),
		.chany_in_68_(sb_2__1__0_chany_top_out_68_[0]),
		.chany_in_69_(sb_2__2__0_chany_bottom_out_69_[0]),
		.chany_in_70_(sb_2__1__0_chany_top_out_70_[0]),
		.chany_in_71_(sb_2__2__0_chany_bottom_out_71_[0]),
		.chany_in_72_(sb_2__1__0_chany_top_out_72_[0]),
		.chany_in_73_(sb_2__2__0_chany_bottom_out_73_[0]),
		.chany_in_74_(sb_2__1__0_chany_top_out_74_[0]),
		.chany_in_75_(sb_2__2__0_chany_bottom_out_75_[0]),
		.chany_in_76_(sb_2__1__0_chany_top_out_76_[0]),
		.chany_in_77_(sb_2__2__0_chany_bottom_out_77_[0]),
		.chany_in_78_(sb_2__1__0_chany_top_out_78_[0]),
		.chany_in_79_(sb_2__2__0_chany_bottom_out_79_[0]),
		.chany_in_80_(sb_2__1__0_chany_top_out_80_[0]),
		.chany_in_81_(sb_2__2__0_chany_bottom_out_81_[0]),
		.chany_in_82_(sb_2__1__0_chany_top_out_82_[0]),
		.chany_in_83_(sb_2__2__0_chany_bottom_out_83_[0]),
		.chany_in_84_(sb_2__1__0_chany_top_out_84_[0]),
		.chany_in_85_(sb_2__2__0_chany_bottom_out_85_[0]),
		.chany_in_86_(sb_2__1__0_chany_top_out_86_[0]),
		.chany_in_87_(sb_2__2__0_chany_bottom_out_87_[0]),
		.chany_in_88_(sb_2__1__0_chany_top_out_88_[0]),
		.chany_in_89_(sb_2__2__0_chany_bottom_out_89_[0]),
		.chany_in_90_(sb_2__1__0_chany_top_out_90_[0]),
		.chany_in_91_(sb_2__2__0_chany_bottom_out_91_[0]),
		.chany_in_92_(sb_2__1__0_chany_top_out_92_[0]),
		.chany_in_93_(sb_2__2__0_chany_bottom_out_93_[0]),
		.chany_in_94_(sb_2__1__0_chany_top_out_94_[0]),
		.chany_in_95_(sb_2__2__0_chany_bottom_out_95_[0]),
		.chany_in_96_(sb_2__1__0_chany_top_out_96_[0]),
		.chany_in_97_(sb_2__2__0_chany_bottom_out_97_[0]),
		.chany_in_98_(sb_2__1__0_chany_top_out_98_[0]),
		.chany_in_99_(sb_2__2__0_chany_bottom_out_99_[0]),
		.chany_in_100_(sb_2__1__0_chany_top_out_100_[0]),
		.chany_in_101_(sb_2__2__0_chany_bottom_out_101_[0]),
		.chany_in_102_(sb_2__1__0_chany_top_out_102_[0]),
		.chany_in_103_(sb_2__2__0_chany_bottom_out_103_[0]),
		.chany_in_104_(sb_2__1__0_chany_top_out_104_[0]),
		.chany_in_105_(sb_2__2__0_chany_bottom_out_105_[0]),
		.chany_in_106_(sb_2__1__0_chany_top_out_106_[0]),
		.chany_in_107_(sb_2__2__0_chany_bottom_out_107_[0]),
		.chany_in_108_(sb_2__1__0_chany_top_out_108_[0]),
		.chany_in_109_(sb_2__2__0_chany_bottom_out_109_[0]),
		.chany_in_110_(sb_2__1__0_chany_top_out_110_[0]),
		.chany_in_111_(sb_2__2__0_chany_bottom_out_111_[0]),
		.chany_in_112_(sb_2__1__0_chany_top_out_112_[0]),
		.chany_in_113_(sb_2__2__0_chany_bottom_out_113_[0]),
		.chany_in_114_(sb_2__1__0_chany_top_out_114_[0]),
		.chany_in_115_(sb_2__2__0_chany_bottom_out_115_[0]),
		.chany_in_116_(sb_2__1__0_chany_top_out_116_[0]),
		.chany_in_117_(sb_2__2__0_chany_bottom_out_117_[0]),
		.chany_in_118_(sb_2__1__0_chany_top_out_118_[0]),
		.chany_in_119_(sb_2__2__0_chany_bottom_out_119_[0]),
		.chany_in_120_(sb_2__1__0_chany_top_out_120_[0]),
		.chany_in_121_(sb_2__2__0_chany_bottom_out_121_[0]),
		.chany_in_122_(sb_2__1__0_chany_top_out_122_[0]),
		.chany_in_123_(sb_2__2__0_chany_bottom_out_123_[0]),
		.chany_in_124_(sb_2__1__0_chany_top_out_124_[0]),
		.chany_in_125_(sb_2__2__0_chany_bottom_out_125_[0]),
		.chany_in_126_(sb_2__1__0_chany_top_out_126_[0]),
		.chany_in_127_(sb_2__2__0_chany_bottom_out_127_[0]),
		.chany_in_128_(sb_2__1__0_chany_top_out_128_[0]),
		.chany_in_129_(sb_2__2__0_chany_bottom_out_129_[0]),
		.chany_in_130_(sb_2__1__0_chany_top_out_130_[0]),
		.chany_in_131_(sb_2__2__0_chany_bottom_out_131_[0]),
		.chany_in_132_(sb_2__1__0_chany_top_out_132_[0]),
		.chany_in_133_(sb_2__2__0_chany_bottom_out_133_[0]),
		.chany_in_134_(sb_2__1__0_chany_top_out_134_[0]),
		.chany_in_135_(sb_2__2__0_chany_bottom_out_135_[0]),
		.chany_in_136_(sb_2__1__0_chany_top_out_136_[0]),
		.chany_in_137_(sb_2__2__0_chany_bottom_out_137_[0]),
		.chany_in_138_(sb_2__1__0_chany_top_out_138_[0]),
		.chany_in_139_(sb_2__2__0_chany_bottom_out_139_[0]),
		.chany_in_140_(sb_2__1__0_chany_top_out_140_[0]),
		.chany_in_141_(sb_2__2__0_chany_bottom_out_141_[0]),
		.chany_in_142_(sb_2__1__0_chany_top_out_142_[0]),
		.chany_in_143_(sb_2__2__0_chany_bottom_out_143_[0]),
		.chany_in_144_(sb_2__1__0_chany_top_out_144_[0]),
		.chany_in_145_(sb_2__2__0_chany_bottom_out_145_[0]),
		.chany_in_146_(sb_2__1__0_chany_top_out_146_[0]),
		.chany_in_147_(sb_2__2__0_chany_bottom_out_147_[0]),
		.chany_in_148_(sb_2__1__0_chany_top_out_148_[0]),
		.chany_in_149_(sb_2__2__0_chany_bottom_out_149_[0]),
		.chany_in_150_(sb_2__1__0_chany_top_out_150_[0]),
		.chany_in_151_(sb_2__2__0_chany_bottom_out_151_[0]),
		.chany_in_152_(sb_2__1__0_chany_top_out_152_[0]),
		.chany_in_153_(sb_2__2__0_chany_bottom_out_153_[0]),
		.chany_in_154_(sb_2__1__0_chany_top_out_154_[0]),
		.chany_in_155_(sb_2__2__0_chany_bottom_out_155_[0]),
		.chany_in_156_(sb_2__1__0_chany_top_out_156_[0]),
		.chany_in_157_(sb_2__2__0_chany_bottom_out_157_[0]),
		.chany_in_158_(sb_2__1__0_chany_top_out_158_[0]),
		.chany_in_159_(sb_2__2__0_chany_bottom_out_159_[0]),
		.chany_in_160_(sb_2__1__0_chany_top_out_160_[0]),
		.chany_in_161_(sb_2__2__0_chany_bottom_out_161_[0]),
		.chany_in_162_(sb_2__1__0_chany_top_out_162_[0]),
		.chany_in_163_(sb_2__2__0_chany_bottom_out_163_[0]),
		.chany_in_164_(sb_2__1__0_chany_top_out_164_[0]),
		.chany_in_165_(sb_2__2__0_chany_bottom_out_165_[0]),
		.chany_in_166_(sb_2__1__0_chany_top_out_166_[0]),
		.chany_in_167_(sb_2__2__0_chany_bottom_out_167_[0]),
		.chany_in_168_(sb_2__1__0_chany_top_out_168_[0]),
		.chany_in_169_(sb_2__2__0_chany_bottom_out_169_[0]),
		.chany_in_170_(sb_2__1__0_chany_top_out_170_[0]),
		.chany_in_171_(sb_2__2__0_chany_bottom_out_171_[0]),
		.chany_in_172_(sb_2__1__0_chany_top_out_172_[0]),
		.chany_in_173_(sb_2__2__0_chany_bottom_out_173_[0]),
		.chany_in_174_(sb_2__1__0_chany_top_out_174_[0]),
		.chany_in_175_(sb_2__2__0_chany_bottom_out_175_[0]),
		.chany_in_176_(sb_2__1__0_chany_top_out_176_[0]),
		.chany_in_177_(sb_2__2__0_chany_bottom_out_177_[0]),
		.chany_in_178_(sb_2__1__0_chany_top_out_178_[0]),
		.chany_in_179_(sb_2__2__0_chany_bottom_out_179_[0]),
		.chany_in_180_(sb_2__1__0_chany_top_out_180_[0]),
		.chany_in_181_(sb_2__2__0_chany_bottom_out_181_[0]),
		.chany_in_182_(sb_2__1__0_chany_top_out_182_[0]),
		.chany_in_183_(sb_2__2__0_chany_bottom_out_183_[0]),
		.chany_in_184_(sb_2__1__0_chany_top_out_184_[0]),
		.chany_in_185_(sb_2__2__0_chany_bottom_out_185_[0]),
		.chany_in_186_(sb_2__1__0_chany_top_out_186_[0]),
		.chany_in_187_(sb_2__2__0_chany_bottom_out_187_[0]),
		.chany_in_188_(sb_2__1__0_chany_top_out_188_[0]),
		.chany_in_189_(sb_2__2__0_chany_bottom_out_189_[0]),
		.chany_in_190_(sb_2__1__0_chany_top_out_190_[0]),
		.chany_in_191_(sb_2__2__0_chany_bottom_out_191_[0]),
		.chany_in_192_(sb_2__1__0_chany_top_out_192_[0]),
		.chany_in_193_(sb_2__2__0_chany_bottom_out_193_[0]),
		.chany_in_194_(sb_2__1__0_chany_top_out_194_[0]),
		.chany_in_195_(sb_2__2__0_chany_bottom_out_195_[0]),
		.chany_in_196_(sb_2__1__0_chany_top_out_196_[0]),
		.chany_in_197_(sb_2__2__0_chany_bottom_out_197_[0]),
		.chany_in_198_(sb_2__1__0_chany_top_out_198_[0]),
		.chany_in_199_(sb_2__2__0_chany_bottom_out_199_[0]),
		.ccff_head(cbx_1__1__1_ccff_tail[0]),
		.chany_out_0_(cby_2__1__1_chany_out_0_[0]),
		.chany_out_1_(cby_2__1__1_chany_out_1_[0]),
		.chany_out_2_(cby_2__1__1_chany_out_2_[0]),
		.chany_out_3_(cby_2__1__1_chany_out_3_[0]),
		.chany_out_4_(cby_2__1__1_chany_out_4_[0]),
		.chany_out_5_(cby_2__1__1_chany_out_5_[0]),
		.chany_out_6_(cby_2__1__1_chany_out_6_[0]),
		.chany_out_7_(cby_2__1__1_chany_out_7_[0]),
		.chany_out_8_(cby_2__1__1_chany_out_8_[0]),
		.chany_out_9_(cby_2__1__1_chany_out_9_[0]),
		.chany_out_10_(cby_2__1__1_chany_out_10_[0]),
		.chany_out_11_(cby_2__1__1_chany_out_11_[0]),
		.chany_out_12_(cby_2__1__1_chany_out_12_[0]),
		.chany_out_13_(cby_2__1__1_chany_out_13_[0]),
		.chany_out_14_(cby_2__1__1_chany_out_14_[0]),
		.chany_out_15_(cby_2__1__1_chany_out_15_[0]),
		.chany_out_16_(cby_2__1__1_chany_out_16_[0]),
		.chany_out_17_(cby_2__1__1_chany_out_17_[0]),
		.chany_out_18_(cby_2__1__1_chany_out_18_[0]),
		.chany_out_19_(cby_2__1__1_chany_out_19_[0]),
		.chany_out_20_(cby_2__1__1_chany_out_20_[0]),
		.chany_out_21_(cby_2__1__1_chany_out_21_[0]),
		.chany_out_22_(cby_2__1__1_chany_out_22_[0]),
		.chany_out_23_(cby_2__1__1_chany_out_23_[0]),
		.chany_out_24_(cby_2__1__1_chany_out_24_[0]),
		.chany_out_25_(cby_2__1__1_chany_out_25_[0]),
		.chany_out_26_(cby_2__1__1_chany_out_26_[0]),
		.chany_out_27_(cby_2__1__1_chany_out_27_[0]),
		.chany_out_28_(cby_2__1__1_chany_out_28_[0]),
		.chany_out_29_(cby_2__1__1_chany_out_29_[0]),
		.chany_out_30_(cby_2__1__1_chany_out_30_[0]),
		.chany_out_31_(cby_2__1__1_chany_out_31_[0]),
		.chany_out_32_(cby_2__1__1_chany_out_32_[0]),
		.chany_out_33_(cby_2__1__1_chany_out_33_[0]),
		.chany_out_34_(cby_2__1__1_chany_out_34_[0]),
		.chany_out_35_(cby_2__1__1_chany_out_35_[0]),
		.chany_out_36_(cby_2__1__1_chany_out_36_[0]),
		.chany_out_37_(cby_2__1__1_chany_out_37_[0]),
		.chany_out_38_(cby_2__1__1_chany_out_38_[0]),
		.chany_out_39_(cby_2__1__1_chany_out_39_[0]),
		.chany_out_40_(cby_2__1__1_chany_out_40_[0]),
		.chany_out_41_(cby_2__1__1_chany_out_41_[0]),
		.chany_out_42_(cby_2__1__1_chany_out_42_[0]),
		.chany_out_43_(cby_2__1__1_chany_out_43_[0]),
		.chany_out_44_(cby_2__1__1_chany_out_44_[0]),
		.chany_out_45_(cby_2__1__1_chany_out_45_[0]),
		.chany_out_46_(cby_2__1__1_chany_out_46_[0]),
		.chany_out_47_(cby_2__1__1_chany_out_47_[0]),
		.chany_out_48_(cby_2__1__1_chany_out_48_[0]),
		.chany_out_49_(cby_2__1__1_chany_out_49_[0]),
		.chany_out_50_(cby_2__1__1_chany_out_50_[0]),
		.chany_out_51_(cby_2__1__1_chany_out_51_[0]),
		.chany_out_52_(cby_2__1__1_chany_out_52_[0]),
		.chany_out_53_(cby_2__1__1_chany_out_53_[0]),
		.chany_out_54_(cby_2__1__1_chany_out_54_[0]),
		.chany_out_55_(cby_2__1__1_chany_out_55_[0]),
		.chany_out_56_(cby_2__1__1_chany_out_56_[0]),
		.chany_out_57_(cby_2__1__1_chany_out_57_[0]),
		.chany_out_58_(cby_2__1__1_chany_out_58_[0]),
		.chany_out_59_(cby_2__1__1_chany_out_59_[0]),
		.chany_out_60_(cby_2__1__1_chany_out_60_[0]),
		.chany_out_61_(cby_2__1__1_chany_out_61_[0]),
		.chany_out_62_(cby_2__1__1_chany_out_62_[0]),
		.chany_out_63_(cby_2__1__1_chany_out_63_[0]),
		.chany_out_64_(cby_2__1__1_chany_out_64_[0]),
		.chany_out_65_(cby_2__1__1_chany_out_65_[0]),
		.chany_out_66_(cby_2__1__1_chany_out_66_[0]),
		.chany_out_67_(cby_2__1__1_chany_out_67_[0]),
		.chany_out_68_(cby_2__1__1_chany_out_68_[0]),
		.chany_out_69_(cby_2__1__1_chany_out_69_[0]),
		.chany_out_70_(cby_2__1__1_chany_out_70_[0]),
		.chany_out_71_(cby_2__1__1_chany_out_71_[0]),
		.chany_out_72_(cby_2__1__1_chany_out_72_[0]),
		.chany_out_73_(cby_2__1__1_chany_out_73_[0]),
		.chany_out_74_(cby_2__1__1_chany_out_74_[0]),
		.chany_out_75_(cby_2__1__1_chany_out_75_[0]),
		.chany_out_76_(cby_2__1__1_chany_out_76_[0]),
		.chany_out_77_(cby_2__1__1_chany_out_77_[0]),
		.chany_out_78_(cby_2__1__1_chany_out_78_[0]),
		.chany_out_79_(cby_2__1__1_chany_out_79_[0]),
		.chany_out_80_(cby_2__1__1_chany_out_80_[0]),
		.chany_out_81_(cby_2__1__1_chany_out_81_[0]),
		.chany_out_82_(cby_2__1__1_chany_out_82_[0]),
		.chany_out_83_(cby_2__1__1_chany_out_83_[0]),
		.chany_out_84_(cby_2__1__1_chany_out_84_[0]),
		.chany_out_85_(cby_2__1__1_chany_out_85_[0]),
		.chany_out_86_(cby_2__1__1_chany_out_86_[0]),
		.chany_out_87_(cby_2__1__1_chany_out_87_[0]),
		.chany_out_88_(cby_2__1__1_chany_out_88_[0]),
		.chany_out_89_(cby_2__1__1_chany_out_89_[0]),
		.chany_out_90_(cby_2__1__1_chany_out_90_[0]),
		.chany_out_91_(cby_2__1__1_chany_out_91_[0]),
		.chany_out_92_(cby_2__1__1_chany_out_92_[0]),
		.chany_out_93_(cby_2__1__1_chany_out_93_[0]),
		.chany_out_94_(cby_2__1__1_chany_out_94_[0]),
		.chany_out_95_(cby_2__1__1_chany_out_95_[0]),
		.chany_out_96_(cby_2__1__1_chany_out_96_[0]),
		.chany_out_97_(cby_2__1__1_chany_out_97_[0]),
		.chany_out_98_(cby_2__1__1_chany_out_98_[0]),
		.chany_out_99_(cby_2__1__1_chany_out_99_[0]),
		.chany_out_100_(cby_2__1__1_chany_out_100_[0]),
		.chany_out_101_(cby_2__1__1_chany_out_101_[0]),
		.chany_out_102_(cby_2__1__1_chany_out_102_[0]),
		.chany_out_103_(cby_2__1__1_chany_out_103_[0]),
		.chany_out_104_(cby_2__1__1_chany_out_104_[0]),
		.chany_out_105_(cby_2__1__1_chany_out_105_[0]),
		.chany_out_106_(cby_2__1__1_chany_out_106_[0]),
		.chany_out_107_(cby_2__1__1_chany_out_107_[0]),
		.chany_out_108_(cby_2__1__1_chany_out_108_[0]),
		.chany_out_109_(cby_2__1__1_chany_out_109_[0]),
		.chany_out_110_(cby_2__1__1_chany_out_110_[0]),
		.chany_out_111_(cby_2__1__1_chany_out_111_[0]),
		.chany_out_112_(cby_2__1__1_chany_out_112_[0]),
		.chany_out_113_(cby_2__1__1_chany_out_113_[0]),
		.chany_out_114_(cby_2__1__1_chany_out_114_[0]),
		.chany_out_115_(cby_2__1__1_chany_out_115_[0]),
		.chany_out_116_(cby_2__1__1_chany_out_116_[0]),
		.chany_out_117_(cby_2__1__1_chany_out_117_[0]),
		.chany_out_118_(cby_2__1__1_chany_out_118_[0]),
		.chany_out_119_(cby_2__1__1_chany_out_119_[0]),
		.chany_out_120_(cby_2__1__1_chany_out_120_[0]),
		.chany_out_121_(cby_2__1__1_chany_out_121_[0]),
		.chany_out_122_(cby_2__1__1_chany_out_122_[0]),
		.chany_out_123_(cby_2__1__1_chany_out_123_[0]),
		.chany_out_124_(cby_2__1__1_chany_out_124_[0]),
		.chany_out_125_(cby_2__1__1_chany_out_125_[0]),
		.chany_out_126_(cby_2__1__1_chany_out_126_[0]),
		.chany_out_127_(cby_2__1__1_chany_out_127_[0]),
		.chany_out_128_(cby_2__1__1_chany_out_128_[0]),
		.chany_out_129_(cby_2__1__1_chany_out_129_[0]),
		.chany_out_130_(cby_2__1__1_chany_out_130_[0]),
		.chany_out_131_(cby_2__1__1_chany_out_131_[0]),
		.chany_out_132_(cby_2__1__1_chany_out_132_[0]),
		.chany_out_133_(cby_2__1__1_chany_out_133_[0]),
		.chany_out_134_(cby_2__1__1_chany_out_134_[0]),
		.chany_out_135_(cby_2__1__1_chany_out_135_[0]),
		.chany_out_136_(cby_2__1__1_chany_out_136_[0]),
		.chany_out_137_(cby_2__1__1_chany_out_137_[0]),
		.chany_out_138_(cby_2__1__1_chany_out_138_[0]),
		.chany_out_139_(cby_2__1__1_chany_out_139_[0]),
		.chany_out_140_(cby_2__1__1_chany_out_140_[0]),
		.chany_out_141_(cby_2__1__1_chany_out_141_[0]),
		.chany_out_142_(cby_2__1__1_chany_out_142_[0]),
		.chany_out_143_(cby_2__1__1_chany_out_143_[0]),
		.chany_out_144_(cby_2__1__1_chany_out_144_[0]),
		.chany_out_145_(cby_2__1__1_chany_out_145_[0]),
		.chany_out_146_(cby_2__1__1_chany_out_146_[0]),
		.chany_out_147_(cby_2__1__1_chany_out_147_[0]),
		.chany_out_148_(cby_2__1__1_chany_out_148_[0]),
		.chany_out_149_(cby_2__1__1_chany_out_149_[0]),
		.chany_out_150_(cby_2__1__1_chany_out_150_[0]),
		.chany_out_151_(cby_2__1__1_chany_out_151_[0]),
		.chany_out_152_(cby_2__1__1_chany_out_152_[0]),
		.chany_out_153_(cby_2__1__1_chany_out_153_[0]),
		.chany_out_154_(cby_2__1__1_chany_out_154_[0]),
		.chany_out_155_(cby_2__1__1_chany_out_155_[0]),
		.chany_out_156_(cby_2__1__1_chany_out_156_[0]),
		.chany_out_157_(cby_2__1__1_chany_out_157_[0]),
		.chany_out_158_(cby_2__1__1_chany_out_158_[0]),
		.chany_out_159_(cby_2__1__1_chany_out_159_[0]),
		.chany_out_160_(cby_2__1__1_chany_out_160_[0]),
		.chany_out_161_(cby_2__1__1_chany_out_161_[0]),
		.chany_out_162_(cby_2__1__1_chany_out_162_[0]),
		.chany_out_163_(cby_2__1__1_chany_out_163_[0]),
		.chany_out_164_(cby_2__1__1_chany_out_164_[0]),
		.chany_out_165_(cby_2__1__1_chany_out_165_[0]),
		.chany_out_166_(cby_2__1__1_chany_out_166_[0]),
		.chany_out_167_(cby_2__1__1_chany_out_167_[0]),
		.chany_out_168_(cby_2__1__1_chany_out_168_[0]),
		.chany_out_169_(cby_2__1__1_chany_out_169_[0]),
		.chany_out_170_(cby_2__1__1_chany_out_170_[0]),
		.chany_out_171_(cby_2__1__1_chany_out_171_[0]),
		.chany_out_172_(cby_2__1__1_chany_out_172_[0]),
		.chany_out_173_(cby_2__1__1_chany_out_173_[0]),
		.chany_out_174_(cby_2__1__1_chany_out_174_[0]),
		.chany_out_175_(cby_2__1__1_chany_out_175_[0]),
		.chany_out_176_(cby_2__1__1_chany_out_176_[0]),
		.chany_out_177_(cby_2__1__1_chany_out_177_[0]),
		.chany_out_178_(cby_2__1__1_chany_out_178_[0]),
		.chany_out_179_(cby_2__1__1_chany_out_179_[0]),
		.chany_out_180_(cby_2__1__1_chany_out_180_[0]),
		.chany_out_181_(cby_2__1__1_chany_out_181_[0]),
		.chany_out_182_(cby_2__1__1_chany_out_182_[0]),
		.chany_out_183_(cby_2__1__1_chany_out_183_[0]),
		.chany_out_184_(cby_2__1__1_chany_out_184_[0]),
		.chany_out_185_(cby_2__1__1_chany_out_185_[0]),
		.chany_out_186_(cby_2__1__1_chany_out_186_[0]),
		.chany_out_187_(cby_2__1__1_chany_out_187_[0]),
		.chany_out_188_(cby_2__1__1_chany_out_188_[0]),
		.chany_out_189_(cby_2__1__1_chany_out_189_[0]),
		.chany_out_190_(cby_2__1__1_chany_out_190_[0]),
		.chany_out_191_(cby_2__1__1_chany_out_191_[0]),
		.chany_out_192_(cby_2__1__1_chany_out_192_[0]),
		.chany_out_193_(cby_2__1__1_chany_out_193_[0]),
		.chany_out_194_(cby_2__1__1_chany_out_194_[0]),
		.chany_out_195_(cby_2__1__1_chany_out_195_[0]),
		.chany_out_196_(cby_2__1__1_chany_out_196_[0]),
		.chany_out_197_(cby_2__1__1_chany_out_197_[0]),
		.chany_out_198_(cby_2__1__1_chany_out_198_[0]),
		.chany_out_199_(cby_2__1__1_chany_out_199_[0]),
		.right_grid_pin_0_(cby_2__1__1_right_grid_pin_0_[0]),
		.left_grid_pin_0_(cby_2__1__1_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_2__1__1_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_2__1__1_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_2__1__1_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_2__1__1_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_2__1__1_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_2__1__1_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_2__1__1_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_2__1__1_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_2__1__1_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_2__1__1_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_2__1__1_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_2__1__1_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_2__1__1_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_2__1__1_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_2__1__1_left_grid_pin_15_[0]),
		.left_grid_pin_16_(cby_2__1__1_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_2__1__1_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_2__1__1_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_2__1__1_left_grid_pin_19_[0]),
		.ccff_tail(cby_2__1__1_ccff_tail[0]));

	direct_interc direct_interc_0_ (
		.in(grid_clb_2_bottom_width_0_height_0__pin_65_[0]),
		.out(direct_interc_0_out[0]));

	direct_interc direct_interc_1_ (
		.in(grid_clb_2_bottom_width_0_height_0__pin_64_[0]),
		.out(direct_interc_1_out[0]));

endmodule
// ----- END Verilog module for fpga_top -----



