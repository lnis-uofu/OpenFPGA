*****************************
*     FPGA SPICE Netlist    *
* Description: Switch Block  [1][1] in FPGA *
*    Author: Xifan TANG     *
* Organization: EPFL/IC/LSI *
* Date: Thu Nov 15 14:26:08 2018
 *
*****************************
***** Switch Box[1][1] Sub-Circuit *****
.subckt sb[1][1] 
***** Inputs/outputs of top side *****
+ 
+ 
+ ***** Inputs/outputs of right side *****
+ 
+ 
+ ***** Inputs/outputs of bottom side *****
+ chany[1][1]_in[0] chany[1][1]_out[1] chany[1][1]_in[2] chany[1][1]_out[3] chany[1][1]_in[4] chany[1][1]_out[5] chany[1][1]_in[6] chany[1][1]_out[7] chany[1][1]_in[8] chany[1][1]_out[9] chany[1][1]_in[10] chany[1][1]_out[11] chany[1][1]_in[12] chany[1][1]_out[13] chany[1][1]_in[14] chany[1][1]_out[15] chany[1][1]_in[16] chany[1][1]_out[17] chany[1][1]_in[18] chany[1][1]_out[19] chany[1][1]_in[20] chany[1][1]_out[21] chany[1][1]_in[22] chany[1][1]_out[23] chany[1][1]_in[24] chany[1][1]_out[25] chany[1][1]_in[26] chany[1][1]_out[27] chany[1][1]_in[28] chany[1][1]_out[29] chany[1][1]_in[30] chany[1][1]_out[31] chany[1][1]_in[32] chany[1][1]_out[33] chany[1][1]_in[34] chany[1][1]_out[35] chany[1][1]_in[36] chany[1][1]_out[37] chany[1][1]_in[38] chany[1][1]_out[39] chany[1][1]_in[40] chany[1][1]_out[41] chany[1][1]_in[42] chany[1][1]_out[43] chany[1][1]_in[44] chany[1][1]_out[45] chany[1][1]_in[46] chany[1][1]_out[47] chany[1][1]_in[48] chany[1][1]_out[49] chany[1][1]_in[50] chany[1][1]_out[51] chany[1][1]_in[52] chany[1][1]_out[53] chany[1][1]_in[54] chany[1][1]_out[55] chany[1][1]_in[56] chany[1][1]_out[57] chany[1][1]_in[58] chany[1][1]_out[59] chany[1][1]_in[60] chany[1][1]_out[61] chany[1][1]_in[62] chany[1][1]_out[63] chany[1][1]_in[64] chany[1][1]_out[65] chany[1][1]_in[66] chany[1][1]_out[67] chany[1][1]_in[68] chany[1][1]_out[69] chany[1][1]_in[70] chany[1][1]_out[71] chany[1][1]_in[72] chany[1][1]_out[73] chany[1][1]_in[74] chany[1][1]_out[75] chany[1][1]_in[76] chany[1][1]_out[77] chany[1][1]_in[78] chany[1][1]_out[79] chany[1][1]_in[80] chany[1][1]_out[81] chany[1][1]_in[82] chany[1][1]_out[83] chany[1][1]_in[84] chany[1][1]_out[85] chany[1][1]_in[86] chany[1][1]_out[87] chany[1][1]_in[88] chany[1][1]_out[89] chany[1][1]_in[90] chany[1][1]_out[91] chany[1][1]_in[92] chany[1][1]_out[93] chany[1][1]_in[94] chany[1][1]_out[95] chany[1][1]_in[96] chany[1][1]_out[97] chany[1][1]_in[98] chany[1][1]_out[99] 
+ grid[2][1]_pin[0][3][1] grid[2][1]_pin[0][3][3] grid[2][1]_pin[0][3][5] grid[2][1]_pin[0][3][7] grid[2][1]_pin[0][3][9] grid[2][1]_pin[0][3][11] grid[2][1]_pin[0][3][13] grid[2][1]_pin[0][3][15] grid[1][1]_pin[0][1][41] grid[1][1]_pin[0][1][45] grid[1][1]_pin[0][1][49] 
+ ***** Inputs/outputs of left side *****
+ chanx[1][1]_in[0] chanx[1][1]_out[1] chanx[1][1]_in[2] chanx[1][1]_out[3] chanx[1][1]_in[4] chanx[1][1]_out[5] chanx[1][1]_in[6] chanx[1][1]_out[7] chanx[1][1]_in[8] chanx[1][1]_out[9] chanx[1][1]_in[10] chanx[1][1]_out[11] chanx[1][1]_in[12] chanx[1][1]_out[13] chanx[1][1]_in[14] chanx[1][1]_out[15] chanx[1][1]_in[16] chanx[1][1]_out[17] chanx[1][1]_in[18] chanx[1][1]_out[19] chanx[1][1]_in[20] chanx[1][1]_out[21] chanx[1][1]_in[22] chanx[1][1]_out[23] chanx[1][1]_in[24] chanx[1][1]_out[25] chanx[1][1]_in[26] chanx[1][1]_out[27] chanx[1][1]_in[28] chanx[1][1]_out[29] chanx[1][1]_in[30] chanx[1][1]_out[31] chanx[1][1]_in[32] chanx[1][1]_out[33] chanx[1][1]_in[34] chanx[1][1]_out[35] chanx[1][1]_in[36] chanx[1][1]_out[37] chanx[1][1]_in[38] chanx[1][1]_out[39] chanx[1][1]_in[40] chanx[1][1]_out[41] chanx[1][1]_in[42] chanx[1][1]_out[43] chanx[1][1]_in[44] chanx[1][1]_out[45] chanx[1][1]_in[46] chanx[1][1]_out[47] chanx[1][1]_in[48] chanx[1][1]_out[49] chanx[1][1]_in[50] chanx[1][1]_out[51] chanx[1][1]_in[52] chanx[1][1]_out[53] chanx[1][1]_in[54] chanx[1][1]_out[55] chanx[1][1]_in[56] chanx[1][1]_out[57] chanx[1][1]_in[58] chanx[1][1]_out[59] chanx[1][1]_in[60] chanx[1][1]_out[61] chanx[1][1]_in[62] chanx[1][1]_out[63] chanx[1][1]_in[64] chanx[1][1]_out[65] chanx[1][1]_in[66] chanx[1][1]_out[67] chanx[1][1]_in[68] chanx[1][1]_out[69] chanx[1][1]_in[70] chanx[1][1]_out[71] chanx[1][1]_in[72] chanx[1][1]_out[73] chanx[1][1]_in[74] chanx[1][1]_out[75] chanx[1][1]_in[76] chanx[1][1]_out[77] chanx[1][1]_in[78] chanx[1][1]_out[79] chanx[1][1]_in[80] chanx[1][1]_out[81] chanx[1][1]_in[82] chanx[1][1]_out[83] chanx[1][1]_in[84] chanx[1][1]_out[85] chanx[1][1]_in[86] chanx[1][1]_out[87] chanx[1][1]_in[88] chanx[1][1]_out[89] chanx[1][1]_in[90] chanx[1][1]_out[91] chanx[1][1]_in[92] chanx[1][1]_out[93] chanx[1][1]_in[94] chanx[1][1]_out[95] chanx[1][1]_in[96] chanx[1][1]_out[97] chanx[1][1]_in[98] chanx[1][1]_out[99] 
+ grid[1][2]_pin[0][2][1] grid[1][2]_pin[0][2][3] grid[1][2]_pin[0][2][5] grid[1][2]_pin[0][2][7] grid[1][2]_pin[0][2][9] grid[1][2]_pin[0][2][11] grid[1][2]_pin[0][2][13] grid[1][2]_pin[0][2][15] grid[1][1]_pin[0][0][40] grid[1][1]_pin[0][0][44] grid[1][1]_pin[0][0][48] 
+ svdd sgnd
***** top side Multiplexers *****
***** right side Multiplexers *****
***** bottom side Multiplexers *****
Xmux_1level_tapbuf_size3[310] grid[1][1]_pin[0][1][41] grid[2][1]_pin[0][3][15] chanx[1][1]_in[2] chany[1][1]_out[1] sram[1962]->outb sram[1962]->out sram[1963]->out sram[1963]->outb sram[1964]->out sram[1964]->outb svdd sgnd mux_1level_tapbuf_size3
***** SRAM bits for MUX[310], level=1, select_path_id=0. *****
*****100*****
Xsram[1962] sram->in sram[1962]->out sram[1962]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1962]->out) 0
.nodeset V(sram[1962]->outb) vsp
Xsram[1963] sram->in sram[1963]->out sram[1963]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1963]->out) 0
.nodeset V(sram[1963]->outb) vsp
Xsram[1964] sram->in sram[1964]->out sram[1964]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1964]->out) 0
.nodeset V(sram[1964]->outb) vsp
Xmux_1level_tapbuf_size3[311] grid[1][1]_pin[0][1][41] grid[2][1]_pin[0][3][15] chanx[1][1]_in[4] chany[1][1]_out[3] sram[1965]->outb sram[1965]->out sram[1966]->out sram[1966]->outb sram[1967]->out sram[1967]->outb svdd sgnd mux_1level_tapbuf_size3
***** SRAM bits for MUX[311], level=1, select_path_id=0. *****
*****100*****
Xsram[1965] sram->in sram[1965]->out sram[1965]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1965]->out) 0
.nodeset V(sram[1965]->outb) vsp
Xsram[1966] sram->in sram[1966]->out sram[1966]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1966]->out) 0
.nodeset V(sram[1966]->outb) vsp
Xsram[1967] sram->in sram[1967]->out sram[1967]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1967]->out) 0
.nodeset V(sram[1967]->outb) vsp
Xmux_1level_tapbuf_size3[312] grid[1][1]_pin[0][1][41] grid[2][1]_pin[0][3][15] chanx[1][1]_in[6] chany[1][1]_out[5] sram[1968]->outb sram[1968]->out sram[1969]->out sram[1969]->outb sram[1970]->out sram[1970]->outb svdd sgnd mux_1level_tapbuf_size3
***** SRAM bits for MUX[312], level=1, select_path_id=0. *****
*****100*****
Xsram[1968] sram->in sram[1968]->out sram[1968]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1968]->out) 0
.nodeset V(sram[1968]->outb) vsp
Xsram[1969] sram->in sram[1969]->out sram[1969]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1969]->out) 0
.nodeset V(sram[1969]->outb) vsp
Xsram[1970] sram->in sram[1970]->out sram[1970]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1970]->out) 0
.nodeset V(sram[1970]->outb) vsp
Xmux_1level_tapbuf_size3[313] grid[1][1]_pin[0][1][41] grid[2][1]_pin[0][3][15] chanx[1][1]_in[8] chany[1][1]_out[7] sram[1971]->outb sram[1971]->out sram[1972]->out sram[1972]->outb sram[1973]->out sram[1973]->outb svdd sgnd mux_1level_tapbuf_size3
***** SRAM bits for MUX[313], level=1, select_path_id=0. *****
*****100*****
Xsram[1971] sram->in sram[1971]->out sram[1971]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1971]->out) 0
.nodeset V(sram[1971]->outb) vsp
Xsram[1972] sram->in sram[1972]->out sram[1972]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1972]->out) 0
.nodeset V(sram[1972]->outb) vsp
Xsram[1973] sram->in sram[1973]->out sram[1973]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1973]->out) 0
.nodeset V(sram[1973]->outb) vsp
Xmux_1level_tapbuf_size3[314] grid[1][1]_pin[0][1][41] grid[2][1]_pin[0][3][15] chanx[1][1]_in[10] chany[1][1]_out[9] sram[1974]->outb sram[1974]->out sram[1975]->out sram[1975]->outb sram[1976]->out sram[1976]->outb svdd sgnd mux_1level_tapbuf_size3
***** SRAM bits for MUX[314], level=1, select_path_id=0. *****
*****100*****
Xsram[1974] sram->in sram[1974]->out sram[1974]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1974]->out) 0
.nodeset V(sram[1974]->outb) vsp
Xsram[1975] sram->in sram[1975]->out sram[1975]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1975]->out) 0
.nodeset V(sram[1975]->outb) vsp
Xsram[1976] sram->in sram[1976]->out sram[1976]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1976]->out) 0
.nodeset V(sram[1976]->outb) vsp
Xmux_1level_tapbuf_size2[315] grid[1][1]_pin[0][1][45] chanx[1][1]_in[12] chany[1][1]_out[11] sram[1977]->outb sram[1977]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[315], level=1, select_path_id=0. *****
*****1*****
Xsram[1977] sram->in sram[1977]->out sram[1977]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1977]->out) 0
.nodeset V(sram[1977]->outb) vsp
Xmux_1level_tapbuf_size2[316] grid[1][1]_pin[0][1][45] chanx[1][1]_in[14] chany[1][1]_out[13] sram[1978]->outb sram[1978]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[316], level=1, select_path_id=0. *****
*****1*****
Xsram[1978] sram->in sram[1978]->out sram[1978]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1978]->out) 0
.nodeset V(sram[1978]->outb) vsp
Xmux_1level_tapbuf_size2[317] grid[1][1]_pin[0][1][45] chanx[1][1]_in[16] chany[1][1]_out[15] sram[1979]->outb sram[1979]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[317], level=1, select_path_id=0. *****
*****1*****
Xsram[1979] sram->in sram[1979]->out sram[1979]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1979]->out) 0
.nodeset V(sram[1979]->outb) vsp
Xmux_1level_tapbuf_size2[318] grid[1][1]_pin[0][1][45] chanx[1][1]_in[18] chany[1][1]_out[17] sram[1980]->outb sram[1980]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[318], level=1, select_path_id=0. *****
*****1*****
Xsram[1980] sram->in sram[1980]->out sram[1980]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1980]->out) 0
.nodeset V(sram[1980]->outb) vsp
Xmux_1level_tapbuf_size2[319] grid[1][1]_pin[0][1][45] chanx[1][1]_in[20] chany[1][1]_out[19] sram[1981]->outb sram[1981]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[319], level=1, select_path_id=0. *****
*****1*****
Xsram[1981] sram->in sram[1981]->out sram[1981]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1981]->out) 0
.nodeset V(sram[1981]->outb) vsp
Xmux_1level_tapbuf_size2[320] grid[1][1]_pin[0][1][49] chanx[1][1]_in[22] chany[1][1]_out[21] sram[1982]->outb sram[1982]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[320], level=1, select_path_id=0. *****
*****1*****
Xsram[1982] sram->in sram[1982]->out sram[1982]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1982]->out) 0
.nodeset V(sram[1982]->outb) vsp
Xmux_1level_tapbuf_size2[321] grid[1][1]_pin[0][1][49] chanx[1][1]_in[24] chany[1][1]_out[23] sram[1983]->outb sram[1983]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[321], level=1, select_path_id=0. *****
*****1*****
Xsram[1983] sram->in sram[1983]->out sram[1983]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1983]->out) 0
.nodeset V(sram[1983]->outb) vsp
Xmux_1level_tapbuf_size2[322] grid[1][1]_pin[0][1][49] chanx[1][1]_in[26] chany[1][1]_out[25] sram[1984]->outb sram[1984]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[322], level=1, select_path_id=0. *****
*****1*****
Xsram[1984] sram->in sram[1984]->out sram[1984]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1984]->out) 0
.nodeset V(sram[1984]->outb) vsp
Xmux_1level_tapbuf_size2[323] grid[1][1]_pin[0][1][49] chanx[1][1]_in[28] chany[1][1]_out[27] sram[1985]->outb sram[1985]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[323], level=1, select_path_id=0. *****
*****1*****
Xsram[1985] sram->in sram[1985]->out sram[1985]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1985]->out) 0
.nodeset V(sram[1985]->outb) vsp
Xmux_1level_tapbuf_size2[324] grid[1][1]_pin[0][1][49] chanx[1][1]_in[30] chany[1][1]_out[29] sram[1986]->outb sram[1986]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[324], level=1, select_path_id=0. *****
*****1*****
Xsram[1986] sram->in sram[1986]->out sram[1986]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1986]->out) 0
.nodeset V(sram[1986]->outb) vsp
Xmux_1level_tapbuf_size2[325] grid[2][1]_pin[0][3][1] chanx[1][1]_in[32] chany[1][1]_out[31] sram[1987]->outb sram[1987]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[325], level=1, select_path_id=0. *****
*****1*****
Xsram[1987] sram->in sram[1987]->out sram[1987]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1987]->out) 0
.nodeset V(sram[1987]->outb) vsp
Xmux_1level_tapbuf_size2[326] grid[2][1]_pin[0][3][1] chanx[1][1]_in[34] chany[1][1]_out[33] sram[1988]->outb sram[1988]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[326], level=1, select_path_id=0. *****
*****1*****
Xsram[1988] sram->in sram[1988]->out sram[1988]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1988]->out) 0
.nodeset V(sram[1988]->outb) vsp
Xmux_1level_tapbuf_size2[327] grid[2][1]_pin[0][3][1] chanx[1][1]_in[36] chany[1][1]_out[35] sram[1989]->outb sram[1989]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[327], level=1, select_path_id=0. *****
*****1*****
Xsram[1989] sram->in sram[1989]->out sram[1989]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1989]->out) 0
.nodeset V(sram[1989]->outb) vsp
Xmux_1level_tapbuf_size2[328] grid[2][1]_pin[0][3][1] chanx[1][1]_in[38] chany[1][1]_out[37] sram[1990]->outb sram[1990]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[328], level=1, select_path_id=0. *****
*****1*****
Xsram[1990] sram->in sram[1990]->out sram[1990]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1990]->out) 0
.nodeset V(sram[1990]->outb) vsp
Xmux_1level_tapbuf_size2[329] grid[2][1]_pin[0][3][1] chanx[1][1]_in[40] chany[1][1]_out[39] sram[1991]->outb sram[1991]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[329], level=1, select_path_id=0. *****
*****1*****
Xsram[1991] sram->in sram[1991]->out sram[1991]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1991]->out) 0
.nodeset V(sram[1991]->outb) vsp
Xmux_1level_tapbuf_size2[330] grid[2][1]_pin[0][3][3] chanx[1][1]_in[42] chany[1][1]_out[41] sram[1992]->outb sram[1992]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[330], level=1, select_path_id=0. *****
*****1*****
Xsram[1992] sram->in sram[1992]->out sram[1992]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1992]->out) 0
.nodeset V(sram[1992]->outb) vsp
Xmux_1level_tapbuf_size2[331] grid[2][1]_pin[0][3][3] chanx[1][1]_in[44] chany[1][1]_out[43] sram[1993]->outb sram[1993]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[331], level=1, select_path_id=0. *****
*****1*****
Xsram[1993] sram->in sram[1993]->out sram[1993]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1993]->out) 0
.nodeset V(sram[1993]->outb) vsp
Xmux_1level_tapbuf_size2[332] grid[2][1]_pin[0][3][3] chanx[1][1]_in[46] chany[1][1]_out[45] sram[1994]->outb sram[1994]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[332], level=1, select_path_id=0. *****
*****1*****
Xsram[1994] sram->in sram[1994]->out sram[1994]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1994]->out) 0
.nodeset V(sram[1994]->outb) vsp
Xmux_1level_tapbuf_size2[333] grid[2][1]_pin[0][3][3] chanx[1][1]_in[48] chany[1][1]_out[47] sram[1995]->outb sram[1995]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[333], level=1, select_path_id=0. *****
*****1*****
Xsram[1995] sram->in sram[1995]->out sram[1995]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1995]->out) 0
.nodeset V(sram[1995]->outb) vsp
Xmux_1level_tapbuf_size2[334] grid[2][1]_pin[0][3][3] chanx[1][1]_in[50] chany[1][1]_out[49] sram[1996]->outb sram[1996]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[334], level=1, select_path_id=0. *****
*****1*****
Xsram[1996] sram->in sram[1996]->out sram[1996]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1996]->out) 0
.nodeset V(sram[1996]->outb) vsp
Xmux_1level_tapbuf_size2[335] grid[2][1]_pin[0][3][5] chanx[1][1]_in[52] chany[1][1]_out[51] sram[1997]->outb sram[1997]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[335], level=1, select_path_id=0. *****
*****1*****
Xsram[1997] sram->in sram[1997]->out sram[1997]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1997]->out) 0
.nodeset V(sram[1997]->outb) vsp
Xmux_1level_tapbuf_size2[336] grid[2][1]_pin[0][3][5] chanx[1][1]_in[54] chany[1][1]_out[53] sram[1998]->outb sram[1998]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[336], level=1, select_path_id=0. *****
*****1*****
Xsram[1998] sram->in sram[1998]->out sram[1998]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1998]->out) 0
.nodeset V(sram[1998]->outb) vsp
Xmux_1level_tapbuf_size2[337] grid[2][1]_pin[0][3][5] chanx[1][1]_in[56] chany[1][1]_out[55] sram[1999]->outb sram[1999]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[337], level=1, select_path_id=0. *****
*****1*****
Xsram[1999] sram->in sram[1999]->out sram[1999]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1999]->out) 0
.nodeset V(sram[1999]->outb) vsp
Xmux_1level_tapbuf_size2[338] grid[2][1]_pin[0][3][5] chanx[1][1]_in[58] chany[1][1]_out[57] sram[2000]->outb sram[2000]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[338], level=1, select_path_id=0. *****
*****1*****
Xsram[2000] sram->in sram[2000]->out sram[2000]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2000]->out) 0
.nodeset V(sram[2000]->outb) vsp
Xmux_1level_tapbuf_size2[339] grid[2][1]_pin[0][3][5] chanx[1][1]_in[60] chany[1][1]_out[59] sram[2001]->outb sram[2001]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[339], level=1, select_path_id=0. *****
*****1*****
Xsram[2001] sram->in sram[2001]->out sram[2001]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2001]->out) 0
.nodeset V(sram[2001]->outb) vsp
Xmux_1level_tapbuf_size2[340] grid[2][1]_pin[0][3][7] chanx[1][1]_in[62] chany[1][1]_out[61] sram[2002]->outb sram[2002]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[340], level=1, select_path_id=0. *****
*****1*****
Xsram[2002] sram->in sram[2002]->out sram[2002]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2002]->out) 0
.nodeset V(sram[2002]->outb) vsp
Xmux_1level_tapbuf_size2[341] grid[2][1]_pin[0][3][7] chanx[1][1]_in[64] chany[1][1]_out[63] sram[2003]->outb sram[2003]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[341], level=1, select_path_id=0. *****
*****1*****
Xsram[2003] sram->in sram[2003]->out sram[2003]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2003]->out) 0
.nodeset V(sram[2003]->outb) vsp
Xmux_1level_tapbuf_size2[342] grid[2][1]_pin[0][3][7] chanx[1][1]_in[66] chany[1][1]_out[65] sram[2004]->outb sram[2004]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[342], level=1, select_path_id=0. *****
*****1*****
Xsram[2004] sram->in sram[2004]->out sram[2004]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2004]->out) 0
.nodeset V(sram[2004]->outb) vsp
Xmux_1level_tapbuf_size2[343] grid[2][1]_pin[0][3][7] chanx[1][1]_in[68] chany[1][1]_out[67] sram[2005]->outb sram[2005]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[343], level=1, select_path_id=0. *****
*****1*****
Xsram[2005] sram->in sram[2005]->out sram[2005]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2005]->out) 0
.nodeset V(sram[2005]->outb) vsp
Xmux_1level_tapbuf_size2[344] grid[2][1]_pin[0][3][7] chanx[1][1]_in[70] chany[1][1]_out[69] sram[2006]->outb sram[2006]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[344], level=1, select_path_id=0. *****
*****1*****
Xsram[2006] sram->in sram[2006]->out sram[2006]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2006]->out) 0
.nodeset V(sram[2006]->outb) vsp
Xmux_1level_tapbuf_size2[345] grid[2][1]_pin[0][3][9] chanx[1][1]_in[72] chany[1][1]_out[71] sram[2007]->outb sram[2007]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[345], level=1, select_path_id=0. *****
*****1*****
Xsram[2007] sram->in sram[2007]->out sram[2007]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2007]->out) 0
.nodeset V(sram[2007]->outb) vsp
Xmux_1level_tapbuf_size2[346] grid[2][1]_pin[0][3][9] chanx[1][1]_in[74] chany[1][1]_out[73] sram[2008]->outb sram[2008]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[346], level=1, select_path_id=0. *****
*****1*****
Xsram[2008] sram->in sram[2008]->out sram[2008]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2008]->out) 0
.nodeset V(sram[2008]->outb) vsp
Xmux_1level_tapbuf_size2[347] grid[2][1]_pin[0][3][9] chanx[1][1]_in[76] chany[1][1]_out[75] sram[2009]->outb sram[2009]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[347], level=1, select_path_id=0. *****
*****1*****
Xsram[2009] sram->in sram[2009]->out sram[2009]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2009]->out) 0
.nodeset V(sram[2009]->outb) vsp
Xmux_1level_tapbuf_size2[348] grid[2][1]_pin[0][3][9] chanx[1][1]_in[78] chany[1][1]_out[77] sram[2010]->outb sram[2010]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[348], level=1, select_path_id=0. *****
*****1*****
Xsram[2010] sram->in sram[2010]->out sram[2010]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2010]->out) 0
.nodeset V(sram[2010]->outb) vsp
Xmux_1level_tapbuf_size2[349] grid[2][1]_pin[0][3][9] chanx[1][1]_in[80] chany[1][1]_out[79] sram[2011]->outb sram[2011]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[349], level=1, select_path_id=0. *****
*****1*****
Xsram[2011] sram->in sram[2011]->out sram[2011]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2011]->out) 0
.nodeset V(sram[2011]->outb) vsp
Xmux_1level_tapbuf_size2[350] grid[2][1]_pin[0][3][11] chanx[1][1]_in[82] chany[1][1]_out[81] sram[2012]->outb sram[2012]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[350], level=1, select_path_id=0. *****
*****1*****
Xsram[2012] sram->in sram[2012]->out sram[2012]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2012]->out) 0
.nodeset V(sram[2012]->outb) vsp
Xmux_1level_tapbuf_size2[351] grid[2][1]_pin[0][3][11] chanx[1][1]_in[84] chany[1][1]_out[83] sram[2013]->outb sram[2013]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[351], level=1, select_path_id=0. *****
*****1*****
Xsram[2013] sram->in sram[2013]->out sram[2013]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2013]->out) 0
.nodeset V(sram[2013]->outb) vsp
Xmux_1level_tapbuf_size2[352] grid[2][1]_pin[0][3][11] chanx[1][1]_in[86] chany[1][1]_out[85] sram[2014]->outb sram[2014]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[352], level=1, select_path_id=0. *****
*****1*****
Xsram[2014] sram->in sram[2014]->out sram[2014]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2014]->out) 0
.nodeset V(sram[2014]->outb) vsp
Xmux_1level_tapbuf_size2[353] grid[2][1]_pin[0][3][11] chanx[1][1]_in[88] chany[1][1]_out[87] sram[2015]->outb sram[2015]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[353], level=1, select_path_id=0. *****
*****1*****
Xsram[2015] sram->in sram[2015]->out sram[2015]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2015]->out) 0
.nodeset V(sram[2015]->outb) vsp
Xmux_1level_tapbuf_size2[354] grid[2][1]_pin[0][3][11] chanx[1][1]_in[90] chany[1][1]_out[89] sram[2016]->outb sram[2016]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[354], level=1, select_path_id=0. *****
*****1*****
Xsram[2016] sram->in sram[2016]->out sram[2016]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2016]->out) 0
.nodeset V(sram[2016]->outb) vsp
Xmux_1level_tapbuf_size2[355] grid[2][1]_pin[0][3][13] chanx[1][1]_in[92] chany[1][1]_out[91] sram[2017]->outb sram[2017]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[355], level=1, select_path_id=0. *****
*****1*****
Xsram[2017] sram->in sram[2017]->out sram[2017]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2017]->out) 0
.nodeset V(sram[2017]->outb) vsp
Xmux_1level_tapbuf_size2[356] grid[2][1]_pin[0][3][13] chanx[1][1]_in[94] chany[1][1]_out[93] sram[2018]->outb sram[2018]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[356], level=1, select_path_id=0. *****
*****1*****
Xsram[2018] sram->in sram[2018]->out sram[2018]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2018]->out) 0
.nodeset V(sram[2018]->outb) vsp
Xmux_1level_tapbuf_size2[357] grid[2][1]_pin[0][3][13] chanx[1][1]_in[96] chany[1][1]_out[95] sram[2019]->outb sram[2019]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[357], level=1, select_path_id=0. *****
*****1*****
Xsram[2019] sram->in sram[2019]->out sram[2019]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2019]->out) 0
.nodeset V(sram[2019]->outb) vsp
Xmux_1level_tapbuf_size2[358] grid[2][1]_pin[0][3][13] chanx[1][1]_in[98] chany[1][1]_out[97] sram[2020]->outb sram[2020]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[358], level=1, select_path_id=0. *****
*****1*****
Xsram[2020] sram->in sram[2020]->out sram[2020]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2020]->out) 0
.nodeset V(sram[2020]->outb) vsp
Xmux_1level_tapbuf_size2[359] grid[2][1]_pin[0][3][13] chanx[1][1]_in[0] chany[1][1]_out[99] sram[2021]->outb sram[2021]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[359], level=1, select_path_id=0. *****
*****1*****
Xsram[2021] sram->in sram[2021]->out sram[2021]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2021]->out) 0
.nodeset V(sram[2021]->outb) vsp
***** left side Multiplexers *****
Xmux_1level_tapbuf_size3[360] grid[1][1]_pin[0][0][40] grid[1][2]_pin[0][2][15] chany[1][1]_in[98] chanx[1][1]_out[1] sram[2022]->outb sram[2022]->out sram[2023]->out sram[2023]->outb sram[2024]->out sram[2024]->outb svdd sgnd mux_1level_tapbuf_size3
***** SRAM bits for MUX[360], level=1, select_path_id=0. *****
*****100*****
Xsram[2022] sram->in sram[2022]->out sram[2022]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2022]->out) 0
.nodeset V(sram[2022]->outb) vsp
Xsram[2023] sram->in sram[2023]->out sram[2023]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2023]->out) 0
.nodeset V(sram[2023]->outb) vsp
Xsram[2024] sram->in sram[2024]->out sram[2024]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2024]->out) 0
.nodeset V(sram[2024]->outb) vsp
Xmux_1level_tapbuf_size3[361] grid[1][1]_pin[0][0][40] grid[1][2]_pin[0][2][15] chany[1][1]_in[0] chanx[1][1]_out[3] sram[2025]->outb sram[2025]->out sram[2026]->out sram[2026]->outb sram[2027]->out sram[2027]->outb svdd sgnd mux_1level_tapbuf_size3
***** SRAM bits for MUX[361], level=1, select_path_id=0. *****
*****100*****
Xsram[2025] sram->in sram[2025]->out sram[2025]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2025]->out) 0
.nodeset V(sram[2025]->outb) vsp
Xsram[2026] sram->in sram[2026]->out sram[2026]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2026]->out) 0
.nodeset V(sram[2026]->outb) vsp
Xsram[2027] sram->in sram[2027]->out sram[2027]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2027]->out) 0
.nodeset V(sram[2027]->outb) vsp
Xmux_1level_tapbuf_size3[362] grid[1][1]_pin[0][0][40] grid[1][2]_pin[0][2][15] chany[1][1]_in[2] chanx[1][1]_out[5] sram[2028]->outb sram[2028]->out sram[2029]->out sram[2029]->outb sram[2030]->out sram[2030]->outb svdd sgnd mux_1level_tapbuf_size3
***** SRAM bits for MUX[362], level=1, select_path_id=0. *****
*****100*****
Xsram[2028] sram->in sram[2028]->out sram[2028]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2028]->out) 0
.nodeset V(sram[2028]->outb) vsp
Xsram[2029] sram->in sram[2029]->out sram[2029]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2029]->out) 0
.nodeset V(sram[2029]->outb) vsp
Xsram[2030] sram->in sram[2030]->out sram[2030]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2030]->out) 0
.nodeset V(sram[2030]->outb) vsp
Xmux_1level_tapbuf_size3[363] grid[1][1]_pin[0][0][40] grid[1][2]_pin[0][2][15] chany[1][1]_in[4] chanx[1][1]_out[7] sram[2031]->outb sram[2031]->out sram[2032]->out sram[2032]->outb sram[2033]->out sram[2033]->outb svdd sgnd mux_1level_tapbuf_size3
***** SRAM bits for MUX[363], level=1, select_path_id=0. *****
*****100*****
Xsram[2031] sram->in sram[2031]->out sram[2031]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2031]->out) 0
.nodeset V(sram[2031]->outb) vsp
Xsram[2032] sram->in sram[2032]->out sram[2032]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2032]->out) 0
.nodeset V(sram[2032]->outb) vsp
Xsram[2033] sram->in sram[2033]->out sram[2033]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2033]->out) 0
.nodeset V(sram[2033]->outb) vsp
Xmux_1level_tapbuf_size3[364] grid[1][1]_pin[0][0][40] grid[1][2]_pin[0][2][15] chany[1][1]_in[6] chanx[1][1]_out[9] sram[2034]->outb sram[2034]->out sram[2035]->out sram[2035]->outb sram[2036]->out sram[2036]->outb svdd sgnd mux_1level_tapbuf_size3
***** SRAM bits for MUX[364], level=1, select_path_id=0. *****
*****100*****
Xsram[2034] sram->in sram[2034]->out sram[2034]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2034]->out) 0
.nodeset V(sram[2034]->outb) vsp
Xsram[2035] sram->in sram[2035]->out sram[2035]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2035]->out) 0
.nodeset V(sram[2035]->outb) vsp
Xsram[2036] sram->in sram[2036]->out sram[2036]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2036]->out) 0
.nodeset V(sram[2036]->outb) vsp
Xmux_1level_tapbuf_size2[365] grid[1][1]_pin[0][0][44] chany[1][1]_in[8] chanx[1][1]_out[11] sram[2037]->outb sram[2037]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[365], level=1, select_path_id=0. *****
*****1*****
Xsram[2037] sram->in sram[2037]->out sram[2037]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2037]->out) 0
.nodeset V(sram[2037]->outb) vsp
Xmux_1level_tapbuf_size2[366] grid[1][1]_pin[0][0][44] chany[1][1]_in[10] chanx[1][1]_out[13] sram[2038]->outb sram[2038]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[366], level=1, select_path_id=0. *****
*****1*****
Xsram[2038] sram->in sram[2038]->out sram[2038]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2038]->out) 0
.nodeset V(sram[2038]->outb) vsp
Xmux_1level_tapbuf_size2[367] grid[1][1]_pin[0][0][44] chany[1][1]_in[12] chanx[1][1]_out[15] sram[2039]->outb sram[2039]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[367], level=1, select_path_id=0. *****
*****1*****
Xsram[2039] sram->in sram[2039]->out sram[2039]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2039]->out) 0
.nodeset V(sram[2039]->outb) vsp
Xmux_1level_tapbuf_size2[368] grid[1][1]_pin[0][0][44] chany[1][1]_in[14] chanx[1][1]_out[17] sram[2040]->outb sram[2040]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[368], level=1, select_path_id=0. *****
*****1*****
Xsram[2040] sram->in sram[2040]->out sram[2040]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2040]->out) 0
.nodeset V(sram[2040]->outb) vsp
Xmux_1level_tapbuf_size2[369] grid[1][1]_pin[0][0][44] chany[1][1]_in[16] chanx[1][1]_out[19] sram[2041]->outb sram[2041]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[369], level=1, select_path_id=0. *****
*****1*****
Xsram[2041] sram->in sram[2041]->out sram[2041]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2041]->out) 0
.nodeset V(sram[2041]->outb) vsp
Xmux_1level_tapbuf_size2[370] grid[1][1]_pin[0][0][48] chany[1][1]_in[18] chanx[1][1]_out[21] sram[2042]->outb sram[2042]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[370], level=1, select_path_id=0. *****
*****1*****
Xsram[2042] sram->in sram[2042]->out sram[2042]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2042]->out) 0
.nodeset V(sram[2042]->outb) vsp
Xmux_1level_tapbuf_size2[371] grid[1][1]_pin[0][0][48] chany[1][1]_in[20] chanx[1][1]_out[23] sram[2043]->outb sram[2043]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[371], level=1, select_path_id=0. *****
*****1*****
Xsram[2043] sram->in sram[2043]->out sram[2043]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2043]->out) 0
.nodeset V(sram[2043]->outb) vsp
Xmux_1level_tapbuf_size2[372] grid[1][1]_pin[0][0][48] chany[1][1]_in[22] chanx[1][1]_out[25] sram[2044]->outb sram[2044]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[372], level=1, select_path_id=0. *****
*****1*****
Xsram[2044] sram->in sram[2044]->out sram[2044]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2044]->out) 0
.nodeset V(sram[2044]->outb) vsp
Xmux_1level_tapbuf_size2[373] grid[1][1]_pin[0][0][48] chany[1][1]_in[24] chanx[1][1]_out[27] sram[2045]->outb sram[2045]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[373], level=1, select_path_id=0. *****
*****1*****
Xsram[2045] sram->in sram[2045]->out sram[2045]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2045]->out) 0
.nodeset V(sram[2045]->outb) vsp
Xmux_1level_tapbuf_size2[374] grid[1][1]_pin[0][0][48] chany[1][1]_in[26] chanx[1][1]_out[29] sram[2046]->outb sram[2046]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[374], level=1, select_path_id=0. *****
*****1*****
Xsram[2046] sram->in sram[2046]->out sram[2046]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2046]->out) 0
.nodeset V(sram[2046]->outb) vsp
Xmux_1level_tapbuf_size2[375] grid[1][2]_pin[0][2][1] chany[1][1]_in[28] chanx[1][1]_out[31] sram[2047]->outb sram[2047]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[375], level=1, select_path_id=0. *****
*****1*****
Xsram[2047] sram->in sram[2047]->out sram[2047]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2047]->out) 0
.nodeset V(sram[2047]->outb) vsp
Xmux_1level_tapbuf_size2[376] grid[1][2]_pin[0][2][1] chany[1][1]_in[30] chanx[1][1]_out[33] sram[2048]->outb sram[2048]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[376], level=1, select_path_id=0. *****
*****1*****
Xsram[2048] sram->in sram[2048]->out sram[2048]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2048]->out) 0
.nodeset V(sram[2048]->outb) vsp
Xmux_1level_tapbuf_size2[377] grid[1][2]_pin[0][2][1] chany[1][1]_in[32] chanx[1][1]_out[35] sram[2049]->outb sram[2049]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[377], level=1, select_path_id=0. *****
*****1*****
Xsram[2049] sram->in sram[2049]->out sram[2049]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2049]->out) 0
.nodeset V(sram[2049]->outb) vsp
Xmux_1level_tapbuf_size2[378] grid[1][2]_pin[0][2][1] chany[1][1]_in[34] chanx[1][1]_out[37] sram[2050]->outb sram[2050]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[378], level=1, select_path_id=0. *****
*****1*****
Xsram[2050] sram->in sram[2050]->out sram[2050]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2050]->out) 0
.nodeset V(sram[2050]->outb) vsp
Xmux_1level_tapbuf_size2[379] grid[1][2]_pin[0][2][1] chany[1][1]_in[36] chanx[1][1]_out[39] sram[2051]->outb sram[2051]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[379], level=1, select_path_id=0. *****
*****1*****
Xsram[2051] sram->in sram[2051]->out sram[2051]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2051]->out) 0
.nodeset V(sram[2051]->outb) vsp
Xmux_1level_tapbuf_size2[380] grid[1][2]_pin[0][2][3] chany[1][1]_in[38] chanx[1][1]_out[41] sram[2052]->outb sram[2052]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[380], level=1, select_path_id=0. *****
*****1*****
Xsram[2052] sram->in sram[2052]->out sram[2052]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2052]->out) 0
.nodeset V(sram[2052]->outb) vsp
Xmux_1level_tapbuf_size2[381] grid[1][2]_pin[0][2][3] chany[1][1]_in[40] chanx[1][1]_out[43] sram[2053]->outb sram[2053]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[381], level=1, select_path_id=0. *****
*****1*****
Xsram[2053] sram->in sram[2053]->out sram[2053]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2053]->out) 0
.nodeset V(sram[2053]->outb) vsp
Xmux_1level_tapbuf_size2[382] grid[1][2]_pin[0][2][3] chany[1][1]_in[42] chanx[1][1]_out[45] sram[2054]->outb sram[2054]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[382], level=1, select_path_id=0. *****
*****1*****
Xsram[2054] sram->in sram[2054]->out sram[2054]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2054]->out) 0
.nodeset V(sram[2054]->outb) vsp
Xmux_1level_tapbuf_size2[383] grid[1][2]_pin[0][2][3] chany[1][1]_in[44] chanx[1][1]_out[47] sram[2055]->outb sram[2055]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[383], level=1, select_path_id=0. *****
*****1*****
Xsram[2055] sram->in sram[2055]->out sram[2055]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2055]->out) 0
.nodeset V(sram[2055]->outb) vsp
Xmux_1level_tapbuf_size2[384] grid[1][2]_pin[0][2][3] chany[1][1]_in[46] chanx[1][1]_out[49] sram[2056]->outb sram[2056]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[384], level=1, select_path_id=0. *****
*****1*****
Xsram[2056] sram->in sram[2056]->out sram[2056]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2056]->out) 0
.nodeset V(sram[2056]->outb) vsp
Xmux_1level_tapbuf_size2[385] grid[1][2]_pin[0][2][5] chany[1][1]_in[48] chanx[1][1]_out[51] sram[2057]->outb sram[2057]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[385], level=1, select_path_id=0. *****
*****1*****
Xsram[2057] sram->in sram[2057]->out sram[2057]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2057]->out) 0
.nodeset V(sram[2057]->outb) vsp
Xmux_1level_tapbuf_size2[386] grid[1][2]_pin[0][2][5] chany[1][1]_in[50] chanx[1][1]_out[53] sram[2058]->outb sram[2058]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[386], level=1, select_path_id=0. *****
*****1*****
Xsram[2058] sram->in sram[2058]->out sram[2058]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2058]->out) 0
.nodeset V(sram[2058]->outb) vsp
Xmux_1level_tapbuf_size2[387] grid[1][2]_pin[0][2][5] chany[1][1]_in[52] chanx[1][1]_out[55] sram[2059]->outb sram[2059]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[387], level=1, select_path_id=0. *****
*****1*****
Xsram[2059] sram->in sram[2059]->out sram[2059]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2059]->out) 0
.nodeset V(sram[2059]->outb) vsp
Xmux_1level_tapbuf_size2[388] grid[1][2]_pin[0][2][5] chany[1][1]_in[54] chanx[1][1]_out[57] sram[2060]->outb sram[2060]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[388], level=1, select_path_id=0. *****
*****1*****
Xsram[2060] sram->in sram[2060]->out sram[2060]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2060]->out) 0
.nodeset V(sram[2060]->outb) vsp
Xmux_1level_tapbuf_size2[389] grid[1][2]_pin[0][2][5] chany[1][1]_in[56] chanx[1][1]_out[59] sram[2061]->outb sram[2061]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[389], level=1, select_path_id=0. *****
*****1*****
Xsram[2061] sram->in sram[2061]->out sram[2061]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2061]->out) 0
.nodeset V(sram[2061]->outb) vsp
Xmux_1level_tapbuf_size2[390] grid[1][2]_pin[0][2][7] chany[1][1]_in[58] chanx[1][1]_out[61] sram[2062]->outb sram[2062]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[390], level=1, select_path_id=0. *****
*****1*****
Xsram[2062] sram->in sram[2062]->out sram[2062]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2062]->out) 0
.nodeset V(sram[2062]->outb) vsp
Xmux_1level_tapbuf_size2[391] grid[1][2]_pin[0][2][7] chany[1][1]_in[60] chanx[1][1]_out[63] sram[2063]->outb sram[2063]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[391], level=1, select_path_id=0. *****
*****1*****
Xsram[2063] sram->in sram[2063]->out sram[2063]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2063]->out) 0
.nodeset V(sram[2063]->outb) vsp
Xmux_1level_tapbuf_size2[392] grid[1][2]_pin[0][2][7] chany[1][1]_in[62] chanx[1][1]_out[65] sram[2064]->outb sram[2064]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[392], level=1, select_path_id=0. *****
*****1*****
Xsram[2064] sram->in sram[2064]->out sram[2064]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2064]->out) 0
.nodeset V(sram[2064]->outb) vsp
Xmux_1level_tapbuf_size2[393] grid[1][2]_pin[0][2][7] chany[1][1]_in[64] chanx[1][1]_out[67] sram[2065]->outb sram[2065]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[393], level=1, select_path_id=0. *****
*****1*****
Xsram[2065] sram->in sram[2065]->out sram[2065]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2065]->out) 0
.nodeset V(sram[2065]->outb) vsp
Xmux_1level_tapbuf_size2[394] grid[1][2]_pin[0][2][7] chany[1][1]_in[66] chanx[1][1]_out[69] sram[2066]->outb sram[2066]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[394], level=1, select_path_id=0. *****
*****1*****
Xsram[2066] sram->in sram[2066]->out sram[2066]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2066]->out) 0
.nodeset V(sram[2066]->outb) vsp
Xmux_1level_tapbuf_size2[395] grid[1][2]_pin[0][2][9] chany[1][1]_in[68] chanx[1][1]_out[71] sram[2067]->outb sram[2067]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[395], level=1, select_path_id=0. *****
*****1*****
Xsram[2067] sram->in sram[2067]->out sram[2067]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2067]->out) 0
.nodeset V(sram[2067]->outb) vsp
Xmux_1level_tapbuf_size2[396] grid[1][2]_pin[0][2][9] chany[1][1]_in[70] chanx[1][1]_out[73] sram[2068]->outb sram[2068]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[396], level=1, select_path_id=0. *****
*****1*****
Xsram[2068] sram->in sram[2068]->out sram[2068]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2068]->out) 0
.nodeset V(sram[2068]->outb) vsp
Xmux_1level_tapbuf_size2[397] grid[1][2]_pin[0][2][9] chany[1][1]_in[72] chanx[1][1]_out[75] sram[2069]->outb sram[2069]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[397], level=1, select_path_id=0. *****
*****1*****
Xsram[2069] sram->in sram[2069]->out sram[2069]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2069]->out) 0
.nodeset V(sram[2069]->outb) vsp
Xmux_1level_tapbuf_size2[398] grid[1][2]_pin[0][2][9] chany[1][1]_in[74] chanx[1][1]_out[77] sram[2070]->outb sram[2070]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[398], level=1, select_path_id=0. *****
*****1*****
Xsram[2070] sram->in sram[2070]->out sram[2070]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2070]->out) 0
.nodeset V(sram[2070]->outb) vsp
Xmux_1level_tapbuf_size2[399] grid[1][2]_pin[0][2][9] chany[1][1]_in[76] chanx[1][1]_out[79] sram[2071]->outb sram[2071]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[399], level=1, select_path_id=0. *****
*****1*****
Xsram[2071] sram->in sram[2071]->out sram[2071]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2071]->out) 0
.nodeset V(sram[2071]->outb) vsp
Xmux_1level_tapbuf_size2[400] grid[1][2]_pin[0][2][11] chany[1][1]_in[78] chanx[1][1]_out[81] sram[2072]->outb sram[2072]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[400], level=1, select_path_id=0. *****
*****1*****
Xsram[2072] sram->in sram[2072]->out sram[2072]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2072]->out) 0
.nodeset V(sram[2072]->outb) vsp
Xmux_1level_tapbuf_size2[401] grid[1][2]_pin[0][2][11] chany[1][1]_in[80] chanx[1][1]_out[83] sram[2073]->outb sram[2073]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[401], level=1, select_path_id=0. *****
*****1*****
Xsram[2073] sram->in sram[2073]->out sram[2073]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2073]->out) 0
.nodeset V(sram[2073]->outb) vsp
Xmux_1level_tapbuf_size2[402] grid[1][2]_pin[0][2][11] chany[1][1]_in[82] chanx[1][1]_out[85] sram[2074]->outb sram[2074]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[402], level=1, select_path_id=0. *****
*****1*****
Xsram[2074] sram->in sram[2074]->out sram[2074]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2074]->out) 0
.nodeset V(sram[2074]->outb) vsp
Xmux_1level_tapbuf_size2[403] grid[1][2]_pin[0][2][11] chany[1][1]_in[84] chanx[1][1]_out[87] sram[2075]->outb sram[2075]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[403], level=1, select_path_id=0. *****
*****1*****
Xsram[2075] sram->in sram[2075]->out sram[2075]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2075]->out) 0
.nodeset V(sram[2075]->outb) vsp
Xmux_1level_tapbuf_size2[404] grid[1][2]_pin[0][2][11] chany[1][1]_in[86] chanx[1][1]_out[89] sram[2076]->outb sram[2076]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[404], level=1, select_path_id=0. *****
*****1*****
Xsram[2076] sram->in sram[2076]->out sram[2076]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2076]->out) 0
.nodeset V(sram[2076]->outb) vsp
Xmux_1level_tapbuf_size2[405] grid[1][2]_pin[0][2][13] chany[1][1]_in[88] chanx[1][1]_out[91] sram[2077]->outb sram[2077]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[405], level=1, select_path_id=0. *****
*****1*****
Xsram[2077] sram->in sram[2077]->out sram[2077]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2077]->out) 0
.nodeset V(sram[2077]->outb) vsp
Xmux_1level_tapbuf_size2[406] grid[1][2]_pin[0][2][13] chany[1][1]_in[90] chanx[1][1]_out[93] sram[2078]->outb sram[2078]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[406], level=1, select_path_id=0. *****
*****1*****
Xsram[2078] sram->in sram[2078]->out sram[2078]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2078]->out) 0
.nodeset V(sram[2078]->outb) vsp
Xmux_1level_tapbuf_size2[407] grid[1][2]_pin[0][2][13] chany[1][1]_in[92] chanx[1][1]_out[95] sram[2079]->outb sram[2079]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[407], level=1, select_path_id=0. *****
*****1*****
Xsram[2079] sram->in sram[2079]->out sram[2079]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2079]->out) 0
.nodeset V(sram[2079]->outb) vsp
Xmux_1level_tapbuf_size2[408] grid[1][2]_pin[0][2][13] chany[1][1]_in[94] chanx[1][1]_out[97] sram[2080]->outb sram[2080]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[408], level=1, select_path_id=0. *****
*****1*****
Xsram[2080] sram->in sram[2080]->out sram[2080]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2080]->out) 0
.nodeset V(sram[2080]->outb) vsp
Xmux_1level_tapbuf_size2[409] grid[1][2]_pin[0][2][13] chany[1][1]_in[96] chanx[1][1]_out[99] sram[2081]->outb sram[2081]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[409], level=1, select_path_id=0. *****
*****1*****
Xsram[2081] sram->in sram[2081]->out sram[2081]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[2081]->out) 0
.nodeset V(sram[2081]->outb) vsp
.eom
