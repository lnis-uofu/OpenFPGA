// Benchmark "TOP" written by ABC on Tue Mar  5 10:04:28 2019

module s38417 ( clock, 
    Pg3234, Pg3233, Pg3232, Pg3231, Pg3230, Pg3229, Pg3228, Pg3227, Pg3226,
    Pg3225, Pg3224, Pg3223, Pg3222, Pg3221, Pg3220, Pg3219, Pg3218, Pg3217,
    Pg3216, Pg3215, Pg3214, Pg3213, Pg3212, Pg2637, Pg1943, Pg1249, Pg563,
    Pg51,
    Pg27380, Pg26149, Pg26135, Pg26104, Pg25489, Pg25442, Pg25435, Pg25420,
    Pg24734, Pg16496, Pg16437, Pg16399, Pg16355, Pg16297, Pg8275, Pg8274,
    Pg8273, Pg8272, Pg8271, Pg8270, Pg8269, Pg8268, Pg8267, Pg8266, Pg8265,
    Pg8264, Pg8263, Pg8262, Pg8261, Pg8260, Pg8259, Pg8258, Pg8251, Pg8249,
    Pg8175, Pg8167, Pg8106, Pg8096, Pg8087, Pg8082, Pg8030, Pg8023, Pg8021,
    Pg8012, Pg8007, Pg7961, Pg7956, Pg7909, Pg7519, Pg7487, Pg7425, Pg7390,
    Pg7357, Pg7334, Pg7302, Pg7264, Pg7229, Pg7194, Pg7161, Pg7084, Pg7052,
    Pg7014, Pg6979, Pg6944, Pg6911, Pg6895, Pg6837, Pg6782, Pg6750, Pg6712,
    Pg6677, Pg6642, Pg6573, Pg6518, Pg6485, Pg6447, Pg6442, Pg6368, Pg6313,
    Pg6231, Pg6225, Pg5796, Pg5747, Pg5738, Pg5695, Pg5686, Pg5657, Pg5648,
    Pg5637, Pg5629, Pg5612, Pg5595, Pg5555, Pg5549, Pg5511, Pg5472, Pg5437,
    Pg5388, Pg4590, Pg4450, Pg4323, Pg4321, Pg4200, Pg4090, Pg4088, Pg3993  );
  input  Pg3234, Pg3233, Pg3232, Pg3231, Pg3230, Pg3229, Pg3228, Pg3227,
    Pg3226, Pg3225, Pg3224, Pg3223, Pg3222, Pg3221, Pg3220, Pg3219, Pg3218,
    Pg3217, Pg3216, Pg3215, Pg3214, Pg3213, Pg3212, Pg2637, Pg1943, Pg1249,
    Pg563, Pg51, clock;
  output Pg27380, Pg26149, Pg26135, Pg26104, Pg25489, Pg25442, Pg25435,
    Pg25420, Pg24734, Pg16496, Pg16437, Pg16399, Pg16355, Pg16297, Pg8275,
    Pg8274, Pg8273, Pg8272, Pg8271, Pg8270, Pg8269, Pg8268, Pg8267, Pg8266,
    Pg8265, Pg8264, Pg8263, Pg8262, Pg8261, Pg8260, Pg8259, Pg8258, Pg8251,
    Pg8249, Pg8175, Pg8167, Pg8106, Pg8096, Pg8087, Pg8082, Pg8030, Pg8023,
    Pg8021, Pg8012, Pg8007, Pg7961, Pg7956, Pg7909, Pg7519, Pg7487, Pg7425,
    Pg7390, Pg7357, Pg7334, Pg7302, Pg7264, Pg7229, Pg7194, Pg7161, Pg7084,
    Pg7052, Pg7014, Pg6979, Pg6944, Pg6911, Pg6895, Pg6837, Pg6782, Pg6750,
    Pg6712, Pg6677, Pg6642, Pg6573, Pg6518, Pg6485, Pg6447, Pg6442, Pg6368,
    Pg6313, Pg6231, Pg6225, Pg5796, Pg5747, Pg5738, Pg5695, Pg5686, Pg5657,
    Pg5648, Pg5637, Pg5629, Pg5612, Pg5595, Pg5555, Pg5549, Pg5511, Pg5472,
    Pg5437, Pg5388, Pg4590, Pg4450, Pg4323, Pg4321, Pg4200, Pg4090, Pg4088,
    Pg3993;
  reg Pg8021, Ng2817, Ng2933, Ng13457, Ng2883, Ng2888, Ng2896, Ng2892,
    Ng2903, Ng2900, Ng2908, Ng2912, Ng2917, Ng2924, Ng2920, Ng2984, Ng2985,
    Ng2929, Ng2879, Ng2934, Ng2935, Ng2938, Ng2941, Ng2944, Ng2947, Ng2953,
    Ng2956, Ng2959, Ng2962, Ng2963, Ng2966, Ng2969, Ng2972, Ng2975, Ng2978,
    Ng2981, Ng2874, Ng1506, Ng1501, Ng1496, Ng1491, Ng1486, Ng1481, Ng1476,
    Ng1471, Ng13439, Pg8251, Ng813, Pg4090, Ng809, Pg4323, Ng805, Pg4590,
    Ng801, Pg6225, Ng797, Pg6442, Ng793, Pg6895, Ng789, Pg7334, Ng785,
    Pg7519, Ng13423, Pg8249, Ng125, Pg4088, Ng121, Pg4321, Ng117, Pg8023,
    Ng113, Pg8175, Ng109, Pg3993, Ng105, Pg4200, Ng101, Pg4450, Ng97,
    Pg8096, Ng13407, Ng2200, Ng2195, Ng2190, Ng2185, Ng2180, Ng2175,
    Ng2170, Ng2165, Ng13455, Ng3210, Ng3211, Ng3084, Ng3085, Ng3086,
    Ng3087, Ng3091, Ng3092, Ng3093, Ng3094, Ng3095, Ng3096, Ng3097, Ng3098,
    Ng3099, Ng3100, Ng3101, Ng3102, Ng3103, Ng3104, Ng3105, Ng3106, Ng3107,
    Ng3108, Ng3155, Ng3158, Ng3161, Ng3164, Ng3167, Ng3170, Ng3173, Ng3176,
    Ng3179, Ng3182, Ng3185, Ng3088, Ng3191, Ng3128, Ng3126, Ng3125, Ng3123,
    Ng3120, Ng3110, Ng3139, Ng3135, Ng3147, Ng185, Ng130, Ng131, Ng129,
    Ng133, Ng134, Ng132, Ng142, Ng143, Ng141, Ng145, Ng146, Ng144, Ng148,
    Ng149, Ng147, Ng151, Ng152, Ng150, Ng154, Ng155, Ng153, Ng157, Ng158,
    Ng156, Ng160, Ng161, Ng159, Ng163, Ng164, Ng162, Ng169, Ng170, Ng168,
    Ng172, Ng173, Ng171, Ng175, Ng176, Ng174, Ng178, Ng179, Ng177, Ng186,
    Ng189, Ng192, Ng231, Ng234, Ng237, Ng195, Ng198, Ng201, Ng240, Ng243,
    Ng246, Ng204, Ng207, Ng210, Ng249, Ng252, Ng255, Ng213, Ng216, Ng219,
    Ng258, Ng261, Ng264, Ng222, Ng225, Ng228, Ng267, Ng270, Ng273, Ng92,
    Ng88, Ng83, Ng79, Ng74, Ng70, Ng65, Ng61, Ng56, Ng52, Ng11497, Ng11498,
    Ng11499, Ng11500, Ng11501, Ng11502, Ng11503, Ng11504, Ng11505, Ng11506,
    Ng11507, Ng11508, Ng408, Ng411, Ng414, Ng417, Ng420, Ng423, Ng427,
    Ng428, Ng426, Ng429, Ng432, Ng435, Ng438, Ng441, Ng444, Ng448, Ng449,
    Ng447, Ng312, Ng313, Ng314, Ng315, Ng316, Ng317, Ng318, Ng319, Ng320,
    Ng322, Ng323, Ng321, Ng403, Ng404, Ng402, Ng450, Ng451, Ng452, Ng453,
    Ng454, Ng279, Ng280, Ng281, Ng282, Ng283, Ng284, Ng285, Ng286, Ng287,
    Ng288, Ng289, Ng290, Ng291, Ng299, Ng305, Ng298, Ng342, Ng349, Ng350,
    Ng351, Ng352, Ng353, Ng357, Ng364, Ng365, Ng366, Ng367, Ng368, Ng372,
    Ng379, Ng380, Ng381, Ng382, Ng383, Ng387, Ng394, Ng395, Ng396, Ng397,
    Ng324, Ng554, Ng557, Ng510, Ng513, Ng523, Ng524, Ng564, Ng569, Ng570,
    Ng571, Ng572, Ng573, Ng574, Ng565, Ng566, Ng567, Ng568, Ng489, Ng486,
    Ng487, Ng488, Ng11512, Ng11515, Ng11516, Ng477, Ng478, Ng479, Ng480,
    Ng484, Ng464, Ng11517, Ng11513, Ng11514, Ng528, Ng535, Ng542, Ng543,
    Ng544, Ng548, Ng549, Ng8284, Ng558, Ng559, Ng576, Ng577, Ng575, Ng579,
    Ng580, Ng578, Ng582, Ng583, Ng581, Ng585, Ng586, Ng584, Ng587, Ng590,
    Ng593, Ng596, Ng599, Ng602, Ng614, Ng617, Ng620, Ng605, Ng608, Ng611,
    Ng490, Ng493, Ng496, Ng506, Ng507, Pg16297, Ng525, Ng529, Ng530, Ng531,
    Ng532, Ng533, Ng534, Ng536, Ng537, Ng538, Ng541, Ng630, Ng659, Ng640,
    Ng633, Ng653, Ng646, Ng660, Ng672, Ng666, Ng679, Ng686, Ng692, Ng699,
    Ng700, Ng698, Ng702, Ng703, Ng701, Ng705, Ng706, Ng704, Ng708, Ng709,
    Ng707, Ng711, Ng712, Ng710, Ng714, Ng715, Ng713, Ng717, Ng718, Ng716,
    Ng720, Ng721, Ng719, Ng723, Ng724, Ng722, Ng726, Ng727, Ng725, Ng729,
    Ng730, Ng728, Ng732, Ng733, Ng731, Ng735, Ng736, Ng734, Ng738, Ng739,
    Ng737, \[1612] , \[1594] , Ng853, Ng818, Ng819, Ng817, Ng821, Ng822,
    Ng820, Ng830, Ng831, Ng829, Ng833, Ng834, Ng832, Ng836, Ng837, Ng835,
    Ng839, Ng840, Ng838, Ng842, Ng843, Ng841, Ng845, Ng846, Ng844, Ng848,
    Ng849, Ng847, Ng851, Ng852, Ng850, Ng857, Ng858, Ng856, Ng860, Ng861,
    Ng859, Ng863, Ng864, Ng862, Ng866, Ng867, Ng865, Ng873, Ng876, Ng879,
    Ng918, Ng921, Ng924, Ng882, Ng885, Ng888, Ng927, Ng930, Ng933, Ng891,
    Ng894, Ng897, Ng936, Ng939, Ng942, Ng900, Ng903, Ng906, Ng945, Ng948,
    Ng951, Ng909, Ng912, Ng915, Ng954, Ng957, Ng960, Ng780, Ng776, Ng771,
    Ng767, Ng762, Ng758, Ng753, Ng749, Ng744, Ng740, Ng11524, Ng11525,
    Ng11526, Ng11527, Ng11528, Ng11529, Ng11530, Ng11531, Ng11532, Ng11533,
    Ng11534, Ng11535, Ng1095, Ng1098, Ng1101, Ng1104, Ng1107, Ng1110,
    Ng1114, Ng1115, Ng1113, Ng1116, Ng1119, Ng1122, Ng1125, Ng1128, Ng1131,
    Ng1135, Ng1136, Ng1134, Ng999, Ng1000, Ng1001, Ng1002, Ng1003, Ng1004,
    Ng1005, Ng1006, Ng1007, Ng1009, Ng1010, Ng1008, Ng1090, Ng1091, Ng1089,
    Ng1137, Ng1138, Ng1139, Ng1140, Ng1141, Ng966, Ng967, Ng968, Ng969,
    Ng970, Ng971, Ng972, Ng973, Ng974, Ng975, Ng976, Ng977, Ng978, Ng986,
    Ng992, Ng985, Ng1029, Ng1036, Ng1037, Ng1038, Ng1039, Ng1040, Ng1044,
    Ng1051, Ng1052, Ng1053, Ng1054, Ng1055, Ng1059, Ng1066, Ng1067, Ng1068,
    Ng1069, Ng1070, Ng1074, Ng1081, Ng1082, Ng1083, Ng1084, Ng1011, Ng1240,
    Ng1243, Ng1196, Ng1199, Ng1209, Ng1210, Ng1250, Ng1255, Ng1256, Ng1257,
    Ng1258, Ng1259, Ng1260, Ng1251, Ng1252, Ng1253, Ng1254, Ng1176, Ng1173,
    Ng1174, Ng1175, Ng11539, Ng11542, Ng11543, Ng1164, Ng1165, Ng1166,
    Ng1167, Ng1171, Ng1151, Ng11544, Ng11540, Ng11541, Ng1214, Ng1221,
    Ng1228, Ng1229, Ng1230, Ng1234, Ng1235, Ng8293, Ng1244, Ng1245, Ng1262,
    Ng1263, Ng1261, Ng1265, Ng1266, Ng1264, Ng1268, Ng1269, Ng1267, Ng1271,
    Ng1272, Ng1270, Ng1273, Ng1276, Ng1279, Ng1282, Ng1285, Ng1288, Ng1300,
    Ng1303, Ng1306, Ng1291, Ng1294, Ng1297, Ng1177, Ng1180, Ng1183, Ng1192,
    Ng1193, Pg16355, Ng1211, Ng1215, Ng1216, Ng1217, Ng1218, Ng1219,
    Ng1220, Ng1222, Ng1223, Ng1224, Ng1227, \[1605] , \[1603] , Ng1315,
    Ng1316, Ng1345, Ng1326, Ng1319, Ng1339, Ng1332, Ng1346, Ng1358, Ng1352,
    Ng1365, Ng1372, Ng1378, Ng1385, Ng1386, Ng1384, Ng1388, Ng1389, Ng1387,
    Ng1391, Ng1392, Ng1390, Ng1394, Ng1395, Ng1393, Ng1397, Ng1398, Ng1396,
    Ng1400, Ng1401, Ng1399, Ng1403, Ng1404, Ng1402, Ng1406, Ng1407, Ng1405,
    Ng1409, Ng1410, Ng1408, Ng1412, Ng1413, Ng1411, Ng1415, Ng1416, Ng1414,
    Ng1418, Ng1419, Ng1417, Ng1421, Ng1422, Ng1420, Ng1424, Ng1425, Ng1423,
    Ng1512, Ng1513, Ng1511, Ng1515, Ng1516, Ng1514, Ng1524, Ng1525, Ng1523,
    Ng1527, Ng1528, Ng1526, Ng1530, Ng1531, Ng1529, Ng1533, Ng1534, Ng1532,
    Ng1536, Ng1537, Ng1535, Ng1539, Ng1540, Ng1538, Ng1542, Ng1543, Ng1541,
    Ng1545, Ng1546, Ng1544, Ng1551, Ng1552, Ng1550, Ng1554, Ng1555, Ng1553,
    Ng1557, Ng1558, Ng1556, Ng1560, Ng1561, Ng1559, Ng1567, Ng1570, Ng1573,
    Ng1612, Ng1615, Ng1618, Ng1576, Ng1579, Ng1582, Ng1621, Ng1624, Ng1627,
    Ng1585, Ng1588, Ng1591, Ng1630, Ng1633, Ng1636, Ng1594, Ng1597, Ng1600,
    Ng1639, Ng1642, Ng1645, Ng1603, Ng1606, Ng1609, Ng1648, Ng1651, Ng1654,
    Ng1466, Ng1462, Ng1457, Ng1453, Ng1448, Ng1444, Ng1439, Ng1435, Ng1430,
    Ng1426, Ng11551, Ng11552, Ng11553, Ng11554, Ng11555, Ng11556, Ng11557,
    Ng11558, Ng11559, Ng11560, Ng11561, Ng11562, Ng1789, Ng1792, Ng1795,
    Ng1798, Ng1801, Ng1804, Ng1808, Ng1809, Ng1807, Ng1810, Ng1813, Ng1816,
    Ng1819, Ng1822, Ng1825, Ng1829, Ng1830, Ng1828, Ng1693, Ng1694, Ng1695,
    Ng1696, Ng1697, Ng1698, Ng1699, Ng1700, Ng1701, Ng1703, Ng1704, Ng1702,
    Ng1784, Ng1785, Ng1783, Ng1831, Ng1832, Ng1833, Ng1834, Ng1835, Ng1660,
    Ng1661, Ng1662, Ng1663, Ng1664, Ng1665, Ng1666, Ng1667, Ng1668, Ng1669,
    Ng1670, Ng1671, Ng1672, Ng1680, Ng1686, Ng1679, Ng1723, Ng1730, Ng1731,
    Ng1732, Ng1733, Ng1734, Ng1738, Ng1745, Ng1746, Ng1747, Ng1748, Ng1749,
    Ng1753, Ng1760, Ng1761, Ng1762, Ng1763, Ng1764, Ng1768, Ng1775, Ng1776,
    Ng1777, Ng1778, Ng1705, Ng1934, Ng1937, Ng1890, Ng1893, Ng1903, Ng1904,
    Ng1944, Ng1949, Ng1950, Ng1951, Ng1952, Ng1953, Ng1954, Ng1945, Ng1946,
    Ng1947, Ng1948, Ng1870, Ng1867, Ng1868, Ng1869, Ng11566, Ng11569,
    Ng11570, Ng1858, Ng1859, Ng1860, Ng1861, Ng1865, Ng1845, Ng11571,
    Ng11567, Ng11568, Ng1908, Ng1915, Ng1922, Ng1923, Ng1924, Ng1928,
    Ng1929, Ng8302, Ng1938, Ng1939, Ng1956, Ng1957, Ng1955, Ng1959, Ng1960,
    Ng1958, Ng1962, Ng1963, Ng1961, Ng1965, Ng1966, Ng1964, Ng1967, Ng1970,
    Ng1973, Ng1976, Ng1979, Ng1982, Ng1994, Ng1997, Ng2000, Ng1985, Ng1988,
    Ng1991, Ng1871, Ng1874, Ng1877, Ng1886, Ng1887, Pg16399, Ng1905,
    Ng1909, Ng1910, Ng1911, Ng1912, Ng1913, Ng1914, Ng1916, Ng1917, Ng1918,
    Ng1921, Ng2010, Ng2039, Ng2020, Ng2013, Ng2033, Ng2026, Ng2040, Ng2052,
    Ng2046, Ng2059, Ng2066, Ng2072, Ng2079, Ng2080, Ng2078, Ng2082, Ng2083,
    Ng2081, Ng2085, Ng2086, Ng2084, Ng2088, Ng2089, Ng2087, Ng2091, Ng2092,
    Ng2090, Ng2094, Ng2095, Ng2093, Ng2097, Ng2098, Ng2096, Ng2100, Ng2101,
    Ng2099, Ng2103, Ng2104, Ng2102, Ng2106, Ng2107, Ng2105, Ng2109, Ng2110,
    Ng2108, Ng2112, Ng2113, Ng2111, Ng2115, Ng2116, Ng2114, Ng2118, Ng2119,
    Ng2117, Ng2206, Ng2207, Ng2205, Ng2209, Ng2210, Ng2208, Ng2218, Ng2219,
    Ng2217, Ng2221, Ng2222, Ng2220, Ng2224, Ng2225, Ng2223, Ng2227, Ng2228,
    Ng2226, Ng2230, Ng2231, Ng2229, Ng2233, Ng2234, Ng2232, Ng2236, Ng2237,
    Ng2235, Ng2239, Ng2240, Ng2238, Ng2245, Ng2246, Ng2244, Ng2248, Ng2249,
    Ng2247, Ng2251, Ng2252, Ng2250, Ng2254, Ng2255, Ng2253, Ng2261, Ng2264,
    Ng2267, Ng2306, Ng2309, Ng2312, Ng2270, Ng2273, Ng2276, Ng2315, Ng2318,
    Ng2321, Ng2279, Ng2282, Ng2285, Ng2324, Ng2327, Ng2330, Ng2288, Ng2291,
    Ng2294, Ng2333, Ng2336, Ng2339, Ng2297, Ng2300, Ng2303, Ng2342, Ng2345,
    Ng2348, Ng2160, Ng2156, Ng2151, Ng2147, Ng2142, Ng2138, Ng2133, Ng2129,
    Ng2124, Ng2120, Ng2256, \[1609] , Ng2257, Ng11578, Ng11579, Ng11580,
    Ng11581, Ng11582, Ng11583, Ng11584, Ng11585, Ng11586, Ng11587, Ng11588,
    Ng11589, Ng2483, Ng2486, Ng2489, Ng2492, Ng2495, Ng2498, Ng2502,
    Ng2503, Ng2501, Ng2504, Ng2507, Ng2510, Ng2513, Ng2516, Ng2519, Ng2523,
    Ng2524, Ng2522, Ng2387, Ng2388, Ng2389, Ng2390, Ng2391, Ng2392, Ng2393,
    Ng2394, Ng2395, Ng2397, Ng2398, Ng2396, Ng2478, Ng2479, Ng2477, Ng2525,
    Ng2526, Ng2527, Ng2528, Ng2529, Ng2354, Ng2355, Ng2356, Ng2357, Ng2358,
    Ng2359, Ng2360, Ng2361, Ng2362, Ng2363, Ng2364, Ng2365, Ng2366, Ng2374,
    Ng2380, Ng2373, Ng2417, Ng2424, Ng2425, Ng2426, Ng2427, Ng2428, Ng2432,
    Ng2439, Ng2440, Ng2441, Ng2442, Ng2443, Ng2447, Ng2454, Ng2455, Ng2456,
    Ng2457, Ng2458, Ng2462, Ng2469, Ng2470, Ng2471, Ng2472, Ng2399, Ng2628,
    Ng2631, Ng2584, Ng2587, Ng2597, Ng2598, Ng2638, Ng2643, Ng2644, Ng2645,
    Ng2646, Ng2647, Ng2648, Ng2639, Ng2640, Ng2641, Ng2642, Ng2564, Ng2561,
    Ng2562, Ng2563, Ng11593, Ng11596, Ng11597, Ng2552, Ng2553, Ng2554,
    Ng2555, Ng2559, Ng2539, Ng11598, Ng11594, Ng11595, Ng2602, Ng2609,
    Ng2616, Ng2617, Ng2618, Ng2622, Ng2623, Ng8311, Ng2632, Ng2633, Ng2650,
    Ng2651, Ng2649, Ng2653, Ng2654, Ng2652, Ng2656, Ng2657, Ng2655, Ng2659,
    Ng2660, Ng2658, Ng2661, Ng2664, Ng2667, Ng2670, Ng2673, Ng2676, Ng2688,
    Ng2691, Ng2694, Ng2679, Ng2682, Ng2685, Ng2565, Ng2568, Ng2571, Ng2580,
    Ng2581, Pg16437, Ng2599, Ng2603, Ng2604, Ng2605, Ng2606, Ng2607,
    Ng2608, Ng2610, Ng2611, Ng2612, Ng2615, Ng2704, Ng2733, Ng2714, Ng2707,
    Ng2727, Ng2720, Ng2734, Ng2746, Ng2740, Ng2753, Ng2760, Ng2766, Ng2773,
    Ng2774, Ng2772, Ng2776, Ng2777, Ng2775, Ng2779, Ng2780, Ng2778, Ng2782,
    Ng2783, Ng2781, Ng2785, Ng2786, Ng2784, Ng2788, Ng2789, Ng2787, Ng2791,
    Ng2792, Ng2790, Ng2794, Ng2795, Ng2793, Ng2797, Ng2798, Ng2796, Ng2800,
    Ng2801, Ng2799, Ng2803, Ng2804, Ng2802, Ng2806, Ng2807, Ng2805, Ng2809,
    Ng2810, Ng2808, Ng2812, Ng2813, Ng2811, Ng3054, Ng3079, Ng13475,
    Ng3043, Ng3044, Ng3045, Ng3046, Ng3047, Ng3048, Ng3049, Ng3050, Ng3051,
    Ng3052, Ng3053, Ng3055, Ng3056, Ng3057, Ng3058, Ng3059, Ng3060, Ng3061,
    Ng3062, Ng3063, Ng3064, Ng3065, Ng3066, Ng3067, Ng3068, Ng3069, Ng3070,
    Ng3071, Ng3072, Ng3073, Ng3074, Ng3075, Ng3076, Ng3077, Ng3078, Ng2997,
    Ng2993, Ng2998, Ng3006, Ng3002, Ng3013, Ng3010, Ng3024, Ng3018, Ng3028,
    Ng3036, Ng3032, Pg5388, Ng2986, Ng2987, Pg8275, Pg8274, Pg8273, Pg8272,
    Pg8268, Pg8269, Pg8270, Pg8271, Ng3083, Pg8267, Ng2992, Pg8266, Pg8265,
    Pg8264, Pg8262, Pg8263, Pg8260, Pg8261, Pg8259, Ng2990, Ng2991, Pg8258;
  wire n4530, n4531_1, n4532, n4533, n4534, n4535, n4536_1, n4537, n4538,
    n4539, n4540, n4541_1, n4542, n4543, n4544, n4545, n4546_1, n4547,
    n4548, n4549, n4550_1, n4551, n4552, n4553, n4554, n4555_1, n4556,
    n4557, n4558, n4559_1, n4560, n4561, n4562, n4563, n4564_1, n4565,
    n4566, n4567, n4568_1, n4569, n4570, n4571, n4572, n4573_1, n4574,
    n4575, n4576, n4577_1, n4578, n4579, n4580, n4581, n4582_1, n4583,
    n4584, n4585, n4586_1, n4588, n4590, n4591_1, n4592, n4593, n4594,
    n4596, n4598, n4600_1, n4601, n4602, n4603, n4604_1, n4606, n4608,
    n4610, n4612, n4613_1, n4614, n4615, n4616, n4618, n4620, n4622, n4624,
    n4625, n4626_1, n4628, n4630, n4632, n4633, n4634, n4636_1, n4638,
    n4639, n4640_1, n4642, n4643, n4644, n4646, n4647, n4648_1, n4649,
    n4650, n4651, n4652_1, n4653, n4654, n4655, n4656_1, n4657, n4658,
    n4659, n4660_1, n4661, n4662, n4663, n4664_1, n4665, n4666, n4667,
    n4668_1, n4669, n4670, n4671, n4672_1, n4673, n4674, n4675, n4676_1,
    n4677, n4678, n4679, n4680_1, n4681, n4682, n4683, n4684_1, n4685,
    n4686, n4687, n4688_1, n4689, n4690, n4691, n4692_1, n4693, n4694,
    n4695, n4696_1, n4697, n4698, n4699, n4700_1, n4701, n4702, n4703,
    n4704_1, n4705, n4706, n4707, n4708_1, n4709, n4710, n4711, n4712_1,
    n4713, n4714, n4715, n4716_1, n4717, n4718, n4719, n4720_1, n4721,
    n4722, n4723, n4724_1, n4725, n4726, n4727, n4728_1, n4729, n4730,
    n4731, n4732_1, n4733, n4734, n4735, n4736, n4737_1, n4738, n4739,
    n4740, n4741, n4742_1, n4743, n4744, n4745, n4746, n4747_1, n4748,
    n4749, n4750, n4751, n4752_1, n4753, n4754, n4755, n4756_1, n4757,
    n4758, n4759, n4760_1, n4761, n4762, n4763, n4764, n4765_1, n4766,
    n4767, n4768, n4769_1, n4770, n4771, n4772, n4773, n4774_1, n4775,
    n4776, n4777, n4778_1, n4779, n4780, n4781, n4782, n4783_1, n4784,
    n4785, n4786, n4787_1, n4788, n4789, n4790, n4791, n4792_1, n4793,
    n4794, n4795, n4796_1, n4797, n4798, n4799, n4800, n4801_1, n4802,
    n4803, n4804, n4805_1, n4806, n4807, n4808, n4809, n4810_1, n4811,
    n4812, n4813, n4814_1, n4815, n4816, n4817, n4818, n4819_1, n4820,
    n4821, n4822, n4823, n4824_1, n4825, n4826, n4827, n4828, n4829_1,
    n4830, n4831, n4832, n4833, n4834_1, n4835, n4836, n4837, n4838_1,
    n4839, n4840, n4841, n4842_1, n4843, n4844, n4845, n4846_1, n4847,
    n4848, n4849, n4850, n4851_1, n4852, n4853, n4854, n4855, n4856_1,
    n4857, n4858, n4859, n4860, n4861_1, n4862, n4863, n4864, n4865,
    n4866_1, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
    n4876_1, n4877, n4878, n4879, n4880_1, n4881, n4882, n4883, n4884_1,
    n4885, n4886, n4887, n4888_1, n4889, n4890, n4891, n4892_1, n4893,
    n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901_1, n4902, n4903,
    n4904, n4905, n4906, n4907, n4908, n4909, n4910_1, n4911, n4912, n4913,
    n4914, n4915_1, n4916, n4917, n4918, n4919_1, n4920, n4921, n4922,
    n4923, n4924_1, n4925, n4926, n4927, n4928_1, n4929, n4930, n4931,
    n4932, n4933_1, n4934, n4935, n4936, n4937, n4938_1, n4939, n4940,
    n4941, n4942, n4943_1, n4944, n4945, n4946, n4947, n4948_1, n4949,
    n4950, n4951, n4952, n4953_1, n4954, n4955, n4956, n4957, n4958_1,
    n4959, n4960, n4961, n4962, n4963_1, n4964, n4965, n4966, n4967,
    n4968_1, n4969, n4970, n4971, n4972, n4973_1, n4974, n4975, n4976,
    n4977, n4978_1, n4979, n4980, n4981, n4982, n4983_1, n4984, n4985,
    n4986, n4987, n4988_1, n4989, n4990, n4991, n4992, n4993_1, n4994,
    n4995, n4996, n4997, n4998_1, n4999, n5000, n5001, n5002, n5003_1,
    n5004, n5005, n5006, n5007, n5008_1, n5009, n5010, n5011, n5012,
    n5013_1, n5014, n5015, n5016, n5017, n5018_1, n5019, n5020, n5021,
    n5022, n5023_1, n5024, n5025, n5026, n5027, n5028_1, n5029, n5030,
    n5031, n5032, n5033_1, n5034, n5035, n5036, n5037, n5038_1, n5039,
    n5040, n5041, n5042, n5043_1, n5044, n5045, n5046, n5047, n5049, n5050,
    n5051, n5052, n5053_1, n5054, n5055, n5056, n5057, n5058_1, n5059,
    n5060, n5061, n5062, n5063_1, n5064, n5065, n5066, n5067_1, n5068,
    n5069, n5070, n5071, n5072_1, n5073, n5074, n5075, n5076, n5077_1,
    n5078, n5079, n5080_1, n5081, n5082, n5083, n5084, n5087, n5089, n5091,
    n5093, n5097, n5099, n5101, n5103, n5105_1, n5106, n5108, n5109, n5111,
    n5112, n5114, n5115_1, n5117, n5118, n5122, n5124, n5126, n5127, n5128,
    n5129, n5131, n5132, n5133, n5135_1, n5136, n5137, n5138, n5139,
    n5140_1, n5142, n5144, n5145_1, n5147, n5149, n5151, n5153, n5154,
    n5156, n5158, n5160_1, n5161, n5163, n5164, n5165_1, n5166, n5168,
    n5170_1, n5171, n5173, n5174, n5175_1, n5176, n5178, n5180_1, n5181,
    n5183, n5184, n5185_1, n5186, n5188, n5190_1, n5191, n5192, n5193,
    n5196, n5198, n5200_1, n5202, n5204, n5206, n5208, n5210_1, n5213,
    n5215_1, n5217, n5219, n5221, n5223, n5225_1, n5227, n5229, n5230_1,
    n5232, n5234, n5236, n5239, n5241, n5243, n5245_1, n5247, n5249, n5251,
    n5253, n5255_1, n5257, n5259, n5261, n5263, n5265_1, n5267, n5269,
    n5271, n5273, n5275_1, n5277, n5279, n5281, n5284, n5286, n5289, n5291,
    n5293, n5295_1, n5297, n5299, n5301, n5303, n5305_1, n5307, n5309,
    n5311, n5312, n5313, n5314, n5315_1, n5316, n5317, n5318, n5319,
    n5320_1, n5321, n5322, n5323, n5325_1, n5327, n5329, n5331, n5333,
    n5335_1, n5337, n5339, n5340_1, n5342, n5344, n5345_1, n5347, n5349,
    n5351, n5352, n5354, n5356, n5358, n5359, n5361, n5363, n5365_1, n5367,
    n5369, n5371, n5373, n5375_1, n5377, n5379, n5381, n5383, n5385_1,
    n5387, n5389, n5391, n5392, n5394, n5396, n5397, n5399, n5401, n5403,
    n5404, n5406, n5408, n5410_1, n5411, n5413, n5415_1, n5417, n5419,
    n5421, n5423, n5425_1, n5427, n5429, n5431, n5433, n5435_1, n5436,
    n5437, n5438, n5439, n5440_1, n5441, n5442, n5443, n5444, n5445_1,
    n5446, n5447, n5448, n5449, n5450_1, n5451, n5452, n5453, n5454,
    n5455_1, n5456, n5457, n5458, n5459, n5460_1, n5461, n5462, n5463,
    n5464, n5465_1, n5466, n5467, n5468, n5469, n5470_1, n5471, n5472,
    n5473, n5474, n5475_1, n5476, n5477, n5478, n5479, n5480_1, n5481,
    n5482, n5483, n5484, n5485_1, n5486, n5487, n5488, n5489, n5490_1,
    n5491, n5492, n5493, n5494, n5495_1, n5496, n5497, n5498, n5499,
    n5500_1, n5501, n5502, n5503, n5504, n5505_1, n5506, n5507, n5508,
    n5509, n5510_1, n5511, n5512, n5513, n5514, n5515_1, n5516, n5517,
    n5518, n5519, n5520_1, n5521, n5522, n5523, n5524, n5525_1, n5526,
    n5527, n5528, n5529, n5530_1, n5531, n5532, n5533, n5534, n5535_1,
    n5536, n5537, n5538, n5539, n5540_1, n5541, n5542, n5543, n5544,
    n5545_1, n5546, n5547, n5548, n5549, n5550_1, n5551, n5552, n5553,
    n5554, n5555_1, n5556, n5557, n5558, n5559, n5560_1, n5561, n5562,
    n5563, n5564, n5565_1, n5566, n5567, n5568, n5569, n5570_1, n5571,
    n5572, n5573, n5574, n5575_1, n5576, n5577, n5578, n5579, n5580_1,
    n5581, n5582, n5583, n5584, n5585_1, n5586, n5587, n5588, n5589,
    n5590_1, n5591, n5592, n5593, n5594, n5595_1, n5596, n5597, n5598,
    n5599, n5600_1, n5601, n5602, n5603, n5604, n5605_1, n5606, n5607,
    n5608, n5609, n5610_1, n5611, n5612, n5613, n5614, n5615_1, n5616,
    n5617, n5618, n5619, n5620_1, n5621, n5622, n5623, n5624, n5625_1,
    n5626, n5627, n5628, n5629, n5630_1, n5631, n5632, n5633, n5634,
    n5635_1, n5636, n5637, n5638, n5639, n5640_1, n5641, n5642, n5643,
    n5644, n5645_1, n5646, n5647, n5648, n5649, n5650_1, n5651, n5652,
    n5653, n5654, n5655_1, n5656, n5657, n5658, n5659, n5660_1, n5661,
    n5662, n5663, n5664, n5665_1, n5666, n5667, n5668, n5669, n5670_1,
    n5671, n5672, n5677, n5679, n5681, n5683, n5685_1, n5687, n5689, n5691,
    n5693, n5695_1, n5697, n5699, n5701, n5703, n5705_1, n5707, n5709,
    n5711, n5713, n5715_1, n5717, n5719, n5721, n5723, n5725_1, n5727,
    n5729, n5731, n5733, n5735_1, n5737, n5739, n5741, n5743, n5745_1,
    n5747, n5817, n5818, n5819_1, n5820, n5821, n5822, n5823_1, n5824,
    n5825, n5826, n5827, n5828_1, n5829, n5830, n5831, n5832, n5833_1,
    n5834, n5835, n5836, n5837, n5838_1, n5839, n5840, n5841, n5842,
    n5843_1, n5844, n5845, n5846, n5847, n5848_1, n5849, n5850, n5851,
    n5852, n5853_1, n5854, n5855, n5856, n5857, n5858_1, n5859, n5860,
    n5861, n5862, n5863_1, n5864, n5865, n5866, n5867, n5868_1, n5869,
    n5870, n5871, n5872, n5873_1, n5874, n5875, n5876, n5877, n5878_1,
    n5879, n5880, n5881, n5882, n5883_1, n5884, n5885, n5886, n5887,
    n5888_1, n5889, n5890, n5891, n5892, n5893_1, n5894, n5895, n5896,
    n5897, n5898_1, n5899, n5900, n5901, n5902, n5903_1, n5904, n5905,
    n5906, n5907, n5908_1, n5909, n5910, n5911, n5912, n5913_1, n5914,
    n5915, n5916, n5917, n5918_1, n5919, n5920, n5921, n5922, n5923_1,
    n5924, n5925, n5926, n5927, n5928_1, n5929, n5930, n5931, n5932,
    n5933_1, n5934, n5935, n5936, n5937, n5938_1, n5939, n5940, n5941,
    n5942, n5943_1, n5944, n5945, n5946, n5947, n5948_1, n5949, n5950,
    n5951, n5952, n5953_1, n5954, n5955, n5956, n5957, n5958_1, n5959,
    n5960, n5961, n5962, n5963_1, n5964, n5965, n5966, n5967, n5968_1,
    n5969, n5970, n5971, n5972, n5973_1, n5974, n5975, n5976, n5977,
    n5978_1, n5979, n5980, n5981, n5982, n5983_1, n5984, n5985, n5986,
    n5987, n5988_1, n5989, n5990, n5991, n5992, n5993_1, n5994, n5995,
    n5996, n5997, n5998_1, n5999, n6000, n6001, n6002, n6003_1, n6004,
    n6005, n6006, n6007, n6008_1, n6009, n6010, n6011, n6012, n6013_1,
    n6014, n6015, n6016, n6017, n6018_1, n6019, n6020, n6021, n6022,
    n6023_1, n6024, n6025, n6026, n6027, n6028_1, n6029, n6030, n6031,
    n6032, n6033_1, n6034, n6035, n6036, n6037, n6038_1, n6039, n6040,
    n6041, n6042, n6043_1, n6044, n6045, n6046, n6047, n6048_1, n6049,
    n6050, n6051, n6052, n6053_1, n6054, n6055, n6056, n6057_1, n6058,
    n6059, n6060, n6061, n6062_1, n6063, n6064, n6065, n6066_1, n6067,
    n6068, n6069, n6070, n6071_1, n6072, n6073, n6074, n6075_1, n6076,
    n6077, n6078, n6079, n6080_1, n6081, n6082, n6083, n6084_1, n6085,
    n6086, n6087, n6088, n6089_1, n6090, n6091, n6092, n6093_1, n6094,
    n6095, n6096, n6097, n6098_1, n6099, n6100, n6101, n6102_1, n6103,
    n6104, n6105, n6106, n6107_1, n6108, n6109, n6110, n6111_1, n6112,
    n6113, n6114, n6115, n6116_1, n6117, n6118, n6119, n6120_1, n6121,
    n6122, n6123, n6124_1, n6125, n6126, n6127, n6128_1, n6129, n6130,
    n6131, n6132, n6133_1, n6134, n6135, n6136, n6137, n6138_1, n6139,
    n6140, n6141, n6142, n6143_1, n6144, n6145, n6146, n6147_1, n6148,
    n6149, n6150, n6151_1, n6152, n6153, n6154, n6155_1, n6156, n6157,
    n6158, n6159_1, n6160, n6161, n6162, n6163_1, n6164, n6165, n6166,
    n6167_1, n6168, n6169, n6170, n6171_1, n6172, n6173, n6174, n6175_1,
    n6176, n6177, n6178, n6179_1, n6180, n6181, n6182, n6183_1, n6184,
    n6185, n6186, n6187_1, n6188, n6189, n6190, n6191_1, n6192, n6193,
    n6194, n6195_1, n6196, n6197, n6198, n6199_1, n6200, n6201, n6202,
    n6203_1, n6204, n6205, n6206, n6207_1, n6208, n6209, n6210, n6211_1,
    n6212, n6213, n6214, n6215_1, n6216, n6217, n6218, n6219_1, n6221,
    n6222, n6223_1, n6225, n6226, n6227_1, n6229, n6230, n6231_1, n6233,
    n6234, n6235_1, n6236, n6237, n6238, n6239_1, n6240, n6241, n6242,
    n6243, n6244_1, n6245, n6246, n6247, n6248, n6249_1, n6250, n6251,
    n6252, n6253, n6254_1, n6255, n6256, n6257, n6258, n6259_1, n6260,
    n6261, n6262, n6263_1, n6264, n6265, n6266, n6267_1, n6268, n6269,
    n6270, n6271, n6272_1, n6273, n6274, n6275, n6276_1, n6277, n6278,
    n6279, n6280, n6281_1, n6282, n6283, n6285_1, n6286, n6287, n6288,
    n6289, n6290_1, n6291, n6292, n6293, n6294_1, n6295, n6296, n6297,
    n6298, n6299_1, n6300, n6301, n6302, n6303_1, n6304, n6305, n6306,
    n6307, n6308_1, n6309, n6310, n6311, n6312_1, n6313, n6314, n6315,
    n6316, n6317_1, n6318, n6319, n6320, n6321_1, n6322, n6323, n6324,
    n6325, n6326_1, n6327, n6328, n6329, n6330, n6331_1, n6332, n6333,
    n6334, n6335, n6336_1, n6337, n6338, n6339, n6340, n6341_1, n6342,
    n6343, n6344, n6345_1, n6346, n6347, n6348, n6349_1, n6350, n6351,
    n6352, n6353_1, n6354, n6355, n6356, n6357, n6358_1, n6359, n6360,
    n6361, n6362, n6363_1, n6364, n6365, n6366, n6367, n6368_1, n6369,
    n6370, n6371, n6372, n6373_1, n6374, n6375, n6376, n6377, n6378_1,
    n6379, n6380, n6381, n6382, n6383_1, n6384, n6385, n6386, n6387_1,
    n6388, n6389, n6390, n6391_1, n6392, n6393, n6394, n6395_1, n6396,
    n6397, n6398, n6399_1, n6400, n6401, n6402, n6403_1, n6404, n6405,
    n6406, n6407, n6408_1, n6409, n6410, n6411, n6412_1, n6413, n6414,
    n6415, n6416, n6417_1, n6418, n6419, n6420, n6421, n6422_1, n6423,
    n6424, n6425, n6426_1, n6427, n6428, n6429, n6430, n6431_1, n6432,
    n6433, n6434, n6435_1, n6436, n6437, n6438, n6439, n6440_1, n6441,
    n6442, n6443, n6444, n6445_1, n6446, n6447, n6448, n6449, n6450_1,
    n6451, n6452, n6453, n6454, n6455_1, n6456, n6457, n6458, n6459,
    n6460_1, n6461, n6462, n6463, n6464, n6465_1, n6466, n6467, n6468,
    n6469, n6470_1, n6471, n6472, n6473, n6474, n6476, n6478, n6479,
    n6480_1, n6481, n6482, n6483, n6484, n6485_1, n6486, n6487, n6488,
    n6489, n6490_1, n6491, n6492, n6493, n6494, n6495_1, n6496, n6497,
    n6498, n6499, n6500_1, n6501, n6502, n6503, n6504, n6505_1, n6506,
    n6507, n6508, n6509, n6510_1, n6511, n6512, n6513, n6514, n6515_1,
    n6516, n6517, n6518, n6520_1, n6521, n6522, n6523, n6524, n6526, n6527,
    n6528, n6529, n6530_1, n6531, n6532, n6533, n6534, n6535_1, n6536,
    n6537, n6538, n6539, n6540_1, n6541, n6542, n6543, n6544, n6545_1,
    n6546, n6547, n6548, n6549, n6550_1, n6551, n6552, n6553, n6554,
    n6555_1, n6556, n6557, n6558, n6559, n6560_1, n6561, n6562, n6563,
    n6564, n6565_1, n6566, n6567, n6568, n6569, n6570_1, n6571, n6572,
    n6573, n6574_1, n6575, n6576, n6577, n6578, n6579_1, n6580, n6581,
    n6582, n6583, n6584_1, n6585, n6586, n6587_1, n6588, n6589, n6591,
    n6595, n6597_1, n6599, n6600, n6601, n6602_1, n6603, n6604, n6605,
    n6606, n6607_1, n6608, n6610, n6612_1, n6614, n6615, n6616, n6617_1,
    n6618, n6619, n6621, n6623, n6625, n6626, n6627_1, n6629, n6631, n6633,
    n6635, n6637_1, n6639, n6641, n6643, n6645, n6647_1, n6649, n6651,
    n6653, n6655, n6657_1, n6659, n6661, n6663, n6664, n6665, n6667_1,
    n6669, n6671, n6673, n6675, n6677_1, n6679, n6681, n6683, n6685,
    n6687_1, n6689, n6691, n6693, n6695, n6697_1, n6699, n6701, n6702_1,
    n6703, n6705, n6707_1, n6709, n6711, n6713, n6715, n6717_1, n6719,
    n6721, n6723, n6725, n6727_1, n6729, n6731, n6733, n6735, n6737_1,
    n6739, n6740, n6741, n6743, n6745, n6747_1, n6749, n6751, n6753, n6755,
    n6757_1, n6759, n6761, n6763, n6765, n6767_1, n6769, n6771, n6773,
    n6775, n6777_1, n6779, n6781, n6783, n6785, n6787_1, n6789, n6791,
    n6793, n6795, n6796, n6798, n6800, n6802_1, n6804, n6806, n6808, n6809,
    n6811, n6813, n6815, n6816, n6818, n6820, n6822_1, n6823, n6825,
    n6827_1, n6829, n6830, n6832_1, n6834, n6836, n6838, n6840, n6842_1,
    n6843, n6845, n6847_1, n6849, n6850, n6852_1, n6854, n6856, n6857_1,
    n6859, n6861, n6863, n6864, n6866, n6868, n6870, n6872_1, n6874, n6876,
    n6877_1, n6879, n6881, n6883, n6884, n6886, n6888, n6890, n6891, n6893,
    n6895, n6897_1, n6898, n6900, n6902_1, n6904, n6906, n6908, n6910,
    n6911, n6913, n6915, n6917_1, n6918, n6920, n6922_1, n6924, n6925,
    n6927, n6929, n6932, n6934, n6936_1, n6938, n6940, n6942, n6944,
    n6946_1, n6948, n6949, n6950, n6951_1, n6952, n6953, n6955, n6957,
    n6959, n6961_1, n6963, n6965, n6967, n6969, n6971_1, n6973, n6975,
    n6977, n6978, n6979, n6980, n6981_1, n6982, n6983, n6985, n6987, n6989,
    n6991_1, n6993, n6995, n6997, n6999, n7001_1, n7003, n7005, n7007,
    n7009, n7011_1, n7013, n7015, n7017, n7019, n7021_1, n7023, n7025,
    n7027, n7029, n7031_1, n7033, n7035, n7037, n7039, n7041_1, n7043,
    n7045, n7047, n7049, n7051_1, n7053, n7055, n7057, n7059, n7061_1,
    n7062, n7063, n7065, n7067, n7069, n7070, n7071_1, n7073, n7075, n7077,
    n7078, n7079, n7081_1, n7083, n7085, n7086_1, n7087, n7089, n7091_1,
    n7093, n7094, n7095, n7097, n7099, n7101_1, n7102, n7103, n7105, n7107,
    n7109, n7110, n7111_1, n7113, n7115, n7117, n7118, n7119, n7121_1,
    n7123, n7125, n7127, n7129, n7131_1, n7132, n7134, n7136_1, n7138,
    n7139, n7141_1, n7143, n7145, n7147, n7149, n7151_1, n7153, n7155,
    n7157, n7158, n7160_1, n7162, n7164, n7165, n7167_1, n7169, n7171,
    n7173, n7175, n7177, n7179, n7181, n7183, n7184_1, n7186, n7188_1,
    n7190, n7191, n7193, n7195, n7197, n7199, n7201, n7203, n7205, n7207,
    n7209_1, n7210, n7212, n7214, n7216, n7217, n7219, n7221, n7223, n7225,
    n7227, n7229, n7231, n7233, n7235, n7236, n7238_1, n7240, n7242_1,
    n7243, n7245, n7247, n7249, n7251, n7253, n7255_1, n7257, n7259, n7261,
    n7262, n7264, n7266, n7268, n7269, n7271, n7273, n7275, n7277, n7279,
    n7281, n7283, n7285, n7287, n7288, n7290, n7292, n7294, n7295, n7297,
    n7299, n7301, n7303, n7305, n7307, n7309, n7311, n7313, n7314, n7316,
    n7318, n7320, n7321, n7323, n7325, n7327, n7329, n7331, n7333, n7335,
    n7337, n7339, n7341, n7343, n7345, n7347, n7349, n7351, n7353, n7355,
    n7357, n7359, n7361, n7363, n7365, n7367, n7369, n7371, n7373, n7375,
    n7377, n7379, n7381, n7383, n7385, n7387, n7389, n7391, n7393, n7395,
    n7397, n7399, n7401, n7403, n7405, n7407, n7409, n7411, n7413, n7415,
    n7417, n7419, n7421, n7423, n7425, n7427, n7429, n7431, n7433, n7435,
    n7437, n7439, n7441, n7443, n7445, n7447, n7449, n7451, n7453, n7455,
    n7457, n7459, n7461, n7463, n7465, n7467, n7469, n7471, n7473, n7475,
    n7477, n7479, n7481, n7483, n7485, n7487, n7489, n7491, n7493, n7495,
    n7497, n7499, n7501, n7503, n7505, n7507, n7509, n7511, n7513, n7515,
    n7517, n7519, n7521, n7523, n7525, n7527, n7529, n7531, n7533, n7535,
    n7537, n7539, n7541, n7543, n7545, n7547, n7549, n7551, n7553, n7555,
    n7557, n7559, n7561, n7563, n7565, n7567, n7569, n7571, n7573, n7575,
    n7577, n7579, n7581, n7583, n7585, n7587, n7589, n7591, n7593, n7595,
    n7597, n7599, n7601, n7603, n7605, n7607, n7609, n7611, n7613, n7615,
    n7617, n7619, n7621, n7622, n7624, n7626, n7628, n7630, n7632, n7634,
    n7636, n7638, n7640, n7642, n7644, n7646, n7648, n7650, n7652, n7654,
    n7656, n7658, n7660, n7662, n7664, n7666, n7668, n7670, n7672, n7674,
    n7676, n7678, n7680, n7682, n7684, n7686, n7688, n7690, n7692, n7694,
    n7696, n7698, n7700, n7702, n7704, n7706, n7708, n7710, n7712, n7714,
    n7716, n7718, n7720, n7722, n7724, n7726, n7728, n7730, n7732, n7734,
    n7736, n7738, n7740, n7742, n7744, n7746, n7748, n7750, n7752, n7754,
    n7756, n7758, n7760, n7762, n7764, n7766, n7768, n7770, n7772, n7774,
    n7776, n7778, n7780, n7782, n7784, n7786, n7788, n7790, n7792, n7794,
    n7796, n7798, n7800, n7802, n7804, n7806, n7808, n7810, n7812, n7814,
    n7816, n7818, n7820, n7822, n7824, n7826, n7828, n7830, n7832, n7834,
    n7836, n7838, n7840, n7842, n7844, n7846, n7848, n7850, n7852, n7854,
    n7856, n7858, n7860, n7862, n7864, n7866, n7868, n7870, n7872, n7874,
    n7876, n7878, n7880, n7882, n7884, n7886, n7888, n7890, n7892, n7894,
    n7896, n7898, n7900, n7902, n7904, n7906, n7908, n7910, n7912, n7914,
    n7916, n7918, n7920, n7922, n7924, n7926, n7928, n7930, n7932, n7934,
    n7936, n7938, n7940, n7942, n7944, n7946, n7948, n7950, n7952, n7954,
    n7956, n7958, n7960, n7962, n7964, n7966, n7968, n7970, n7972, n7974,
    n7976, n7978, n7980, n7982, n7984, n7986, n7988, n7990, n7992, n7994,
    n7996, n7998, n8000, n8002, n8004, n8006, n8008, n8010, n8012, n8014,
    n8016, n8018, n8020, n8022, n8024, n8026, n8028, n8030, n8032, n8034,
    n8036, n8038, n8040, n8042, n8044, n8046, n8048, n8050, n8052, n8054,
    n8056, n8058, n8060, n8062, n8064, n8066, n8068, n8070, n8072, n8074,
    n8076, n8078, n8080, n8082, n8084, n8086, n8088, n8090, n8092, n8094,
    n8096, n8098, n8100, n8102, n8104, n8106, n8108, n8110, n8112, n8114,
    n8116, n8118, n8120, n8122, n8124, n8126, n8128, n8130, n8132, n8134,
    n8136, n8138, n8140, n8142, n8144, n8146, n8148, n8150, n8152, n8154,
    n8156, n8158, n8160, n8162, n8164, n8166, n8168, n8170, n8172, n8174,
    n8176, n8178, n8180, n8182, n8184, n8186, n8188, n8190, n8192, n8194,
    n8196, n8198, n8200, n8202, n8204, n8206, n8208, n8210, n8212, n8214,
    n8216, n8218, n8220, n8222, n8224, n8226, n8228, n8230, n8232, n8234,
    n8236, n8238, n8240, n8242, n8244, n8246, n8248, n8250, n8252, n8254,
    n8256, n8258, n8260, n8262, n8264, n8266, n8268, n8270, n8272, n8274,
    n8276, n8278, n8280, n8282, n8284, n8286, n8288, n8290, n8292, n8294,
    n8296, n8298, n8300, n8302, n8304, n8306, n8308, n8310, n8312, n8314,
    n8316, n8318, n8320, n8322, n8324, n8326, n8328, n8330, n8332, n8334,
    n8336, n8338, n8340, n8342, n8344, n8346, n8348, n8350, n8352, n8354,
    n8356, n8358, n8360, n8362, n8364, n8366, n8368, n8370, n8372, n8374,
    n8376, n8378, n8380, n8382, n8384, n8386, n8388, n8390, n8392, n8394,
    n8396, n8398, n8400, n8402, n8404, n8406, n8408, n8410, n8412, n8414,
    n8416, n8418, n8420, n8422, n8424, n8426, n8428, n8430, n8432, n8434,
    n8436, n8438, n8440, n8442, n8444, n8446, n8448, n8450, n8451, n8452,
    n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
    n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
    n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
    n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
    n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
    n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
    n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
    n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
    n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
    n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
    n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
    n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
    n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
    n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
    n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8603,
    n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
    n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
    n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
    n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
    n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
    n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
    n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
    n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
    n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
    n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
    n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
    n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
    n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
    n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
    n8745, n8746, n8747, n8748, n8749, n8750, n8752, n8753, n8754, n8755,
    n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
    n8766, n8767, n270_1, n274_1, n279_1, n284_1, n289_1, n294_1, n299_1,
    n304_1, n309_1, n314_1, n319_1, n324_1, n329, n334_1, n339, n344,
    n349_1, n353_1, n358_1, n362_1, n366_1, n370_1, n374_1, n378_1, n382_1,
    n386, n390_1, n394, n398_1, n402_1, n406, n410_1, n414_1, n418_1,
    n422_1, n426_1, n430_1, n435_1, n440_1, n445_1, n450_1, n455_1, n460_1,
    n465, n470_1, n475_1, n480_1, n483_1, n488_1, n491_1, n496_1, n499_1,
    n504_1, n507, n512_1, n515_1, n520_1, n523_1, n528_1, n531_1, n536_1,
    n539_1, n544_1, n547_1, n552_1, n555_1, n560_1, n563_1, n568_1, n571_1,
    n576_1, n579, n584_1, n587_1, n592_1, n595_1, n600_1, n603_1, n608_1,
    n611_1, n616, n619_1, n624_1, n629_1, n634_1, n639_1, n644_1, n649_1,
    n654_1, n659_1, n664_1, n669_1, n674, n679_1, n684_1, n689_1, n694,
    n699_1, n704_1, n709_1, n714_1, n719_1, n724_1, n729, n734_1, n739_1,
    n744_1, n749_1, n754_1, n759_1, n764_1, n769_1, n774, n779, n784_1,
    n789_1, n794_1, n799_1, n804_1, n809_1, n814_1, n819_1, n824_1, n829_1,
    n834_1, n839_1, n844_1, n848_1, n853_1, n858_1, n863_1, n868_1, n872_1,
    n876_1, n880_1, n884_1, n888_1, n893_1, n898_1, n903_1, n908_1, n913_1,
    n918_1, n923_1, n928, n933_1, n938_1, n943_1, n948_1, n953_1, n958,
    n963_1, n968_1, n973_1, n978_1, n983_1, n988_1, n993_1, n998, n1003,
    n1008_1, n1013_1, n1018, n1023_1, n1028_1, n1033, n1038_1, n1043_1,
    n1048, n1053, n1058_1, n1063, n1068_1, n1073_1, n1078_1, n1083_1,
    n1088_1, n1093_1, n1098_1, n1103_1, n1108, n1113_1, n1118_1, n1123_1,
    n1128_1, n1133_1, n1138_1, n1143_1, n1148_1, n1153_1, n1158_1, n1163_1,
    n1168_1, n1173_1, n1178, n1183_1, n1188_1, n1193_1, n1198_1, n1203_1,
    n1208_1, n1213_1, n1218_1, n1223_1, n1228_1, n1233_1, n1238_1, n1243_1,
    n1248_1, n1253_1, n1258_1, n1263_1, n1268, n1273_1, n1278, n1283_1,
    n1288, n1293_1, n1298, n1303, n1308_1, n1313, n1318, n1323_1, n1328_1,
    n1333_1, n1338_1, n1343_1, n1348, n1353, n1358_1, n1363_1, n1368,
    n1373_1, n1378_1, n1383, n1388, n1393, n1398_1, n1403, n1408_1, n1413,
    n1418_1, n1423_1, n1428_1, n1433_1, n1438_1, n1443_1, n1448_1, n1453,
    n1458_1, n1463_1, n1468_1, n1473_1, n1478_1, n1483_1, n1488_1, n1493,
    n1498, n1503, n1508, n1513_1, n1518_1, n1523_1, n1528, n1533_1,
    n1537_1, n1542_1, n1546_1, n1551_1, n1555_1, n1560_1, n1564, n1569_1,
    n1573, n1578, n1582_1, n1587, n1591, n1596, n1600_1, n1604_1, n1608,
    n1613, n1618_1, n1623_1, n1627_1, n1631, n1635, n1639_1, n1643,
    n1647_1, n1651, n1655, n1659_1, n1663_1, n1667, n1671_1, n1675_1,
    n1679_1, n1683_1, n1687_1, n1691_1, n1695, n1699_1, n1703, n1707,
    n1711_1, n1715, n1719, n1724_1, n1729_1, n1734_1, n1739_1, n1743,
    n1747, n1752_1, n1756, n1761_1, n1765, n1770_1, n1774_1, n1779_1,
    n1783_1, n1788, n1792_1, n1797_1, n1801_1, n1806_1, n1811_1, n1816_1,
    n1821_1, n1825_1, n1829, n1833, n1838, n1843_1, n1848, n1853_1,
    n1858_1, n1863, n1867_1, n1871_1, n1875_1, n1879_1, n1883_1, n1888,
    n1892, n1897_1, n1902_1, n1906_1, n1911_1, n1915_1, n1920_1, n1925,
    n1930_1, n1935_1, n1940_1, n1945_1, n1950, n1955, n1960_1, n1965,
    n1970_1, n1975, n1980, n1985, n1990_1, n1995_1, n2000_1, n2005_1,
    n2010, n2015_1, n2020_1, n2025_1, n2030, n2035_1, n2040, n2045_1,
    n2050_1, n2054_1, n2059_1, n2064_1, n2067, n2072_1, n2077_1, n2082,
    n2087_1, n2092_1, n2097_1, n2102_1, n2107_1, n2112, n2117_1, n2122_1,
    n2127_1, n2132, n2137, n2142_1, n2147_1, n2152_1, n2157_1, n2162_1,
    n2167_1, n2172_1, n2177, n2182_1, n2187_1, n2192_1, n2197, n2202,
    n2207_1, n2212_1, n2217_1, n2222, n2227_1, n2232, n2237_1, n2242,
    n2247_1, n2252, n2257_1, n2262, n2267, n2272, n2277, n2282, n2287,
    n2292, n2297_1, n2302, n2307, n2312, n2317, n2322, n2327_1, n2332_1,
    n2337, n2342, n2347, n2352, n2357, n2362_1, n2367_1, n2372, n2377,
    n2382, n2387, n2391, n2395_1, n2399, n2404, n2409, n2414, n2419,
    n2424_1, n2429_1, n2434, n2439, n2444_1, n2449, n2454, n2459, n2464,
    n2469, n2474, n2479, n2484, n2489_1, n2494, n2499_1, n2504_1, n2509,
    n2514_1, n2519_1, n2524_1, n2529, n2534_1, n2539, n2544, n2549, n2554,
    n2559, n2564, n2569, n2574, n2579, n2584_1, n2589, n2594, n2599_1,
    n2604, n2609, n2614, n2619_1, n2624, n2629, n2634, n2639, n2644, n2649,
    n2654, n2659, n2664, n2669, n2674, n2679, n2684, n2689, n2694_1,
    n2699_1, n2704_1, n2709, n2714_1, n2719, n2724_1, n2729_1, n2734_1,
    n2739_1, n2744_1, n2749_1, n2754_1, n2759_1, n2764_1, n2769_1, n2774_1,
    n2779_1, n2784_1, n2789_1, n2794_1, n2799_1, n2804_1, n2809_1, n2814_1,
    n2819_1, n2824_1, n2829_1, n2834_1, n2839_1, n2844_1, n2849_1, n2854_1,
    n2859_1, n2864_1, n2869_1, n2874_1, n2879_1, n2884_1, n2889, n2894,
    n2899, n2904, n2909_1, n2914_1, n2919_1, n2924_1, n2929_1, n2934_1,
    n2939_1, n2944_1, n2949_1, n2954_1, n2959_1, n2964_1, n2969_1, n2974_1,
    n2979_1, n2984_1, n2989_1, n2994_1, n2999, n3004_1, n3009_1, n3014,
    n3019_1, n3024_1, n3029_1, n3034_1, n3039_1, n3043_1, n3048_1, n3052_1,
    n3057_1, n3061_1, n3066_1, n3070, n3075, n3079_1, n3084_1, n3088_1,
    n3093_1, n3097_1, n3102, n3106_1, n3110_1, n3114_1, n3119_1, n3124_1,
    n3129_1, n3133_1, n3137_1, n3141_1, n3145_1, n3149_1, n3153_1, n3157_1,
    n3161_1, n3165_1, n3169_1, n3173_1, n3177_1, n3181_1, n3185_1, n3189_1,
    n3193_1, n3197_1, n3201_1, n3205_1, n3209_1, n3213_1, n3217_1, n3221_1,
    n3225_1, n3230_1, n3235_1, n3240_1, n3245_1, n3249_1, n3253_1, n3258_1,
    n3262_1, n3267_1, n3271_1, n3276_1, n3280_1, n3285_1, n3289_1, n3294_1,
    n3298_1, n3303_1, n3307_1, n3312_1, n3317_1, n3322_1, n3327_1, n3331_1,
    n3335_1, n3339_1, n3344_1, n3349_1, n3354_1, n3359_1, n3364_1, n3369_1,
    n3373_1, n3377_1, n3381_1, n3385_1, n3389_1, n3394_1, n3398_1, n3403_1,
    n3408_1, n3412_1, n3417_1, n3421_1, n3426_1, n3431_1, n3436_1, n3441_1,
    n3446_1, n3451_1, n3456_1, n3461_1, n3466_1, n3471_1, n3476_1, n3481_1,
    n3486_1, n3491_1, n3496_1, n3501_1, n3506_1, n3511_1, n3516_1, n3521_1,
    n3526_1, n3531_1, n3536_1, n3541_1, n3546_1, n3551_1, n3556_1, n3560_1,
    n3565_1, n3570_1, n3573_1, n3578_1, n3583_1, n3588_1, n3593_1, n3598_1,
    n3603_1, n3608_1, n3613_1, n3618_1, n3623_1, n3628_1, n3632_1, n3636_1,
    n3641_1, n3646_1, n3651_1, n3656_1, n3661_1, n3666_1, n3671_1, n3676_1,
    n3681_1, n3686_1, n3691_1, n3696_1, n3701_1, n3706_1, n3711_1, n3716_1,
    n3721_1, n3726_1, n3731_1, n3736_1, n3741_1, n3746_1, n3751_1, n3756_1,
    n3761, n3766_1, n3771, n3776_1, n3781_1, n3786, n3791, n3796_1, n3801,
    n3806, n3811_1, n3816, n3821, n3826_1, n3831_1, n3836_1, n3841_1,
    n3846_1, n3851_1, n3856_1, n3861_1, n3866, n3871_1, n3876_1, n3881_1,
    n3886_1, n3891, n3896, n3901, n3906, n3911, n3916_1, n3921, n3926_1,
    n3931, n3936, n3941_1, n3946, n3951, n3956, n3961_1, n3966, n3971,
    n3976, n3981, n3986, n3991, n3996_1, n4001_1, n4006_1, n4011_1,
    n4016_1, n4021, n4026, n4031_1, n4036, n4041_1, n4046, n4051, n4056,
    n4061, n4066_1, n4071_1, n4076, n4081_1, n4086_1, n4091, n4096_1,
    n4101, n4106, n4111_1, n4116_1, n4121, n4126, n4131, n4136_1, n4141,
    n4146, n4151, n4156, n4161, n4166, n4171, n4176, n4181_1, n4186,
    n4191_1, n4196, n4201, n4206, n4211, n4216, n4221, n4226, n4231,
    n4236_1, n4241_1, n4246, n4251, n4256, n4261_1, n4266, n4271, n4276,
    n4281_1, n4286, n4291_1, n4296, n4301, n4306_1, n4311_1, n4316, n4321,
    n4326, n4331_1, n4336_1, n4341_1, n4346, n4351, n4356, n4361, n4366,
    n4371, n4376, n4381, n4386, n4391, n4396, n4401, n4406, n4411, n4416,
    n4421, n4426, n4431, n4436, n4441, n4446_1, n4451_1, n4456_1, n4461,
    n4466, n4471, n4476, n4481, n4486, n4491, n4496, n4501, n4506_1, n4511,
    n4516, n4521, n4526, n4531, n4536, n4541, n4546, n4550, n4555, n4559,
    n4564, n4568, n4573, n4577, n4582, n4586, n4591, n4595, n4600, n4604,
    n4609, n4613, n4617, n4621, n4626, n4631, n4636, n4640, n4644_1, n4648,
    n4652, n4656, n4660, n4664, n4668, n4672, n4676, n4680, n4684, n4688,
    n4692, n4696, n4700, n4704, n4708, n4712, n4716, n4720, n4724, n4728,
    n4732, n4737, n4742, n4747, n4752, n4756, n4760, n4765, n4769, n4774,
    n4778, n4783, n4787, n4792, n4796, n4801, n4805, n4810, n4814, n4819,
    n4824, n4829, n4834, n4838, n4842, n4846, n4851, n4856, n4861, n4866,
    n4871_1, n4876, n4880, n4884, n4888, n4892, n4896_1, n4901, n4905_1,
    n4910, n4915, n4919, n4924, n4928, n4933, n4938, n4943, n4948, n4953,
    n4958, n4963, n4968, n4973, n4978, n4983, n4988, n4993, n4998, n5003,
    n5008, n5013, n5018, n5023, n5028, n5033, n5038, n5043, n5048, n5053,
    n5058, n5063, n5067, n5072, n5077, n5080, n5085, n5090, n5095, n5100,
    n5105, n5110, n5115, n5120, n5125, n5130, n5135, n5140, n5145, n5150,
    n5155, n5160, n5165, n5170, n5175, n5180, n5185, n5190, n5195, n5200,
    n5205, n5210, n5215, n5220, n5225, n5230, n5235, n5240, n5245, n5250,
    n5255, n5260, n5265, n5270, n5275, n5280, n5285, n5290, n5295, n5300,
    n5305, n5310, n5315, n5320, n5325, n5330, n5335, n5340, n5345, n5350,
    n5355, n5360, n5365, n5370, n5375, n5380, n5385, n5390, n5395, n5400,
    n5405, n5410, n5415, n5420, n5425, n5430, n5435, n5440, n5445, n5450,
    n5455, n5460, n5465, n5470, n5475, n5480, n5485, n5490, n5495, n5500,
    n5505, n5510, n5515, n5520, n5525, n5530, n5535, n5540, n5545, n5550,
    n5555, n5560, n5565, n5570, n5575, n5580, n5585, n5590, n5595, n5600,
    n5605, n5610, n5615, n5620, n5625, n5630, n5635, n5640, n5645, n5650,
    n5655, n5660, n5665, n5670, n5675, n5680, n5685, n5690, n5695, n5700,
    n5705, n5710, n5715, n5720, n5725, n5730, n5735, n5740, n5745, n5750,
    n5755, n5760, n5765, n5770, n5775, n5780, n5785, n5790, n5795, n5800,
    n5805, n5810, n5815, n5819, n5823, n5828, n5833, n5838, n5843, n5848,
    n5853, n5858, n5863, n5868, n5873, n5878, n5883, n5888, n5893, n5898,
    n5903, n5908, n5913, n5918, n5923, n5928, n5933, n5938, n5943, n5948,
    n5953, n5958, n5963, n5968, n5973, n5978, n5983, n5988, n5993, n5998,
    n6003, n6008, n6013, n6018, n6023, n6028, n6033, n6038, n6043, n6048,
    n6053, n6057, n6062, n6066, n6071, n6075, n6080, n6084, n6089, n6093,
    n6098, n6102, n6107, n6111, n6116, n6120, n6124, n6128, n6133, n6138,
    n6143, n6147, n6151, n6155, n6159, n6163, n6167, n6171, n6175, n6179,
    n6183, n6187, n6191, n6195, n6199, n6203, n6207, n6211, n6215, n6219,
    n6223, n6227, n6231, n6235, n6239, n6244, n6249, n6254, n6259, n6263,
    n6267, n6272, n6276, n6281, n6285, n6290, n6294, n6299, n6303, n6308,
    n6312, n6317, n6321, n6326, n6331, n6336, n6341, n6345, n6349, n6353,
    n6358, n6363, n6368, n6373, n6378, n6383, n6387, n6391, n6395, n6399,
    n6403, n6408, n6412, n6417, n6422, n6426, n6431, n6435, n6440, n6445,
    n6450, n6455, n6460, n6465, n6470, n6475, n6480, n6485, n6490, n6495,
    n6500, n6505, n6510, n6515, n6520, n6525, n6530, n6535, n6540, n6545,
    n6550, n6555, n6560, n6565, n6570, n6574, n6579, n6584, n6587, n6592,
    n6597, n6602, n6607, n6612, n6617, n6622, n6627, n6632, n6637, n6642,
    n6647, n6652, n6657, n6662, n6667, n6672, n6677, n6682, n6687, n6692,
    n6697, n6702, n6707, n6712, n6717, n6722, n6727, n6732, n6737, n6742,
    n6747, n6752, n6757, n6762, n6767, n6772, n6777, n6782, n6787, n6792,
    n6797, n6802, n6807, n6812, n6817, n6822, n6827, n6832, n6837, n6842,
    n6847, n6852, n6857, n6862, n6867, n6872, n6877, n6882, n6887, n6892,
    n6897, n6902, n6907, n6912, n6917, n6922, n6926, n6931, n6936, n6941,
    n6946, n6951, n6956, n6961, n6966, n6971, n6976, n6981, n6986, n6991,
    n6996, n7001, n7006, n7011, n7016, n7021, n7026, n7031, n7036, n7041,
    n7046, n7051, n7056, n7061, n7066, n7071, n7076, n7081, n7086, n7091,
    n7096, n7101, n7106, n7111, n7116, n7121, n7126, n7131, n7136, n7141,
    n7146, n7151, n7156, n7160, n7163, n7167, n7172, n7176, n7180, n7184,
    n7188, n7192, n7196, n7200, n7204, n7209, n7213, n7218, n7222, n7226,
    n7230, n7234, n7238, n7242, n7246, n7250, n7255, n7260;
  assign Pg27380 = ~n893_1;
  assign Pg26149 = ~n6140;
  assign Pg26135 = ~n853_1;
  assign Pg26104 = ~n6148;
  assign Pg25489 = ~n7621;
  assign n858_1 = ~Pg3233 | Pg3230;
  assign Pg25435 = ~n863_1;
  assign Pg24734 = ~n868_1;
  assign Pg16496 = ~n4652_1;
  assign n4530 = ~Pg8269 ^ ~Pg8268;
  assign n4531_1 = ~Pg8271 ^ ~Pg8270;
  assign n4532 = ~n4530 ^ ~n4531_1;
  assign n4533 = ~Pg8262 ^ ~Pg8264;
  assign n4534 = ~Pg8265 ^ ~Pg8266;
  assign n4535 = ~n4533 ^ ~n4534;
  assign n4536_1 = ~Pg8259 ^ ~Pg8261;
  assign n4537 = ~Pg8260 ^ ~Pg8263;
  assign n4538 = ~n4536_1 ^ ~n4537;
  assign n4539 = ~Pg8272 ^ ~Pg8273;
  assign n4540 = ~Pg8275 ^ ~Pg8274;
  assign n4541_1 = ~n4539 ^ ~n4540;
  assign n4542 = (~Ng1315 | ~Ng324) & (~\[1605]  | ~Ng394);
  assign n4543 = n4542 & (~\[1603]  | ~Ng396);
  assign n4544 = (~Ng1315 | ~Ng383) & (~\[1605]  | ~Ng379);
  assign n4545 = n4544 & (~\[1603]  | ~Ng381);
  assign n4546_1 = (~Ng1315 | ~Ng1011) & (~\[1605]  | ~Ng1081);
  assign n4547 = n4546_1 & (~\[1603]  | ~Ng1083);
  assign n4548 = (~Ng1315 | ~Ng368) & (~\[1605]  | ~Ng364);
  assign n4549 = n4548 & (~\[1603]  | ~Ng366);
  assign n4550_1 = (~Ng1315 | ~Ng1070) & (~\[1605]  | ~Ng1066);
  assign n4551 = n4550_1 & (~\[1603]  | ~Ng1068);
  assign n4552 = (~Ng1315 | ~Ng1705) & (~\[1605]  | ~Ng1775);
  assign n4553 = n4552 & (~\[1603]  | ~Ng1777);
  assign n4554 = (~Ng1315 | ~Ng353) & (~\[1605]  | ~Ng349);
  assign n4555_1 = n4554 & (~\[1603]  | ~Ng351);
  assign n4556 = (~Ng1315 | ~Ng1055) & (~\[1605]  | ~Ng1051);
  assign n4557 = n4556 & (~\[1603]  | ~Ng1053);
  assign n4558 = (~Ng1315 | ~Ng1764) & (~\[1605]  | ~Ng1760);
  assign n4559_1 = n4558 & (~\[1603]  | ~Ng1762);
  assign n4560 = (~Ng1315 | ~Ng2399) & (~\[1605]  | ~Ng2469);
  assign n4561 = n4560 & (~\[1603]  | ~Ng2471);
  assign n4562 = (~Ng1315 | ~Ng1040) & (~\[1605]  | ~Ng1036);
  assign n4563 = n4562 & (~\[1603]  | ~Ng1038);
  assign n4564_1 = (~Ng1315 | ~Ng1749) & (~\[1605]  | ~Ng1745);
  assign n4565 = n4564_1 & (~\[1603]  | ~Ng1747);
  assign n4566 = (~Ng1315 | ~Ng2458) & (~\[1605]  | ~Ng2454);
  assign n4567 = n4566 & (~\[1603]  | ~Ng2456);
  assign n4568_1 = (~Ng1315 | ~Ng1734) & (~\[1605]  | ~Ng1730);
  assign n4569 = n4568_1 & (~\[1603]  | ~Ng1732);
  assign n4570 = (~Ng1315 | ~Ng2443) & (~\[1605]  | ~Ng2439);
  assign n4571 = n4570 & (~\[1603]  | ~Ng2441);
  assign n4572 = (~Ng1315 | ~Ng2428) & (~\[1605]  | ~Ng2424);
  assign n4573_1 = n4572 & (~\[1603]  | ~Ng2426);
  assign n4574 = (~Ng1315 | ~Ng496) & (~\[1605]  | ~Ng490);
  assign n4575 = n4574 & (~\[1603]  | ~Ng493);
  assign n4576 = (~Ng1315 | ~Ng1183) & (~\[1605]  | ~Ng1177);
  assign n4577_1 = n4576 & (~\[1603]  | ~Ng1180);
  assign n4578 = (~Ng1315 | ~Ng1877) & (~\[1605]  | ~Ng1871);
  assign n4579 = n4578 & (~\[1603]  | ~Ng1874);
  assign n4580 = (~Ng1315 | ~Ng2571) & (~\[1605]  | ~Ng2565);
  assign n4581 = n4580 & (~\[1603]  | ~Ng2568);
  assign n4582_1 = (~Ng853 | Ng447) & (~\[1612]  | Ng448);
  assign n4583 = n4582_1 & (~\[1594]  | Ng449);
  assign n4584 = (~Ng853 | Ng402) & (~\[1612]  | Ng403);
  assign n4585 = n4584 & (~\[1594]  | Ng404);
  assign n4586_1 = (~\[1605]  | Ng479) & (~\[1603]  | Ng477);
  assign n1888 = n4586_1 & (~Ng1315 | Ng478);
  assign n4588 = (~\[1605]  | Ng464) & (~\[1603]  | Ng480);
  assign n1902_1 = n4588 & (~Ng1315 | Ng484);
  assign n4590 = (~Ng853 | Ng1134) & (~\[1612]  | Ng1135);
  assign n4591_1 = n4590 & (~\[1594]  | Ng1136);
  assign n4592 = (~Ng853 | Ng1089) & (~\[1612]  | Ng1090);
  assign n4593 = n4592 & (~\[1594]  | Ng1091);
  assign n4594 = (~\[1605]  | Ng1166) & (~\[1603]  | Ng1164);
  assign n3394_1 = n4594 & (~Ng1315 | Ng1165);
  assign n4596 = (~\[1605]  | Ng488) & (~\[1603]  | Ng486);
  assign n1911_1 = n4596 & (~Ng1315 | Ng487);
  assign n4598 = (~\[1605]  | Ng1151) & (~\[1603]  | Ng1167);
  assign n3408_1 = n4598 & (~Ng1315 | Ng1171);
  assign n4600_1 = (~Ng853 | Ng1828) & (~\[1612]  | Ng1829);
  assign n4601 = n4600_1 & (~\[1594]  | Ng1830);
  assign n4602 = (~Ng853 | Ng1783) & (~\[1612]  | Ng1784);
  assign n4603 = n4602 & (~\[1594]  | Ng1785);
  assign n4604_1 = (~\[1605]  | Ng1860) & (~\[1603]  | Ng1858);
  assign n4901 = n4604_1 & (~Ng1315 | Ng1859);
  assign n4606 = (~Ng1315 | ~Ng573) & (~\[1605]  | ~Ng569);
  assign n1739_1 = n4606 & (~\[1603]  | ~Ng571);
  assign n4608 = (~\[1605]  | Ng1175) & (~\[1603]  | Ng1173);
  assign n3417_1 = n4608 & (~Ng1315 | Ng1174);
  assign n4610 = (~\[1605]  | Ng1845) & (~\[1603]  | Ng1861);
  assign n4915 = n4610 & (~Ng1315 | Ng1865);
  assign n4612 = (~Ng853 | Ng2522) & (~\[1612]  | Ng2523);
  assign n4613_1 = n4612 & (~\[1594]  | Ng2524);
  assign n4614 = (~Ng853 | Ng2477) & (~\[1612]  | Ng2478);
  assign n4615 = n4614 & (~\[1594]  | Ng2479);
  assign n4616 = (~\[1605]  | Ng2554) & (~\[1603]  | Ng2552);
  assign n6408 = n4616 & (~Ng1315 | Ng2553);
  assign n4618 = (~Ng1315 | ~Ng1259) & (~\[1605]  | ~Ng1255);
  assign n3245_1 = n4618 & (~\[1603]  | ~Ng1257);
  assign n4620 = (~\[1605]  | Ng1869) & (~\[1603]  | Ng1867);
  assign n4924 = n4620 & (~Ng1315 | Ng1868);
  assign n4622 = (~\[1605]  | Ng2539) & (~\[1603]  | Ng2555);
  assign n6422 = n4622 & (~Ng1315 | Ng2559);
  assign n4624 = (~Ng853 | Ng321) & (~\[1612]  | Ng322);
  assign n4625 = n4624 & (~\[1594]  | Ng323);
  assign n4626_1 = (~Ng1315 | ~Ng1953) & (~\[1605]  | ~Ng1949);
  assign n4752 = n4626_1 & (~\[1603]  | ~Ng1951);
  assign n4628 = (~\[1605]  | Ng2563) & (~\[1603]  | Ng2561);
  assign n6431 = n4628 & (~Ng1315 | Ng2562);
  assign n4630 = (~Ng1315 | ~Ng489) & (~\[1605]  | ~Ng565);
  assign n1875_1 = n4630 & (~\[1603]  | ~Ng567);
  assign n4632 = (~Ng853 | Ng1008) & (~\[1612]  | Ng1009);
  assign n4633 = n4632 & (~\[1594]  | Ng1010);
  assign n4634 = (~Ng1315 | ~Ng2647) & (~\[1605]  | ~Ng2643);
  assign n6259 = n4634 & (~\[1603]  | ~Ng2645);
  assign n4636_1 = (~Ng1315 | ~Ng1176) & (~\[1605]  | ~Ng1251);
  assign n3381_1 = n4636_1 & (~\[1603]  | ~Ng1253);
  assign n4638 = (~Ng853 | Ng1702) & (~\[1612]  | Ng1703);
  assign n4639 = n4638 & (~\[1594]  | Ng1704);
  assign n4640_1 = (~Ng1315 | ~Ng1870) & (~\[1605]  | ~Ng1945);
  assign n4888 = n4640_1 & (~\[1603]  | ~Ng1947);
  assign n4642 = (~Ng853 | Ng2396) & (~\[1612]  | Ng2397);
  assign n4643 = n4642 & (~\[1594]  | Ng2398);
  assign n4644 = (~Ng1315 | ~Ng2564) & (~\[1605]  | ~Ng2639);
  assign n6395 = n4644 & (~\[1603]  | ~Ng2641);
  assign n4646 = (~Ng853 | Ng141) & (~\[1594]  | Ng143);
  assign n4647 = n4646 & (~\[1612]  | Ng142);
  assign n4648_1 = (~Ng853 | Ng144) & (~\[1594]  | Ng146);
  assign n4649 = n4648_1 & (~\[1612]  | Ng145);
  assign n4650 = (~Ng853 | Ng829) & (~\[1594]  | Ng831);
  assign n4651 = n4650 & (~\[1612]  | Ng830);
  assign n4652_1 = Ng2987 & (~Pg5388 | Ng2986);
  assign n4653 = (~Ng853 | Ng147) & (~\[1594]  | Ng149);
  assign n4654 = n4653 & (~\[1612]  | Ng148);
  assign n4655 = (~Ng853 | Ng832) & (~\[1594]  | Ng834);
  assign n4656_1 = n4655 & (~\[1612]  | Ng833);
  assign n4657 = (~Ng853 | Ng1523) & (~\[1594]  | Ng1525);
  assign n4658 = n4657 & (~\[1612]  | Ng1524);
  assign n4659 = (~Ng853 | Ng150) & (~\[1594]  | Ng152);
  assign n4660_1 = n4659 & (~\[1612]  | Ng151);
  assign n4661 = (~\[1594]  | ~Ng216) & (~Ng853 | ~Ng219);
  assign n4662 = n4661 & (~\[1612]  | ~Ng213);
  assign n4663 = (~Ng853 | Ng835) & (~\[1594]  | Ng837);
  assign n4664_1 = n4663 & (~\[1612]  | Ng836);
  assign n4665 = (~Ng853 | Ng1526) & (~\[1594]  | Ng1528);
  assign n4666 = n4665 & (~\[1612]  | Ng1527);
  assign n4667 = (~Ng853 | Ng2217) & (~\[1594]  | Ng2219);
  assign n4668_1 = n4667 & (~\[1612]  | Ng2218);
  assign n4669 = (~Ng853 | Ng153) & (~\[1612]  | Ng154);
  assign n4670 = n4669 & (~\[1594]  | Ng155);
  assign n4671 = (~\[1612]  | ~Ng222) & (~\[1594]  | ~Ng225);
  assign n4672_1 = n4671 & (~Ng853 | ~Ng228);
  assign n4673 = (~Ng853 | Ng838) & (~\[1612]  | Ng839);
  assign n4674 = n4673 & (~\[1594]  | Ng840);
  assign n4675 = (~\[1612]  | ~Ng900) & (~\[1594]  | ~Ng903);
  assign n4676_1 = n4675 & (~Ng853 | ~Ng906);
  assign n4677 = (~Ng853 | Ng1529) & (~\[1612]  | Ng1530);
  assign n4678 = n4677 & (~\[1594]  | Ng1531);
  assign n4679 = (~Ng853 | Ng2220) & (~\[1612]  | Ng2221);
  assign n4680_1 = n4679 & (~\[1594]  | Ng2222);
  assign n4681 = (~Ng853 | Ng156) & (~\[1612]  | Ng157);
  assign n4682 = n4681 & (~\[1594]  | Ng158);
  assign n4683 = (~Ng853 | ~Ng237) & (~\[1612]  | ~Ng231);
  assign n4684_1 = n4683 & (~\[1594]  | ~Ng234);
  assign n4685 = (~Ng1315 | Ng698) & (~\[1605]  | Ng699);
  assign n4686 = n4685 & (~\[1603]  | Ng700);
  assign n4687 = (~Ng1315 | Ng725) & (~\[1605]  | Ng726);
  assign n4688_1 = n4687 & (~\[1603]  | Ng727);
  assign n4689 = (~Ng853 | Ng841) & (~\[1612]  | Ng842);
  assign n4690 = n4689 & (~\[1594]  | Ng843);
  assign n4691 = (~Ng853 | ~Ng915) & (~\[1612]  | ~Ng909);
  assign n4692_1 = n4691 & (~\[1594]  | ~Ng912);
  assign n4693 = (~Ng853 | Ng1532) & (~\[1612]  | Ng1533);
  assign n4694 = n4693 & (~\[1594]  | Ng1534);
  assign n4695 = (~Ng853 | ~Ng1600) & (~\[1612]  | ~Ng1594);
  assign n4696_1 = n4695 & (~\[1594]  | ~Ng1597);
  assign n4697 = (~Ng853 | Ng2223) & (~\[1612]  | Ng2224);
  assign n4698 = n4697 & (~\[1594]  | Ng2225);
  assign n4699 = (~Ng853 | Ng159) & (~\[1612]  | Ng160);
  assign n4700_1 = n4699 & (~\[1594]  | Ng161);
  assign n4701 = (~Ng853 | ~Ng246) & (~\[1612]  | ~Ng240);
  assign n4702 = n4701 & (~\[1594]  | ~Ng243);
  assign n4703 = (~Ng1315 | Ng701) & (~\[1605]  | Ng702);
  assign n4704_1 = n4703 & (~\[1603]  | Ng703);
  assign n4705 = (~Ng853 | Ng844) & (~\[1612]  | Ng845);
  assign n4706 = n4705 & (~\[1594]  | Ng846);
  assign n4707 = (~Ng853 | ~Ng924) & (~\[1612]  | ~Ng918);
  assign n4708_1 = n4707 & (~\[1594]  | ~Ng921);
  assign n4709 = (~Ng1315 | Ng1384) & (~\[1605]  | Ng1385);
  assign n4710 = n4709 & (~\[1603]  | Ng1386);
  assign n4711 = (~Ng1315 | Ng1411) & (~\[1605]  | Ng1412);
  assign n4712_1 = n4711 & (~\[1603]  | Ng1413);
  assign n4713 = (~Ng853 | Ng1535) & (~\[1612]  | Ng1536);
  assign n4714 = n4713 & (~\[1594]  | Ng1537);
  assign n4715 = (~Ng853 | ~Ng1609) & (~\[1612]  | ~Ng1603);
  assign n4716_1 = n4715 & (~\[1594]  | ~Ng1606);
  assign n4717 = (~Ng853 | Ng2226) & (~\[1612]  | Ng2227);
  assign n4718 = n4717 & (~\[1594]  | Ng2228);
  assign n4719 = (~Ng853 | ~Ng2294) & (~\[1612]  | ~Ng2288);
  assign n4720_1 = n4719 & (~\[1594]  | ~Ng2291);
  assign n4721 = (~Ng853 | Ng129) & (~\[1612]  | Ng130);
  assign n4722 = n4721 & (~\[1594]  | Ng131);
  assign n4723 = (~Ng853 | Ng162) & (~\[1612]  | Ng163);
  assign n4724_1 = n4723 & (~\[1594]  | Ng164);
  assign n4725 = (~Ng853 | ~Ng255) & (~\[1612]  | ~Ng249);
  assign n4726 = n4725 & (~\[1594]  | ~Ng252);
  assign n4727 = (~Ng1315 | Ng704) & (~\[1605]  | Ng705);
  assign n4728_1 = n4727 & (~\[1603]  | Ng706);
  assign n4729 = (~Ng853 | Ng847) & (~\[1612]  | Ng848);
  assign n4730 = n4729 & (~\[1594]  | Ng849);
  assign n4731 = (~Ng853 | ~Ng933) & (~\[1612]  | ~Ng927);
  assign n4732_1 = n4731 & (~\[1594]  | ~Ng930);
  assign n4733 = (~Ng1315 | Ng1387) & (~\[1605]  | Ng1388);
  assign n4734 = n4733 & (~\[1603]  | Ng1389);
  assign n4735 = (~Ng853 | Ng1538) & (~\[1612]  | Ng1539);
  assign n4736 = n4735 & (~\[1594]  | Ng1540);
  assign n4737_1 = (~Ng853 | ~Ng1618) & (~\[1612]  | ~Ng1612);
  assign n4738 = n4737_1 & (~\[1594]  | ~Ng1615);
  assign n4739 = (~Ng1315 | Ng2078) & (~\[1605]  | Ng2079);
  assign n4740 = n4739 & (~\[1603]  | Ng2080);
  assign n4741 = (~Ng1315 | Ng2105) & (~\[1605]  | Ng2106);
  assign n4742_1 = n4741 & (~\[1603]  | Ng2107);
  assign n4743 = (~Ng853 | Ng2229) & (~\[1612]  | Ng2230);
  assign n4744 = n4743 & (~\[1594]  | Ng2231);
  assign n4745 = (~Ng853 | ~Ng2303) & (~\[1612]  | ~Ng2297);
  assign n4746 = n4745 & (~\[1594]  | ~Ng2300);
  assign n4747_1 = (~Ng853 | Ng132) & (~\[1612]  | Ng133);
  assign n4748 = n4747_1 & (~\[1594]  | Ng134);
  assign n4749 = (~Ng853 | ~Ng264) & (~\[1612]  | ~Ng258);
  assign n4750 = n4749 & (~\[1594]  | ~Ng261);
  assign n4751 = (~Ng853 | Ng11499) & (~\[1612]  | Ng11497);
  assign n4752_1 = n4751 & (~\[1594]  | Ng11498);
  assign n4753 = (~Ng853 | ~Ng435) & (~\[1612]  | ~Ng429);
  assign n4754 = n4753 & (~\[1594]  | ~Ng432);
  assign n4755 = (~Ng1315 | Ng707) & (~\[1605]  | Ng708);
  assign n4756_1 = n4755 & (~\[1603]  | Ng709);
  assign n4757 = (~Ng853 | Ng817) & (~\[1612]  | Ng818);
  assign n4758 = n4757 & (~\[1594]  | Ng819);
  assign n4759 = (~Ng853 | Ng850) & (~\[1612]  | Ng851);
  assign n4760_1 = n4759 & (~\[1594]  | Ng852);
  assign n4761 = (~Ng853 | ~Ng942) & (~\[1612]  | ~Ng936);
  assign n4762 = n4761 & (~\[1594]  | ~Ng939);
  assign n4763 = (~Ng1315 | Ng1390) & (~\[1605]  | Ng1391);
  assign n4764 = n4763 & (~\[1603]  | Ng1392);
  assign n4765_1 = (~Ng853 | Ng1541) & (~\[1612]  | Ng1542);
  assign n4766 = n4765_1 & (~\[1594]  | Ng1543);
  assign n4767 = (~Ng853 | ~Ng1627) & (~\[1612]  | ~Ng1621);
  assign n4768 = n4767 & (~\[1594]  | ~Ng1624);
  assign n4769_1 = (~Ng1315 | Ng2081) & (~\[1605]  | Ng2082);
  assign n4770 = n4769_1 & (~\[1603]  | Ng2083);
  assign n4771 = (~Ng853 | Ng2232) & (~\[1612]  | Ng2233);
  assign n4772 = n4771 & (~\[1594]  | Ng2234);
  assign n4773 = (~Ng853 | ~Ng2312) & (~\[1612]  | ~Ng2306);
  assign n4774_1 = n4773 & (~\[1594]  | ~Ng2309);
  assign n4775 = (~Ng1315 | Ng2772) & (~\[1605]  | Ng2773);
  assign n4776 = n4775 & (~\[1603]  | Ng2774);
  assign n4777 = (~Ng1315 | Ng2799) & (~\[1605]  | Ng2800);
  assign n4778_1 = n4777 & (~\[1603]  | Ng2801);
  assign n4779 = (~Ng853 | ~Ng192) & (~\[1612]  | ~Ng186);
  assign n4780 = n4779 & (~\[1594]  | ~Ng189);
  assign n4781 = (~Ng853 | ~Ng273) & (~\[1612]  | ~Ng267);
  assign n4782 = n4781 & (~\[1594]  | ~Ng270);
  assign n4783_1 = (~Ng853 | Ng11502) & (~\[1612]  | Ng11500);
  assign n4784 = n4783_1 & (~\[1594]  | Ng11501);
  assign n4785 = (~Ng853 | ~Ng444) & (~\[1612]  | ~Ng438);
  assign n4786 = n4785 & (~\[1594]  | ~Ng441);
  assign n4787_1 = (~Ng1315 | Ng710) & (~\[1605]  | Ng711);
  assign n4788 = n4787_1 & (~\[1603]  | Ng712);
  assign n4789 = (~Ng853 | Ng820) & (~\[1612]  | Ng821);
  assign n4790 = n4789 & (~\[1594]  | Ng822);
  assign n4791 = (~Ng853 | ~Ng951) & (~\[1612]  | ~Ng945);
  assign n4792_1 = n4791 & (~\[1594]  | ~Ng948);
  assign n4793 = (~Ng853 | Ng11526) & (~\[1612]  | Ng11524);
  assign n4794 = n4793 & (~\[1594]  | Ng11525);
  assign n4795 = (~Ng853 | ~Ng1122) & (~\[1612]  | ~Ng1116);
  assign n4796_1 = n4795 & (~\[1594]  | ~Ng1119);
  assign n4797 = (~Ng1315 | Ng1393) & (~\[1605]  | Ng1394);
  assign n4798 = n4797 & (~\[1603]  | Ng1395);
  assign n4799 = (~Ng853 | Ng1511) & (~\[1612]  | Ng1512);
  assign n4800 = n4799 & (~\[1594]  | Ng1513);
  assign n4801_1 = (~Ng853 | Ng1544) & (~\[1612]  | Ng1545);
  assign n4802 = n4801_1 & (~\[1594]  | Ng1546);
  assign n4803 = (~Ng853 | ~Ng1636) & (~\[1612]  | ~Ng1630);
  assign n4804 = n4803 & (~\[1594]  | ~Ng1633);
  assign n4805_1 = (~Ng1315 | Ng2084) & (~\[1605]  | Ng2085);
  assign n4806 = n4805_1 & (~\[1603]  | Ng2086);
  assign n4807 = (~Ng853 | Ng2235) & (~\[1612]  | Ng2236);
  assign n4808 = n4807 & (~\[1594]  | Ng2237);
  assign n4809 = (~Ng853 | ~Ng2321) & (~\[1612]  | ~Ng2315);
  assign n4810_1 = n4809 & (~\[1594]  | ~Ng2318);
  assign n4811 = (~Ng1315 | Ng2775) & (~\[1605]  | Ng2776);
  assign n4812 = n4811 & (~\[1603]  | Ng2777);
  assign n4813 = (~Ng853 | ~Ng201) & (~\[1612]  | ~Ng195);
  assign n4814_1 = n4813 & (~\[1594]  | ~Ng198);
  assign n4815 = (~Ng853 | Ng11505) & (~\[1612]  | Ng11503);
  assign n4816 = n4815 & (~\[1594]  | Ng11504);
  assign n4817 = (~Ng1315 | Ng713) & (~\[1605]  | Ng714);
  assign n4818 = n4817 & (~\[1603]  | Ng715);
  assign n4819_1 = (~Ng1315 | Ng731) & (~\[1605]  | Ng732);
  assign n4820 = n4819_1 & (~\[1603]  | Ng733);
  assign n4821 = (~Ng853 | ~Ng879) & (~\[1612]  | ~Ng873);
  assign n4822 = n4821 & (~\[1594]  | ~Ng876);
  assign n4823 = (~Ng853 | ~Ng960) & (~\[1612]  | ~Ng954);
  assign n4824_1 = n4823 & (~\[1594]  | ~Ng957);
  assign n4825 = (~Ng853 | Ng11529) & (~\[1612]  | Ng11527);
  assign n4826 = n4825 & (~\[1594]  | Ng11528);
  assign n4827 = (~Ng853 | ~Ng1131) & (~\[1612]  | ~Ng1125);
  assign n4828 = n4827 & (~\[1594]  | ~Ng1128);
  assign n4829_1 = (~Ng1315 | Ng1396) & (~\[1605]  | Ng1397);
  assign n4830 = n4829_1 & (~\[1603]  | Ng1398);
  assign n4831 = (~Ng853 | Ng1514) & (~\[1612]  | Ng1515);
  assign n4832 = n4831 & (~\[1594]  | Ng1516);
  assign n4833 = (~Ng853 | ~Ng1645) & (~\[1612]  | ~Ng1639);
  assign n4834_1 = n4833 & (~\[1594]  | ~Ng1642);
  assign n4835 = (~Ng853 | Ng11553) & (~\[1612]  | Ng11551);
  assign n4836 = n4835 & (~\[1594]  | Ng11552);
  assign n4837 = (~Ng853 | ~Ng1816) & (~\[1612]  | ~Ng1810);
  assign n4838_1 = n4837 & (~\[1594]  | ~Ng1813);
  assign n4839 = (~Ng1315 | Ng2087) & (~\[1605]  | Ng2088);
  assign n4840 = n4839 & (~\[1603]  | Ng2089);
  assign n4841 = (~Ng853 | Ng2205) & (~\[1612]  | Ng2206);
  assign n4842_1 = n4841 & (~\[1594]  | Ng2207);
  assign n4843 = (~Ng853 | Ng2238) & (~\[1612]  | Ng2239);
  assign n4844 = n4843 & (~\[1594]  | Ng2240);
  assign n4845 = (~Ng853 | ~Ng2330) & (~\[1612]  | ~Ng2324);
  assign n4846_1 = n4845 & (~\[1594]  | ~Ng2327);
  assign n4847 = (~Ng1315 | Ng2778) & (~\[1605]  | Ng2779);
  assign n4848 = n4847 & (~\[1603]  | Ng2780);
  assign n4849 = (~Ng853 | ~Ng210) & (~\[1612]  | ~Ng204);
  assign n4850 = n4849 & (~\[1594]  | ~Ng207);
  assign n4851_1 = (~Ng853 | Ng11508) & (~\[1612]  | Ng11506);
  assign n4852 = n4851_1 & (~\[1594]  | Ng11507);
  assign n4853 = (~Ng1315 | Ng716) & (~\[1605]  | Ng717);
  assign n4854 = n4853 & (~\[1603]  | Ng718);
  assign n4855 = (~Ng853 | ~Ng888) & (~\[1612]  | ~Ng882);
  assign n4856_1 = n4855 & (~\[1594]  | ~Ng885);
  assign n4857 = (~Ng853 | Ng11532) & (~\[1612]  | Ng11530);
  assign n4858 = n4857 & (~\[1594]  | Ng11531);
  assign n4859 = (~Ng1315 | Ng1399) & (~\[1605]  | Ng1400);
  assign n4860 = n4859 & (~\[1603]  | Ng1401);
  assign n4861_1 = (~Ng1315 | Ng1417) & (~\[1605]  | Ng1418);
  assign n4862 = n4861_1 & (~\[1603]  | Ng1419);
  assign n4863 = (~Ng853 | ~Ng1573) & (~\[1612]  | ~Ng1567);
  assign n4864 = n4863 & (~\[1594]  | ~Ng1570);
  assign n4865 = (~Ng853 | ~Ng1654) & (~\[1612]  | ~Ng1648);
  assign n4866_1 = n4865 & (~\[1594]  | ~Ng1651);
  assign n4867 = (~Ng853 | Ng11556) & (~\[1612]  | Ng11554);
  assign n4868 = n4867 & (~\[1594]  | Ng11555);
  assign n4869 = (~Ng853 | ~Ng1825) & (~\[1612]  | ~Ng1819);
  assign n4870 = n4869 & (~\[1594]  | ~Ng1822);
  assign n4871 = (~Ng1315 | Ng2090) & (~\[1605]  | Ng2091);
  assign n4872 = n4871 & (~\[1603]  | Ng2092);
  assign n4873 = (~Ng853 | Ng2208) & (~\[1612]  | Ng2209);
  assign n4874 = n4873 & (~\[1594]  | Ng2210);
  assign n4875 = (~Ng853 | ~Ng2339) & (~\[1612]  | ~Ng2333);
  assign n4876_1 = n4875 & (~\[1594]  | ~Ng2336);
  assign n4877 = (~Ng853 | Ng11580) & (~\[1612]  | Ng11578);
  assign n4878 = n4877 & (~\[1594]  | Ng11579);
  assign n4879 = (~Ng853 | ~Ng2510) & (~\[1612]  | ~Ng2504);
  assign n4880_1 = n4879 & (~\[1594]  | ~Ng2507);
  assign n4881 = (~Ng1315 | Ng2781) & (~\[1605]  | Ng2782);
  assign n4882 = n4881 & (~\[1603]  | Ng2783);
  assign n4883 = (~Ng853 | Ng168) & (~\[1594]  | Ng170);
  assign n4884_1 = n4883 & (~\[1612]  | Ng169);
  assign n4885 = (~Ng1315 | Ng719) & (~\[1605]  | Ng720);
  assign n4886 = n4885 & (~\[1603]  | Ng721);
  assign n4887 = (~Ng853 | ~Ng897) & (~\[1612]  | ~Ng891);
  assign n4888_1 = n4887 & (~\[1594]  | ~Ng894);
  assign n4889 = (~Ng853 | Ng11535) & (~\[1612]  | Ng11533);
  assign n4890 = n4889 & (~\[1594]  | Ng11534);
  assign n4891 = (~Ng1315 | Ng1402) & (~\[1605]  | Ng1403);
  assign n4892_1 = n4891 & (~\[1603]  | Ng1404);
  assign n4893 = (~Ng853 | ~Ng1582) & (~\[1612]  | ~Ng1576);
  assign n4894 = n4893 & (~\[1594]  | ~Ng1579);
  assign n4895 = (~Ng853 | Ng11559) & (~\[1612]  | Ng11557);
  assign n4896 = n4895 & (~\[1594]  | Ng11558);
  assign n4897 = (~Ng1315 | Ng2093) & (~\[1605]  | Ng2094);
  assign n4898 = n4897 & (~\[1603]  | Ng2095);
  assign n4899 = (~Ng1315 | Ng2111) & (~\[1605]  | Ng2112);
  assign n4900 = n4899 & (~\[1603]  | Ng2113);
  assign n4901_1 = (~Ng853 | ~Ng2267) & (~\[1612]  | ~Ng2261);
  assign n4902 = n4901_1 & (~\[1594]  | ~Ng2264);
  assign n4903 = (~Ng853 | ~Ng2348) & (~\[1612]  | ~Ng2342);
  assign n4904 = n4903 & (~\[1594]  | ~Ng2345);
  assign n4905 = (~Ng853 | Ng11583) & (~\[1612]  | Ng11581);
  assign n4906 = n4905 & (~\[1594]  | Ng11582);
  assign n4907 = (~Ng853 | ~Ng2519) & (~\[1612]  | ~Ng2513);
  assign n4908 = n4907 & (~\[1594]  | ~Ng2516);
  assign n4909 = (~Ng1315 | Ng2784) & (~\[1605]  | Ng2785);
  assign n4910_1 = n4909 & (~\[1603]  | Ng2786);
  assign n4911 = (~Ng1315 | Ng722) & (~\[1605]  | Ng723);
  assign n4912 = n4911 & (~\[1603]  | Ng724);
  assign n4913 = (~Ng853 | Ng856) & (~\[1594]  | Ng858);
  assign n4914 = n4913 & (~\[1612]  | Ng857);
  assign n4915_1 = (~Ng1315 | Ng1405) & (~\[1605]  | Ng1406);
  assign n4916 = n4915_1 & (~\[1603]  | Ng1407);
  assign n4917 = (~Ng853 | ~Ng1591) & (~\[1612]  | ~Ng1585);
  assign n4918 = n4917 & (~\[1594]  | ~Ng1588);
  assign n4919_1 = (~Ng853 | Ng11562) & (~\[1612]  | Ng11560);
  assign n4920 = n4919_1 & (~\[1594]  | Ng11561);
  assign n4921 = (~Ng1315 | Ng2096) & (~\[1605]  | Ng2097);
  assign n4922 = n4921 & (~\[1603]  | Ng2098);
  assign n4923 = (~Ng853 | ~Ng2276) & (~\[1612]  | ~Ng2270);
  assign n4924_1 = n4923 & (~\[1594]  | ~Ng2273);
  assign n4925 = (~Ng853 | Ng11586) & (~\[1612]  | Ng11584);
  assign n4926 = n4925 & (~\[1594]  | Ng11585);
  assign n4927 = (~Ng1315 | Ng2787) & (~\[1605]  | Ng2788);
  assign n4928_1 = n4927 & (~\[1603]  | Ng2789);
  assign n4929 = (~Ng1315 | Ng2805) & (~\[1605]  | Ng2806);
  assign n4930 = n4929 & (~\[1603]  | Ng2807);
  assign n4931 = (~Ng1315 | Ng1408) & (~\[1605]  | Ng1409);
  assign n4932 = n4931 & (~\[1603]  | Ng1410);
  assign n4933_1 = (~Ng853 | Ng1550) & (~\[1612]  | Ng1551);
  assign n4934 = n4933_1 & (~\[1594]  | Ng1552);
  assign n4935 = (~Ng1315 | Ng2099) & (~\[1605]  | Ng2100);
  assign n4936 = n4935 & (~\[1603]  | Ng2101);
  assign n4937 = (~Ng853 | ~Ng2285) & (~\[1612]  | ~Ng2279);
  assign n4938_1 = n4937 & (~\[1594]  | ~Ng2282);
  assign n4939 = (~Ng853 | Ng11589) & (~\[1612]  | Ng11587);
  assign n4940 = n4939 & (~\[1594]  | Ng11588);
  assign n4941 = (~Ng1315 | Ng2790) & (~\[1605]  | Ng2791);
  assign n4942 = n4941 & (~\[1603]  | Ng2792);
  assign n4943_1 = (~Ng1315 | Ng2102) & (~\[1605]  | Ng2103);
  assign n4944 = n4943_1 & (~\[1603]  | Ng2104);
  assign n4945 = (~Ng853 | Ng2244) & (~\[1612]  | Ng2245);
  assign n4946 = n4945 & (~\[1594]  | Ng2246);
  assign n4947 = (~Ng1315 | Ng2793) & (~\[1605]  | Ng2794);
  assign n4948_1 = n4947 & (~\[1603]  | Ng2795);
  assign n4949 = (~Ng853 | Ng314) & (~\[1612]  | Ng312);
  assign n4950 = n4949 & (~\[1594]  | Ng313);
  assign n4951 = (~Ng1315 | Ng2796) & (~\[1605]  | Ng2797);
  assign n4952 = n4951 & (~\[1603]  | Ng2798);
  assign n4953_1 = (~Ng853 | Ng317) & (~\[1612]  | Ng315);
  assign n4954 = n4953_1 & (~\[1594]  | Ng316);
  assign n4955 = (~Ng853 | Ng1001) & (~\[1612]  | Ng999);
  assign n4956 = n4955 & (~\[1594]  | Ng1000);
  assign n4957 = (~Ng853 | Ng320) & (~\[1612]  | Ng318);
  assign n4958_1 = n4957 & (~\[1594]  | Ng319);
  assign n4959 = (~Ng853 | Ng1004) & (~\[1612]  | Ng1002);
  assign n4960 = n4959 & (~\[1594]  | Ng1003);
  assign n4961 = (~Ng853 | Ng1695) & (~\[1612]  | Ng1693);
  assign n4962 = n4961 & (~\[1594]  | Ng1694);
  assign n4963_1 = (~Ng1315 | ~Ng620) & (~\[1605]  | ~Ng614);
  assign n4964 = n4963_1 & (~\[1603]  | ~Ng617);
  assign n4965 = (~Ng853 | Ng1007) & (~\[1612]  | Ng1005);
  assign n4966 = n4965 & (~\[1594]  | Ng1006);
  assign n4967 = (~Ng853 | Ng1698) & (~\[1612]  | Ng1696);
  assign n4968_1 = n4967 & (~\[1594]  | Ng1697);
  assign n4969 = (~Ng853 | Ng2389) & (~\[1612]  | Ng2387);
  assign n4970 = n4969 & (~\[1594]  | Ng2388);
  assign n4971 = (~Ng1315 | ~Ng1306) & (~\[1605]  | ~Ng1300);
  assign n4972 = n4971 & (~\[1603]  | ~Ng1303);
  assign n4973_1 = (~Ng853 | Ng1701) & (~\[1612]  | Ng1699);
  assign n4974 = n4973_1 & (~\[1594]  | Ng1700);
  assign n4975 = (~Ng853 | Ng2392) & (~\[1612]  | Ng2390);
  assign n4976 = n4975 & (~\[1594]  | Ng2391);
  assign n4977 = (~Ng1315 | ~Ng2000) & (~\[1605]  | ~Ng1994);
  assign n4978_1 = n4977 & (~\[1603]  | ~Ng1997);
  assign n4979 = (~Ng853 | Ng2395) & (~\[1612]  | Ng2393);
  assign n4980 = n4979 & (~\[1594]  | Ng2394);
  assign n4981 = (~Ng1315 | ~Ng2694) & (~\[1605]  | ~Ng2688);
  assign n4982 = n4981 & (~\[1603]  | ~Ng2691);
  assign n4983_1 = (~Ng1315 | Ng575) & (~\[1605]  | Ng576);
  assign n4984 = n4983_1 & (~\[1603]  | Ng577);
  assign n4985 = (~Ng1315 | Ng578) & (~\[1605]  | Ng579);
  assign n4986 = n4985 & (~\[1603]  | Ng580);
  assign n4987 = (~Ng1315 | Ng1261) & (~\[1605]  | Ng1262);
  assign n4988_1 = n4987 & (~\[1603]  | Ng1263);
  assign n4989 = (~Ng853 | ~Ng414) & (~\[1612]  | ~Ng408);
  assign n4990 = n4989 & (~\[1594]  | ~Ng411);
  assign n4991 = (~Ng1315 | Ng581) & (~\[1605]  | Ng582);
  assign n4992 = n4991 & (~\[1603]  | Ng583);
  assign n4993_1 = (~Ng1315 | Ng1264) & (~\[1605]  | Ng1265);
  assign n4994 = n4993_1 & (~\[1603]  | Ng1266);
  assign n4995 = (~Ng1315 | Ng1955) & (~\[1605]  | Ng1956);
  assign n4996 = n4995 & (~\[1603]  | Ng1957);
  assign n4997 = (~Ng853 | ~Ng423) & (~\[1612]  | ~Ng417);
  assign n4998_1 = n4997 & (~\[1594]  | ~Ng420);
  assign n4999 = (~Ng1315 | Ng584) & (~\[1605]  | Ng585);
  assign n5000 = n4999 & (~\[1603]  | Ng586);
  assign n5001 = (~Ng853 | ~Ng1101) & (~\[1612]  | ~Ng1095);
  assign n5002 = n5001 & (~\[1594]  | ~Ng1098);
  assign n5003_1 = (~Ng1315 | Ng1267) & (~\[1605]  | Ng1268);
  assign n5004 = n5003_1 & (~\[1603]  | Ng1269);
  assign n5005 = (~Ng1315 | Ng1958) & (~\[1605]  | Ng1959);
  assign n5006 = n5005 & (~\[1603]  | Ng1960);
  assign n5007 = (~Ng1315 | Ng2649) & (~\[1605]  | Ng2650);
  assign n5008_1 = n5007 & (~\[1603]  | Ng2651);
  assign n5009 = (~Ng853 | ~Ng1110) & (~\[1612]  | ~Ng1104);
  assign n5010 = n5009 & (~\[1594]  | ~Ng1107);
  assign n5011 = (~Ng1315 | Ng1270) & (~\[1605]  | Ng1271);
  assign n5012 = n5011 & (~\[1603]  | Ng1272);
  assign n5013_1 = (~Ng853 | ~Ng1795) & (~\[1612]  | ~Ng1789);
  assign n5014 = n5013_1 & (~\[1594]  | ~Ng1792);
  assign n5015 = (~Ng1315 | Ng1961) & (~\[1605]  | Ng1962);
  assign n5016 = n5015 & (~\[1603]  | Ng1963);
  assign n5017 = (~Ng1315 | Ng2652) & (~\[1605]  | Ng2653);
  assign n5018_1 = n5017 & (~\[1603]  | Ng2654);
  assign n5019 = (~Ng853 | Ng171) & (~\[1594]  | Ng173);
  assign n5020 = n5019 & (~\[1612]  | Ng172);
  assign n5021 = (~Ng853 | ~Ng1804) & (~\[1612]  | ~Ng1798);
  assign n5022 = n5021 & (~\[1594]  | ~Ng1801);
  assign n5023_1 = (~Ng1315 | Ng1964) & (~\[1605]  | Ng1965);
  assign n5024 = n5023_1 & (~\[1603]  | Ng1966);
  assign n5025 = (~Ng853 | ~Ng2489) & (~\[1612]  | ~Ng2483);
  assign n5026 = n5025 & (~\[1594]  | ~Ng2486);
  assign n5027 = (~Ng1315 | Ng2655) & (~\[1605]  | Ng2656);
  assign n5028_1 = n5027 & (~\[1603]  | Ng2657);
  assign n5029 = (~Ng853 | Ng174) & (~\[1612]  | Ng175);
  assign n5030 = n5029 & (~\[1594]  | Ng176);
  assign n5031 = (~Ng853 | Ng859) & (~\[1612]  | Ng860);
  assign n5032 = n5031 & (~\[1594]  | Ng861);
  assign n5033_1 = (~Ng853 | ~Ng2498) & (~\[1612]  | ~Ng2492);
  assign n5034 = n5033_1 & (~\[1594]  | ~Ng2495);
  assign n5035 = (~Ng1315 | Ng2658) & (~\[1605]  | Ng2659);
  assign n5036 = n5035 & (~\[1603]  | Ng2660);
  assign n5037 = (~Ng853 | Ng862) & (~\[1612]  | Ng863);
  assign n5038_1 = n5037 & (~\[1594]  | Ng864);
  assign n5039 = (~Ng853 | Ng1553) & (~\[1612]  | Ng1554);
  assign n5040 = n5039 & (~\[1594]  | Ng1555);
  assign n5041 = (~Ng853 | Ng1556) & (~\[1612]  | Ng1557);
  assign n5042 = n5041 & (~\[1594]  | Ng1558);
  assign n5043_1 = (~Ng853 | Ng2247) & (~\[1612]  | Ng2248);
  assign n5044 = n5043_1 & (~\[1594]  | Ng2249);
  assign n5045 = (~Ng853 | Ng2250) & (~\[1612]  | Ng2251);
  assign n5046 = n5045 & (~\[1594]  | Ng2252);
  assign n5047 = Ng2879 & (~Pg8021 | Ng2929);
  assign n358_1 = ~n5047;
  assign n5049 = (~Ng853 | Ng426) & (~\[1612]  | Ng427);
  assign n5050 = n5049 & (~\[1594]  | Ng428);
  assign n5051 = (~Ng853 | Ng1113) & (~\[1612]  | Ng1114);
  assign n5052 = n5051 & (~\[1594]  | Ng1115);
  assign n5053_1 = (~Ng1315 | ~Ng611) & (~\[1605]  | ~Ng605);
  assign n5054 = n5053_1 & (~\[1603]  | ~Ng608);
  assign n5055 = (~Ng853 | Ng1807) & (~\[1612]  | Ng1808);
  assign n5056 = n5055 & (~\[1594]  | Ng1809);
  assign n5057 = (~Ng1315 | ~Ng1297) & (~\[1605]  | ~Ng1291);
  assign n5058_1 = n5057 & (~\[1603]  | ~Ng1294);
  assign n5059 = (~Ng853 | Ng2501) & (~\[1612]  | Ng2502);
  assign n5060 = n5059 & (~\[1594]  | Ng2503);
  assign n5061 = (~Ng1315 | ~Ng1991) & (~\[1605]  | ~Ng1985);
  assign n5062 = n5061 & (~\[1603]  | ~Ng1988);
  assign n5063_1 = (~Ng1315 | ~Ng2685) & (~\[1605]  | ~Ng2679);
  assign n5064 = n5063_1 & (~\[1603]  | ~Ng2682);
  assign n5065 = ~Ng557 & (Ng525 | Ng510);
  assign n5066 = ~Ng510 & (Ng525 | Ng557);
  assign n5067_1 = ~Ng1243 & (Ng1211 | Ng1196);
  assign n5068 = ~Ng1196 & (Ng1211 | Ng1243);
  assign n5069 = ~Ng1937 & (Ng1905 | Ng1890);
  assign n5070 = ~Ng1890 & (Ng1905 | Ng1937);
  assign n5071 = ~Ng2631 & (Ng2599 | Ng2584);
  assign n5072_1 = ~Ng2584 & (Ng2599 | Ng2631);
  assign n5073 = n1739_1 | ~Ng185 | ~Ng524;
  assign n5074 = (~Ng1315 | ~Ng593) & (~\[1605]  | ~Ng587);
  assign n5075 = n5073 & n5074 & (~\[1603]  | ~Ng590);
  assign n5076 = n3245_1 | ~Ng185 | ~Ng1210;
  assign n5077_1 = (~Ng1315 | ~Ng1279) & (~\[1605]  | ~Ng1273);
  assign n5078 = n5076 & n5077_1 & (~\[1603]  | ~Ng1276);
  assign n5079 = n4752 | ~Ng185 | ~Ng1904;
  assign n5080_1 = (~Ng1315 | ~Ng1973) & (~\[1605]  | ~Ng1967);
  assign n5081 = n5079 & n5080_1 & (~\[1603]  | ~Ng1970);
  assign n5082 = n6259 | ~Ng185 | ~Ng2598;
  assign n5083 = (~Ng1315 | ~Ng2667) & (~\[1605]  | ~Ng2661);
  assign n5084 = n5082 & n5083 & (~\[1603]  | ~Ng2664);
  assign n274_1 = ~Pg51 & Ng13457;
  assign n279_1 = ~Pg51 & Ng2817;
  assign n5087 = n6275 & (~Ng659 | n6276_1);
  assign n2127_1 = ~n5087;
  assign n5089 = n6275 & (~Ng1345 | n6276_1);
  assign n3646_1 = ~n5089;
  assign n5091 = n6275 & (~Ng2039 | n6276_1);
  assign n5140 = ~n5091;
  assign n5093 = n6275 & (~Ng2733 | n6276_1);
  assign n6647 = ~n5093;
  assign n284_1 = Pg51 | Ng2933;
  assign n6922 = Ng3079 | Pg3234;
  assign n5097 = n6270 & (n6271 | ~Ng554);
  assign n1724_1 = ~n5097;
  assign n5099 = n6270 & (n6271 | ~Ng1240);
  assign n3230_1 = ~n5099;
  assign n5101 = n6270 & (n6271 | ~Ng1934);
  assign n4737 = ~n5101;
  assign n5103 = n6270 & (n6271 | ~Ng2628);
  assign n6244 = ~n5103;
  assign n5105_1 = n6274 ^ ~Ng640;
  assign n5106 = ~\[1603]  | ~Ng630;
  assign n2132 = n5105_1 & n5106;
  assign n5108 = n6273 ^ ~Ng1326;
  assign n5109 = ~\[1603]  | ~Ng1316;
  assign n3651_1 = n5108 & n5109;
  assign n5111 = n6272_1 ^ ~Ng2020;
  assign n5112 = ~\[1603]  | ~Ng2010;
  assign n5145 = n5111 & n5112;
  assign n5114 = n6269 ^ ~Ng2714;
  assign n5115_1 = ~\[1603]  | ~Ng2704;
  assign n6652 = n5114 & n5115_1;
  assign n5117 = n6258 | Pg8021;
  assign n5118 = ~Ng2883 ^ ~Ng13457;
  assign n289_1 = n5117 | n5118;
  assign n6912 = ~Pg3234 & Ng13475;
  assign n6917 = ~Pg3234 & Ng3054;
  assign n5122 = ~n6266 ^ ~Ng633;
  assign n2137 = n5122 & n5106;
  assign n5124 = ~n6264 ^ ~Ng1319;
  assign n3656_1 = n5124 & n5109;
  assign n5126 = ~n4950 | n4954 | n4958_1;
  assign n5127 = Ng2896 | Ng2900 | Ng2908 | Ng2892 | Ng2903;
  assign n5128 = n5126 & (n5127 | ~n6231_1);
  assign n5129 = ~n6262 ^ ~Ng2013;
  assign n5150 = n5129 & n5112;
  assign n5131 = ~n4956 | n4960 | n4966;
  assign n5132 = n5131 & (n5127 | ~n6227_1);
  assign n5133 = ~n6260 ^ ~Ng2707;
  assign n6657 = n5133 & n5115_1;
  assign n5135_1 = ~n4962 | n4968_1 | n4974;
  assign n5136 = n5135_1 & (n5127 | ~n6223_1);
  assign n5137 = ~n4970 | n4976 | n4980;
  assign n5138 = n5137 & (n5127 | ~n6219_1);
  assign n5139 = n5117 & (Pg8021 | n6237);
  assign n5140_1 = ~n6258 ^ ~Ng2912;
  assign n324_1 = n5139 | n5140_1;
  assign n5142 = n6192 & (~n8750 | (~n4575 & ~n5054));
  assign n2059_1 = ~n5142;
  assign n5144 = n6234 & (Pg3234 | n6233);
  assign n5145_1 = ~n6256 ^ ~Ng3018;
  assign n7141 = n5144 | n5145_1;
  assign n5147 = n6187_1 & (~n8750 | (~n4577_1 & ~n5058_1));
  assign n3565_1 = ~n5147;
  assign n5149 = n6182 & (~n8750 | (~n4579 & ~n5062));
  assign n5072 = ~n5149;
  assign n5151 = ~Ng2888 ^ ~n6268;
  assign n294_1 = ~n5117 & n5151;
  assign n5153 = ~\[1605]  | ~Ng630;
  assign n5154 = \[1605]  & n6579_1;
  assign n2377 = n5153 & (Ng738 | n5154);
  assign n5156 = n6177 & (~n8750 | (~n4581 & ~n5064));
  assign n6579 = ~n5156;
  assign n5158 = \[1603]  & n6579_1;
  assign n2382 = n5106 & (Ng739 | n5158);
  assign n5160_1 = ~\[1605]  | ~Ng1316;
  assign n5161 = \[1605]  & n6578;
  assign n3896 = n5160_1 & (Ng1424 | n5161);
  assign n5163 = n8547 & n8548 & (~\[1605]  | Ng729);
  assign n5164 = n4820 & n5163 & (~\[1603]  | Ng730);
  assign n5165_1 = ~Ng1315 | ~Ng630;
  assign n5166 = Ng1315 & n6579_1;
  assign n2387 = n5165_1 & (Ng737 | n5166);
  assign n5168 = \[1603]  & n6578;
  assign n3901 = n5109 & (Ng1425 | n5168);
  assign n5170_1 = ~\[1605]  | ~Ng2010;
  assign n5171 = \[1605]  & n6577;
  assign n5390 = n5170_1 & (Ng2118 | n5171);
  assign n5173 = n8544 & n8545 & (~\[1605]  | Ng1415);
  assign n5174 = n4862 & n5173 & (~\[1603]  | Ng1416);
  assign n5175_1 = ~Ng1315 | ~Ng1316;
  assign n5176 = Ng1315 & n6578;
  assign n3906 = n5175_1 & (Ng1423 | n5176);
  assign n5178 = \[1603]  & n6577;
  assign n5395 = n5112 & (Ng2119 | n5178);
  assign n5180_1 = ~\[1605]  | ~Ng2704;
  assign n5181 = \[1605]  & n6575;
  assign n6897 = n5180_1 & (Ng2812 | n5181);
  assign n5183 = n8541 & n8542 & (~\[1605]  | Ng2109);
  assign n5184 = n4900 & n5183 & (~\[1603]  | Ng2110);
  assign n5185_1 = ~Ng1315 | ~Ng2010;
  assign n5186 = Ng1315 & n6577;
  assign n5400 = n5185_1 & (Ng2117 | n5186);
  assign n5188 = \[1603]  & n6575;
  assign n6902 = n5115_1 & (Ng2813 | n5188);
  assign n5190_1 = n8538 & n8539 & (~\[1605]  | Ng2803);
  assign n5191 = n4930 & n5190_1 & (~\[1603]  | Ng2804);
  assign n5192 = ~Ng1315 | ~Ng2704;
  assign n5193 = Ng1315 & n6575;
  assign n6907 = n5192 & (Ng2811 | n5193);
  assign n868_1 = ~n858_1 & (n5978_1 | Ng3123);
  assign n5196 = ~Ng653 ^ ~n6267_1;
  assign n2142_1 = n5196 & n5106;
  assign n5198 = ~Ng1339 ^ ~n6265;
  assign n3661_1 = n5198 & n5109;
  assign n5200_1 = ~n6572 ^ ~Ng3006;
  assign n7116 = n5200_1 & ~n6234;
  assign n5202 = ~Ng2033 ^ ~n6263_1;
  assign n5155 = n5202 & n5112;
  assign n5204 = ~Ng2727 ^ ~n6261;
  assign n6662 = n5204 & n5115_1;
  assign n5206 = ~Ng2917 ^ ~n6259_1;
  assign n329 = ~n5139 & n5206;
  assign n5208 = ~n6254_1 ^ ~Ng2896;
  assign n299_1 = ~n5117 & n5208;
  assign n5210_1 = ~Ng3028 ^ ~n6257;
  assign n7146 = ~n5144 & n5210_1;
  assign n863_1 = ~n858_1 & (n5978_1 | Ng3125);
  assign n5213 = ~n6250 ^ ~Ng646;
  assign n2147_1 = n5213 & n5106;
  assign n5215_1 = ~n6247 ^ ~Ng1332;
  assign n3666_1 = n5215_1 & n5109;
  assign n5217 = ~n6244_1 ^ ~Ng2026;
  assign n5160 = n5217 & n5112;
  assign n5219 = ~n6240 ^ ~Ng2720;
  assign n6667 = n5219 & n5115_1;
  assign n5221 = n6253 ^ ~Ng3002;
  assign n7121 = n5221 & ~n6234;
  assign n5223 = ~n6235_1 ^ ~Ng3036;
  assign n7151 = ~n5144 & n5223;
  assign n5225_1 = ~Ng2892 ^ ~n6255;
  assign n304_1 = ~n5117 & n5225_1;
  assign n5227 = ~n6238 ^ ~Ng2924;
  assign n334_1 = ~n5139 & n5227;
  assign n5229 = n6252 ^ ~Ng88;
  assign n5230_1 = n6521 | n5127;
  assign n1263_1 = n5229 & n5230_1;
  assign n5232 = n6249_1 ^ ~Ng776;
  assign n2769_1 = n5232 & n5230_1;
  assign n5234 = n6246 ^ ~Ng1462;
  assign n4276 = n5234 & n5230_1;
  assign n5236 = n6243 ^ ~Ng2156;
  assign n5770 = n5236 & n5230_1;
  assign n853_1 = n6039 & n6038_1 & n6037 & n6035 & n6036 & n6040 & n6041 & n6042;
  assign n5239 = ~Ng660 ^ ~n6251;
  assign n2152_1 = n5239 & n5106;
  assign n5241 = ~Ng1346 ^ ~n6248;
  assign n3671_1 = n5241 & n5109;
  assign n5243 = Ng3013 ^ ~n6573;
  assign n7126 = n5243 & ~n6234;
  assign n5245_1 = ~Ng2040 ^ ~n6245;
  assign n5165 = n5245_1 & n5112;
  assign n5247 = ~Ng2734 ^ ~n6241;
  assign n6672 = n5247 & n5115_1;
  assign n5249 = ~Ng2920 ^ ~n6239_1;
  assign n339 = ~n5139 & n5249;
  assign n5251 = ~n6574_1 ^ ~Ng2903;
  assign n309_1 = ~n5117 & n5251;
  assign n5253 = ~Ng3032 ^ ~n6236;
  assign n7156 = ~n5144 & n5253;
  assign n5255_1 = ~n6215_1 ^ ~Ng83;
  assign n1268 = n5255_1 & n5230_1;
  assign n5257 = ~n6211_1 ^ ~Ng771;
  assign n2774_1 = n5257 & n5230_1;
  assign n5259 = ~n6207_1 ^ ~Ng1457;
  assign n4281_1 = n5259 & n5230_1;
  assign n5261 = ~n6203_1 ^ ~Ng2151;
  assign n5775 = n5261 & n5230_1;
  assign n5263 = ~n6213 ^ ~Ng672;
  assign n2157_1 = n5263 & n5106;
  assign n5265_1 = ~n6209 ^ ~Ng1358;
  assign n3676_1 = n5265_1 & n5109;
  assign n5267 = ~n6205 ^ ~Ng2052;
  assign n5170 = n5267 & n5112;
  assign n5269 = ~n6201 ^ ~Ng2746;
  assign n6677 = n5269 & n5115_1;
  assign n5271 = n6197 ^ ~Ng3010;
  assign n7131 = n5271 & ~n6234;
  assign n5273 = ~Ng2900 ^ ~n6199_1;
  assign n314_1 = ~n5117 & n5273;
  assign n5275_1 = ~Ng79 ^ ~n6216;
  assign n1273_1 = n5275_1 & n5230_1;
  assign n5277 = ~Ng767 ^ ~n6212;
  assign n2779_1 = n5277 & n5230_1;
  assign n5279 = ~Ng1453 ^ ~n6208;
  assign n4286 = n5279 & n5230_1;
  assign n5281 = ~Ng2147 ^ ~n6204;
  assign n5780 = n5281 & n5230_1;
  assign n893_1 = ~n858_1 & n5977 & (Ng185 | n5978_1);
  assign n5284 = ~Ng666 ^ ~n6214;
  assign n2162_1 = n5284 & n5106;
  assign n5286 = ~Ng1352 ^ ~n6210;
  assign n3681_1 = n5286 & n5109;
  assign n7136 = ~n6234 & ~n6584_1;
  assign n5289 = ~Ng2046 ^ ~n6206;
  assign n5175 = n5289 & n5112;
  assign n5291 = ~Ng2740 ^ ~n6202;
  assign n6682 = n5291 & n5115_1;
  assign n5293 = ~Ng2908 ^ ~n6200;
  assign n319_1 = ~n5117 & n5293;
  assign n5295_1 = ~n6175_1 ^ ~Ng74;
  assign n1278 = n5295_1 & n5230_1;
  assign n5297 = ~n6168 ^ ~Ng762;
  assign n2784_1 = n5297 & n5230_1;
  assign n5299 = ~n6161 ^ ~Ng1448;
  assign n4291_1 = n5299 & n5230_1;
  assign n5301 = ~n6154 ^ ~Ng2142;
  assign n5785 = n5301 & n5230_1;
  assign n5303 = ~n6564 ^ ~Ng679;
  assign n2167_1 = n5303 & n5106;
  assign n5305_1 = ~n6560_1 ^ ~Ng1365;
  assign n3686_1 = n5305_1 & n5109;
  assign n5307 = ~n6556 ^ ~Ng2059;
  assign n5180 = n5307 & n5112;
  assign n5309 = ~n6550_1 ^ ~Ng2753;
  assign n6687 = n5309 & n5115_1;
  assign n5311 = n5918_1 & n5916 & n5917;
  assign n5312 = n4672_1 ^ ~n5947;
  assign n5313 = n5311 & n5312;
  assign n5314 = n5898_1 & n5896 & n5897;
  assign n5315_1 = n4692_1 ^ ~n5940;
  assign n5316 = n5314 & n5315_1;
  assign n5317 = n5878_1 & n5876 & n5877;
  assign n5318 = n4716_1 ^ ~n5933_1;
  assign n5319 = n5317 & n5318;
  assign n5320_1 = n5858_1 & n5856 & n5857;
  assign n5321 = n4746 ^ ~n5926;
  assign n5322 = n5320_1 & n5321;
  assign n5323 = ~Ng70 ^ ~n6176;
  assign n1283_1 = n5323 & n5230_1;
  assign n5325_1 = ~Ng758 ^ ~n6169;
  assign n2789_1 = n5325_1 & n5230_1;
  assign n5327 = ~Ng1444 ^ ~n6162;
  assign n4296 = n5327 & n5230_1;
  assign n5329 = ~Ng2138 ^ ~n6155_1;
  assign n5790 = n5329 & n5230_1;
  assign n5331 = ~Ng686 ^ ~n6109;
  assign n2172_1 = n5331 & n5106;
  assign n5333 = ~Ng1372 ^ ~n6087;
  assign n3691_1 = n5333 & n5109;
  assign n5335_1 = ~Ng2066 ^ ~n6065;
  assign n5185 = n5335_1 & n5112;
  assign n5337 = ~Ng2760 ^ ~n6043_1;
  assign n6692 = n5337 & n5115_1;
  assign n5339 = n6571 | ~n4583 | ~Ng2257;
  assign n5340_1 = \[1612]  & ~n6174;
  assign n1443_1 = (~\[1612]  | n5339) & (n5340_1 | Ng448);
  assign n5342 = \[1594]  & ~n6174;
  assign n1448_1 = (~\[1594]  | n5339) & (Ng449 | n5342);
  assign n5344 = n6570_1 | ~n4591_1 | ~Ng2257;
  assign n5345_1 = \[1612]  & ~n6167_1;
  assign n2949_1 = (~\[1612]  | n5344) & (n5345_1 | Ng1135);
  assign n5347 = Ng853 & ~n6174;
  assign n1453 = (~Ng853 | n5339) & (n5347 | Ng447);
  assign n5349 = \[1594]  & ~n6167_1;
  assign n2954_1 = (~\[1594]  | n5344) & (Ng1136 | n5349);
  assign n5351 = n6569 | ~n4601 | ~Ng2257;
  assign n5352 = \[1612]  & ~n6160;
  assign n4456_1 = (~\[1612]  | n5351) & (n5352 | Ng1829);
  assign n5354 = Ng853 & ~n6167_1;
  assign n2959_1 = (~Ng853 | n5344) & (n5354 | Ng1134);
  assign n5356 = \[1594]  & ~n6160;
  assign n4461 = (~\[1594]  | n5351) & (Ng1830 | n5356);
  assign n5358 = n6568 | ~n4613_1 | ~Ng2257;
  assign n5359 = \[1612]  & ~n6153;
  assign n5963 = (~\[1612]  | n5358) & (n5359 | Ng2523);
  assign n5361 = Ng853 & ~n6160;
  assign n4466 = (~Ng853 | n5351) & (n5361 | Ng1828);
  assign n5363 = \[1594]  & ~n6153;
  assign n5968 = (~\[1594]  | n5358) & (Ng2524 | n5363);
  assign n5365_1 = Ng853 & ~n6153;
  assign n5973 = (~Ng853 | n5358) & (n5365_1 | Ng2522);
  assign n5367 = ~n6033_1 ^ ~Ng65;
  assign n1288 = n5367 & n5230_1;
  assign n5369 = ~n6029 ^ ~Ng753;
  assign n2794_1 = n5369 & n5230_1;
  assign n5371 = ~n6025 ^ ~Ng1439;
  assign n4301 = n5371 & n5230_1;
  assign n5373 = ~n6021 ^ ~Ng2133;
  assign n5795 = n5373 & n5230_1;
  assign n5375_1 = ~Ng692 ^ ~n6110;
  assign n2177 = n5375_1 & n5106;
  assign n5377 = ~Ng1378 ^ ~n6088;
  assign n3696_1 = n5377 & n5109;
  assign n5379 = ~Ng2072 ^ ~n6066_1;
  assign n5190 = n5379 & n5112;
  assign n5381 = ~Ng2766 ^ ~n6044;
  assign n6697 = n5381 & n5115_1;
  assign n5383 = ~Ng61 ^ ~n6034;
  assign n1293_1 = n5383 & n5230_1;
  assign n5385_1 = ~Ng749 ^ ~n6030;
  assign n2799_1 = n5385_1 & n5230_1;
  assign n5387 = ~Ng1435 ^ ~n6026;
  assign n4306_1 = n5387 & n5230_1;
  assign n5389 = ~Ng2129 ^ ~n6022;
  assign n5800 = n5389 & n5230_1;
  assign n5391 = ~\[1612]  | n6530_1;
  assign n5392 = n4990 & ~n5663 & Ng2257;
  assign n1398_1 = n5391 & (Ng427 | (\[1612]  & n5392));
  assign n5394 = ~\[1594]  | n6530_1;
  assign n1403 = n5394 & (Ng428 | (\[1594]  & n5392));
  assign n5396 = ~\[1612]  | n6529;
  assign n5397 = n5002 & ~n5666 & Ng2257;
  assign n2904 = n5396 & (Ng1114 | (\[1612]  & n5397));
  assign n5399 = ~Ng853 | n6530_1;
  assign n1408_1 = n5399 & (Ng426 | (Ng853 & n5392));
  assign n5401 = ~\[1594]  | n6529;
  assign n2909_1 = n5401 & (Ng1115 | (\[1594]  & n5397));
  assign n5403 = ~\[1612]  | n6528;
  assign n5404 = n5014 & ~n5669 & Ng2257;
  assign n4411 = n5403 & (Ng1808 | (\[1612]  & n5404));
  assign n5406 = ~Ng853 | n6529;
  assign n2914_1 = n5406 & (Ng1113 | (Ng853 & n5397));
  assign n5408 = ~\[1594]  | n6528;
  assign n4416 = n5408 & (Ng1809 | (\[1594]  & n5404));
  assign n5410_1 = ~\[1612]  | n6527;
  assign n5411 = n5026 & ~n5672 & Ng2257;
  assign n5918 = n5410_1 & (Ng2502 | (\[1612]  & n5411));
  assign n5413 = ~Ng853 | n6528;
  assign n4421 = n5413 & (Ng1807 | (Ng853 & n5404));
  assign n5415_1 = ~\[1594]  | n6527;
  assign n5923 = n5415_1 & (Ng2503 | (\[1594]  & n5411));
  assign n5417 = ~Ng853 | n6527;
  assign n5928 = n5417 & (Ng2501 | (Ng853 & n5411));
  assign n5419 = ~n5971 ^ ~Ng56;
  assign n1298 = n5419 & n5230_1;
  assign n5421 = ~n5968_1 ^ ~Ng744;
  assign n2804_1 = n5421 & n5230_1;
  assign n5423 = ~n5965 ^ ~Ng1430;
  assign n4311_1 = n5423 & n5230_1;
  assign n5425_1 = ~n5962 ^ ~Ng2124;
  assign n5805 = n5425_1 & n5230_1;
  assign n5427 = ~Ng52 ^ ~n5972;
  assign n1303 = n5427 & n5230_1;
  assign n5429 = ~Ng740 ^ ~n5969;
  assign n2809_1 = n5429 & n5230_1;
  assign n5431 = ~Ng1426 ^ ~n5966;
  assign n4316 = n5431 & n5230_1;
  assign n5433 = ~Ng2120 ^ ~n5963_1;
  assign n5810 = n5433 & n5230_1;
  assign n5435_1 = n5542 | n5920;
  assign n5436 = n4585 | n6013_1;
  assign n5437 = n5435_1 & n5436 & (~n4958_1 | ~n5542);
  assign n5438 = n5544 | n5900;
  assign n5439 = n4593 | n6005;
  assign n5440_1 = n5438 & n5439 & (~n4966 | ~n5544);
  assign n5441 = n5546 | n5880;
  assign n5442 = n4603 | n5997;
  assign n5443 = n5441 & n5442 & (~n4974 | ~n5546);
  assign n5444 = n5548 | n5860;
  assign n5445_1 = n4615 | n5989;
  assign n5446 = n5444 & n5445_1 & (~n4980 | ~n5548);
  assign n5447 = n4672_1 ^ ~n5311;
  assign n5448 = ~n5030 & ~n5923_1;
  assign n5449 = (n5448 | ~n5828_1) & (n5447 | ~n5925);
  assign n5450_1 = ~n4684_1 ^ ~n6379;
  assign n5451 = Ng101 & ~n5923_1;
  assign n5452 = (n5451 | ~n5828_1) & (n5450_1 | ~n5925);
  assign n5453 = n4692_1 ^ ~n5314;
  assign n5454 = ~n5038_1 & ~n5903_1;
  assign n5455_1 = (n5454 | ~n5829) & (n5453 | ~n5905);
  assign n5456 = ~n4702 ^ ~n6378_1;
  assign n5457 = Ng109 & ~n5923_1;
  assign n5458 = (n5457 | ~n5828_1) & (n5456 | ~n5925);
  assign n5459 = ~n4708_1 ^ ~n6355;
  assign n5460_1 = Ng789 & ~n5903_1;
  assign n5461 = (n5460_1 | ~n5829) & (n5459 | ~n5905);
  assign n5462 = n4716_1 ^ ~n5317;
  assign n5463 = ~n5042 & ~n5883_1;
  assign n5464 = (n5463 | ~n5830) & (n5462 | ~n5885);
  assign n5465_1 = ~n4732_1 ^ ~n6354;
  assign n5466 = Ng797 & ~n5903_1;
  assign n5467 = (n5466 | ~n5829) & (n5465_1 | ~n5905);
  assign n5468 = ~n4738 ^ ~n6331_1;
  assign n5469 = Ng1476 & ~n5883_1;
  assign n5470_1 = (n5469 | ~n5830) & (n5468 | ~n5885);
  assign n5471 = n4746 ^ ~n5320_1;
  assign n5472 = ~n5046 & ~n5863_1;
  assign n5473 = (n5472 | ~n5831) & (n5471 | ~n5865);
  assign n5474 = ~n4768 ^ ~n6330;
  assign n5475_1 = Ng1486 & ~n5883_1;
  assign n5476 = (n5475_1 | ~n5830) & (n5474 | ~n5885);
  assign n5477 = ~n4774_1 ^ ~n6307;
  assign n5478 = Ng2170 & ~n5863_1;
  assign n5479 = (n5478 | ~n5831) & (n5477 | ~n5865);
  assign n5480_1 = n4782 ^ ~n5313;
  assign n5481 = ~n5020 & ~n5923_1;
  assign n5482 = (n5481 | ~n5828_1) & (n5480_1 | ~n5925);
  assign n5483 = ~n4810_1 ^ ~n6306;
  assign n5484 = Ng2180 & ~n5863_1;
  assign n5485_1 = (n5484 | ~n5831) & (n5483 | ~n5865);
  assign n5486 = ~n4814_1 ^ ~n6380;
  assign n5487 = Ng105 & ~n5923_1;
  assign n5488 = (n5487 | ~n5828_1) & (n5486 | ~n5925);
  assign n5489 = n4824_1 ^ ~n5316;
  assign n5490_1 = ~n5032 & ~n5903_1;
  assign n5491 = (n5490_1 | ~n5829) & (n5489 | ~n5905);
  assign n5492 = ~n4856_1 ^ ~n6356;
  assign n5493 = Ng793 & ~n5903_1;
  assign n5494 = (n5493 | ~n5829) & (n5492 | ~n5905);
  assign n5495_1 = n4866_1 ^ ~n5319;
  assign n5496 = ~n5040 & ~n5883_1;
  assign n5497 = (n5496 | ~n5830) & (n5495_1 | ~n5885);
  assign n5498 = ~n4894 ^ ~n6332;
  assign n5499 = Ng1481 & ~n5883_1;
  assign n5500_1 = (n5499 | ~n5830) & (n5498 | ~n5885);
  assign n5501 = n4904 ^ ~n5322;
  assign n5502 = ~n5044 & ~n5863_1;
  assign n5503 = (n5502 | ~n5831) & (n5501 | ~n5865);
  assign n5504 = ~n4924_1 ^ ~n6308_1;
  assign n5505_1 = Ng2175 & ~n5863_1;
  assign n5506 = (n5505_1 | ~n5831) & (n5504 | ~n5865);
  assign n5507 = ~n4854 | n4964;
  assign n5508 = ~n4964 & ~n5981;
  assign n5509 = n5507 & ~n5826 & (n4854 | n5508);
  assign n5510_1 = n5981 & n5054;
  assign n5511 = ~n5826 & (n5510_1 | ~n6981_1);
  assign n5512 = n5981 & n4964;
  assign n5513 = ~n5826 & (n5512 | ~n6982);
  assign n5514 = ~n4818 | n5054;
  assign n5515_1 = n5514 & ~n5826 & (n4818 | ~n8450);
  assign n5516 = ~n5826 & (n5510_1 | ~n6980);
  assign n5517 = ~n4686 | n4964;
  assign n5518 = n5517 & ~n5826 & (n4686 | n5508);
  assign n5519 = ~n4788 | n4964;
  assign n5520_1 = n5519 & ~n5826 & (n4788 | n5508);
  assign n5521 = ~n4886 | n5054;
  assign n5522 = n5521 & ~n5826 & (n4886 | ~n8450);
  assign n5523 = Pg563 | n5979 | Ng559 | ~n6600;
  assign n5524 = ~n6016 & (n5523 | (Ng8284 & ~n5825));
  assign n5525_1 = ~n4916 | n5058_1;
  assign n5526 = n5525_1 & ~n5823_1 & (n4916 | ~n8451);
  assign n5527 = ~n4892_1 | n4972;
  assign n5528 = ~n4972 & ~n5955;
  assign n5529 = n5527 & ~n5823_1 & (n4892_1 | n5528);
  assign n5530_1 = n5955 & n5058_1;
  assign n5531 = ~n5823_1 & (n5530_1 | ~n6951_1);
  assign n5532 = n5955 & n4972;
  assign n5533 = ~n5823_1 & (n5532 | ~n6952);
  assign n5534 = ~n4860 | n5058_1;
  assign n5535_1 = n5534 & ~n5823_1 & (n4860 | ~n8451);
  assign n5536 = ~n5823_1 & (n5530_1 | ~n6950);
  assign n5537 = ~n4710 | n4972;
  assign n5538 = n5537 & ~n5823_1 & (n4710 | n5528);
  assign n5539 = ~n4830 | n4972;
  assign n5540_1 = n5539 & ~n5823_1 & (n4830 | n5528);
  assign n5541 = (~n5911 & (n4958_1 | n6514)) | (~n4958_1 & n6514);
  assign n5542 = ~n4950 & ~n8584 & (n4954 | n5541);
  assign n5543 = (~n5891 & (n4966 | n6504)) | (~n4966 & n6504);
  assign n5544 = ~n4956 & ~n8583 & (n4960 | n5543);
  assign n5545_1 = (~n5871 & (n4974 | n6494)) | (~n4974 & n6494);
  assign n5546 = ~n4962 & ~n8582 & (n4968_1 | n5545_1);
  assign n5547 = (~n5851 & (n4980 | n6484)) | (~n4980 & n6484);
  assign n5548 = ~n4970 & ~n8581 & (n4976 | n5547);
  assign n5549 = ~n6601 | Pg1249 | Ng1245;
  assign n5550_1 = ~n5958_1 & (n5549 | (Ng8293 & ~n5822));
  assign n5551 = ~n5914 & (~n4958_1 | n5908_1 | ~n6514);
  assign n5552 = ~n4950 & ~n8577 & (n4954 | n5551);
  assign n5553 = ~n5894 & (~n4966 | n5888_1 | ~n6504);
  assign n5554 = ~n4956 & ~n8572 & (n4960 | n5553);
  assign n5555_1 = ~n5874 & (~n4974 | n5868_1 | ~n6494);
  assign n5556 = ~n4962 & ~n8567 & (n4968_1 | n5555_1);
  assign n5557 = ~n5854 & (~n4980 | n5848_1 | ~n6484);
  assign n5558 = ~n4970 & ~n8562 & (n4976 | n5557);
  assign n5559 = (~n4872 & n8452) | (n4978_1 & (n4872 | n8452));
  assign n5560_1 = n5559 & ~n5820;
  assign n5561 = (~n4936 & ~n8453) | (n5062 & (n4936 | ~n8453));
  assign n5562 = n5561 & ~n5820;
  assign n5563 = (~n4922 & n8452) | (n4978_1 & (n4922 | n8452));
  assign n5564 = n5563 & ~n5820;
  assign n5565_1 = n5062 & ~n5840;
  assign n5566 = ~n5820 & (n5565_1 | ~n6617_1);
  assign n5567 = n4978_1 & ~n5840;
  assign n5568 = ~n5820 & (n5567 | ~n6618);
  assign n5569 = (~n4898 & ~n8453) | (n5062 & (n4898 | ~n8453));
  assign n5570_1 = n5569 & ~n5820;
  assign n5571 = ~n5820 & (n5565_1 | ~n6616);
  assign n5572 = (~n4740 & n8452) | (n4978_1 & (n4740 | n8452));
  assign n5573 = n5572 & ~n5820;
  assign n5574 = ~n6602_1 | Pg1943 | Ng1939;
  assign n5575_1 = ~n5843_1 & (n5574 | (Ng8302 & ~n5819_1));
  assign n5576 = n5591 | ~Ng8311;
  assign n5577 = n5576 | ~n8554;
  assign n5578 = (~n4910_1 & n8454) | (n4982 & (n4910_1 | n8454));
  assign n5579 = ~n5576 & n5578;
  assign n5580_1 = (~n4948_1 & ~n8455) | (n5064 & (n4948_1 | ~n8455));
  assign n5581 = ~n5576 & n5580_1;
  assign n5582 = (~n4942 & n8454) | (n4982 & (n4942 | n8454));
  assign n5583 = ~n5576 & n5582;
  assign n5584 = n5064 & ~n5833_1;
  assign n5585_1 = ~n5576 & (n5584 | ~n6606);
  assign n5586 = n4982 & ~n5833_1;
  assign n5587 = ~n5576 & (n5586 | ~n6607_1);
  assign n5588 = (~n4928_1 & ~n8455) | (n5064 & (n4928_1 | ~n8455));
  assign n5589 = ~n5576 & n5588;
  assign n5590_1 = ~n5576 & (n5584 | ~n6605);
  assign n5591 = ~n6603 | Pg2637 | Ng2633;
  assign n5592 = ~n5836 & (n5591 | (Ng8311 & ~n5817));
  assign n5593 = Ng2874 ^ ~Ng2981;
  assign n5594 = Ng2978 ^ ~Ng2975;
  assign n5595_1 = ~Ng2874 ^ ~Ng2981;
  assign n5596 = ~Ng2978 ^ ~Ng2975;
  assign n5597 = (n5593 | n5594) & (n5595_1 | n5596);
  assign n5598 = Ng2972 ^ ~Ng2969;
  assign n5599 = Ng2966 ^ ~Ng2963;
  assign n5600_1 = ~Ng2972 ^ ~Ng2969;
  assign n5601 = ~Ng2966 ^ ~Ng2963;
  assign n5602 = (n5598 | n5599) & (n5600_1 | n5601);
  assign n5603 = Ng2959 ^ ~Ng2956;
  assign n5604 = Ng2953 ^ ~Ng2947;
  assign n5605_1 = ~Ng2959 ^ ~Ng2956;
  assign n5606 = ~Ng2953 ^ ~Ng2947;
  assign n5607 = (n5603 | n5604) & (n5605_1 | n5606);
  assign n5608 = Ng2944 ^ ~Ng2941;
  assign n5609 = Ng2938 ^ ~Ng2935;
  assign n5610_1 = ~Ng2944 ^ ~Ng2941;
  assign n5611 = ~Ng2938 ^ ~Ng2935;
  assign n5612 = (n5608 | n5609) & (n5610_1 | n5611);
  assign n5613 = ~n5826 & (n5512 | ~n6978);
  assign n5614 = ~n5826 & (n5510_1 | ~n6979);
  assign n5615_1 = n5509 ^ ~n5522;
  assign n5616 = n5515_1 ^ ~n5520_1;
  assign n5617 = ~n5509 ^ ~n5522;
  assign n5618 = ~n5515_1 ^ ~n5520_1;
  assign n5619 = (n5615_1 | n5616) & (n5617 | n5618);
  assign n5620_1 = n5516 ^ ~n5518;
  assign n5621 = n5511 ^ ~n5513;
  assign n5622 = ~n5516 ^ ~n5518;
  assign n5623 = ~n5511 ^ ~n5513;
  assign n5624 = (n5620_1 | n5621) & (n5622 | n5623);
  assign n5625_1 = ~n5823_1 & (n5532 | ~n6948);
  assign n5626 = ~n5823_1 & (n5530_1 | ~n6949);
  assign n5627 = n5535_1 ^ ~n5540_1;
  assign n5628 = n5526 ^ ~n5529;
  assign n5629 = ~n5535_1 ^ ~n5540_1;
  assign n5630_1 = ~n5526 ^ ~n5529;
  assign n5631 = (n5627 | n5628) & (n5629 | n5630_1);
  assign n5632 = n5536 ^ ~n5538;
  assign n5633 = n5531 ^ ~n5533;
  assign n5634 = ~n5536 ^ ~n5538;
  assign n5635_1 = ~n5531 ^ ~n5533;
  assign n5636 = (n5632 | n5633) & (n5634 | n5635_1);
  assign n5637 = ~n5820 & (n5567 | ~n6614);
  assign n5638 = ~n5820 & (n5565_1 | ~n6615);
  assign n5639 = n5560_1 ^ ~n5570_1;
  assign n5640_1 = n5562 ^ ~n5564;
  assign n5641 = ~n5560_1 ^ ~n5570_1;
  assign n5642 = ~n5562 ^ ~n5564;
  assign n5643 = (n5639 | n5640_1) & (n5641 | n5642);
  assign n5644 = n5571 ^ ~n5573;
  assign n5645_1 = n5566 ^ ~n5568;
  assign n5646 = ~n5571 ^ ~n5573;
  assign n5647 = ~n5566 ^ ~n5568;
  assign n5648 = (n5644 | n5645_1) & (n5646 | n5647);
  assign n5649 = ~n5576 & (n5586 | ~n6599);
  assign n5650_1 = ~n5576 & (n5584 | ~n6604);
  assign n5651 = n5579 ^ ~n5589;
  assign n5652 = n5581 ^ ~n5583;
  assign n5653 = ~n5579 ^ ~n5589;
  assign n5654 = ~n5581 ^ ~n5583;
  assign n5655_1 = (n5651 | n5652) & (n5653 | n5654);
  assign n5656 = ~n5590_1 ^ ~n5577;
  assign n5657 = n5585_1 ^ ~n5587;
  assign n5658 = n5577 ^ ~n5590_1;
  assign n5659 = ~n5585_1 ^ ~n5587;
  assign n5660_1 = (n5656 | n5657) & (n5658 | n5659);
  assign n5661 = n6515_1 | ~n4998_1 | ~n5662;
  assign n5662 = n6170 & ~n5020 & ~n5030;
  assign n5663 = n5661 & (n5662 | n4998_1);
  assign n5664 = n6505_1 | ~n5010 | ~n5665_1;
  assign n5665_1 = n6163_1 & ~n5032 & ~n5038_1;
  assign n5666 = n5664 & (n5665_1 | n5010);
  assign n5667 = n6495_1 | ~n5022 | ~n5668;
  assign n5668 = n6156 & ~n5040 & ~n5042;
  assign n5669 = n5667 & (n5668 | n5022);
  assign n5670_1 = n6485_1 | ~n5034 | ~n5671;
  assign n5671 = n6149 & ~n5044 & ~n5046;
  assign n5672 = n5670_1 & (n5671 | n5034);
  assign n6133 = ~n5034;
  assign n4626 = ~n5022;
  assign n3119_1 = ~n5010;
  assign n1613 = ~n4998_1;
  assign n5677 = n5834 & (~Ng2584 | n5835);
  assign n7101 = ~n5677;
  assign n5679 = (~n5071 | ~n8458) & (n5649 | n5836);
  assign n7096 = ~n5679;
  assign n5681 = (~n5071 | ~n8459) & (n5650_1 | n5836);
  assign n7091 = ~n5681;
  assign n5683 = n5837 & (~n5071 | ~n8460);
  assign n7086 = ~n5683;
  assign n5685_1 = n5837 & (~n5071 | ~n8461);
  assign n7081 = ~n5685_1;
  assign n5687 = ~n5818 & (~n5071 | ~n8462);
  assign n7076 = ~n5687;
  assign n5689 = ~n5592 & (~n5071 | ~n8463);
  assign n7071 = ~n5689;
  assign n5691 = ~n5592 & (~n5071 | ~n8464);
  assign n7066 = ~n5691;
  assign n5693 = ~n5818 & (~n5071 | ~n8465);
  assign n7061 = ~n5693;
  assign n5695_1 = n5841 & (~Ng1890 | n5842);
  assign n7056 = ~n5695_1;
  assign n5697 = (~n5069 | ~n8468) & (n5637 | n5843_1);
  assign n7051 = ~n5697;
  assign n5699 = (~n5069 | ~n8469) & (n5638 | n5843_1);
  assign n7046 = ~n5699;
  assign n5701 = n5844 & (~n5069 | ~n8470);
  assign n7041 = ~n5701;
  assign n5703 = n5844 & (~n5069 | ~n8471);
  assign n7036 = ~n5703;
  assign n5705_1 = ~n5821 & (~n5069 | ~n8472);
  assign n7031 = ~n5705_1;
  assign n5707 = ~n5575_1 & (~n5069 | ~n8473);
  assign n7026 = ~n5707;
  assign n5709 = ~n5575_1 & (~n5069 | ~n8474);
  assign n7021 = ~n5709;
  assign n5711 = ~n5821 & (~n5069 | ~n8475);
  assign n7016 = ~n5711;
  assign n5713 = n5956 & (~Ng1196 | n5957);
  assign n7011 = ~n5713;
  assign n5715_1 = (~n5067_1 | ~n8502) & (n5625_1 | n5958_1);
  assign n7006 = ~n5715_1;
  assign n5717 = (~n5067_1 | ~n8503) & (n5626 | n5958_1);
  assign n7001 = ~n5717;
  assign n5719 = n5959 & (~n5067_1 | ~n8504);
  assign n6996 = ~n5719;
  assign n5721 = n5959 & (~n5067_1 | ~n8505);
  assign n6991 = ~n5721;
  assign n5723 = ~n5824 & (~n5067_1 | ~n8506);
  assign n6986 = ~n5723;
  assign n5725_1 = ~n5550_1 & (~n5067_1 | ~n8507);
  assign n6981 = ~n5725_1;
  assign n5727 = ~n5550_1 & (~n5067_1 | ~n8508);
  assign n6976 = ~n5727;
  assign n5729 = ~n5824 & (~n5067_1 | ~n8509);
  assign n6971 = ~n5729;
  assign n5731 = n5982 & (~Ng510 | n5983_1);
  assign n6966 = ~n5731;
  assign n5733 = (~n5065 | ~n8512) & (n5613 | n6016);
  assign n6961 = ~n5733;
  assign n5735_1 = (~n5065 | ~n8513) & (n5614 | n6016);
  assign n6956 = ~n5735_1;
  assign n5737 = n6017 & (~n5065 | ~n8514);
  assign n6951 = ~n5737;
  assign n5739 = n6017 & (~n5065 | ~n8515);
  assign n6946 = ~n5739;
  assign n5741 = ~n5827 & (~n5065 | ~n8516);
  assign n6941 = ~n5741;
  assign n5743 = ~n5524 & (~n5065 | ~n8517);
  assign n6936 = ~n5743;
  assign n5745_1 = ~n5524 & (~n5065 | ~n8518);
  assign n6931 = ~n5745_1;
  assign n5747 = ~n5827 & (~n5065 | ~n8519);
  assign n6926 = ~n5747;
  assign n6637 = ~Ng2366;
  assign n6627 = ~Ng2364;
  assign n6622 = ~Ng2362;
  assign n6617 = ~Ng2360;
  assign n6612 = ~Ng2358;
  assign n6607 = ~Ng2356;
  assign n6602 = ~Ng2354;
  assign n6597 = ~Ng2528;
  assign n6592 = ~Ng2526;
  assign n6116 = ~Ng2165;
  assign n6107 = ~Ng2170;
  assign n6098 = ~Ng2175;
  assign n6089 = ~Ng2180;
  assign n6080 = ~Ng2185;
  assign n6071 = ~Ng2190;
  assign n6062 = ~Ng2195;
  assign n6053 = ~Ng2200;
  assign n5130 = ~Ng1672;
  assign n5120 = ~Ng1670;
  assign n5115 = ~Ng1668;
  assign n5110 = ~Ng1666;
  assign n5105 = ~Ng1664;
  assign n5100 = ~Ng1662;
  assign n5095 = ~Ng1660;
  assign n5090 = ~Ng1834;
  assign n5085 = ~Ng1832;
  assign n4609 = ~Ng1471;
  assign n4600 = ~Ng1476;
  assign n4591 = ~Ng1481;
  assign n4582 = ~Ng1486;
  assign n4573 = ~Ng1491;
  assign n4564 = ~Ng1496;
  assign n4555 = ~Ng1501;
  assign n4546 = ~Ng1506;
  assign n3623_1 = ~Ng978;
  assign n3613_1 = ~Ng976;
  assign n3608_1 = ~Ng974;
  assign n3603_1 = ~Ng972;
  assign n3598_1 = ~Ng970;
  assign n3593_1 = ~Ng968;
  assign n3588_1 = ~Ng966;
  assign n3583_1 = ~Ng1140;
  assign n3578_1 = ~Ng1138;
  assign n3102 = ~Ng785;
  assign n3093_1 = ~Ng789;
  assign n3084_1 = ~Ng793;
  assign n3075 = ~Ng797;
  assign n3066_1 = ~Ng801;
  assign n3057_1 = ~Ng805;
  assign n3048_1 = ~Ng809;
  assign n3039_1 = ~Ng813;
  assign n2117_1 = ~Ng291;
  assign n2107_1 = ~Ng289;
  assign n2102_1 = ~Ng287;
  assign n2097_1 = ~Ng285;
  assign n2092_1 = ~Ng283;
  assign n2087_1 = ~Ng281;
  assign n2082 = ~Ng279;
  assign n2077_1 = ~Ng453;
  assign n2072_1 = ~Ng451;
  assign n1596 = ~Ng97;
  assign n1587 = ~Ng101;
  assign n1578 = ~Ng105;
  assign n1569_1 = ~Ng109;
  assign n1560_1 = ~Ng113;
  assign n1551_1 = ~Ng117;
  assign n1542_1 = ~Ng121;
  assign n1533_1 = ~Ng125;
  assign n5817 = n5833_1 & n5838_1 & (~\[1605]  | Ng2809);
  assign n5818 = ~n5836 & (n5576 | n5817);
  assign n5819_1 = n5840 & n5845 & (~\[1605]  | Ng2115);
  assign n5820 = n5574 | ~Ng8302;
  assign n5821 = ~n5843_1 & (n5819_1 | n5820);
  assign n5822 = ~n5955 & n5960 & (~\[1605]  | Ng1421);
  assign n5823_1 = n5549 | ~Ng8293;
  assign n5824 = ~n5958_1 & (n5822 | n5823_1);
  assign n5825 = ~n5981 & n6018_1 & (~\[1605]  | Ng735);
  assign n5826 = n5523 | ~Ng8284;
  assign n5827 = ~n6016 & (n5825 | n5826);
  assign n5828_1 = ~n5925 & (~n5923_1 | ~n5947);
  assign n5829 = ~n5905 & (~n5903_1 | ~n5940);
  assign n5830 = ~n5885 & (~n5883_1 | ~n5933_1);
  assign n5831 = ~n5865 & (~n5863_1 | ~n5926);
  assign n5832 = n4952 | n4930 | n4882 | n4812 | n4778_1 | n4848;
  assign n5833_1 = ~n4928_1 | ~n4776 | ~n4910_1 | ~n8457 | ~n4942 | n5832;
  assign n5834 = (~Ng2631 | n8556) & n8557;
  assign n5835 = n5655_1 ^ ~n5660_1;
  assign n5836 = n5071 | ~n5072_1;
  assign n5837 = ~n5591 | n5836;
  assign n5838_1 = (~Ng1315 | Ng2808) & (~\[1603]  | Ng2810);
  assign n5839 = n4944 | n4900 | n4840 | n4770 | n4742_1 | n4806;
  assign n5840 = ~n4898 | ~n4740 | ~n4872 | ~n8467 | ~n4922 | n5839;
  assign n5841 = (~Ng1937 | n8559) & n8560;
  assign n5842 = n5643 ^ ~n5648;
  assign n5843_1 = n5069 | ~n5070;
  assign n5844 = ~n5574 | n5843_1;
  assign n5845 = (~Ng1315 | Ng2114) & (~\[1603]  | Ng2116);
  assign n5846 = (n6297 | ~n6298) & (n6299_1 | n6300);
  assign n5847 = n4846_1 ^ ~Ng2190;
  assign n5848_1 = ~n5849 & (~n8481 | (n5846 & n5847));
  assign n5849 = n4946 | ~Ng2257;
  assign n5850 = n6300 | n6482 | ~n6298 | n6299_1 | n5847 | n5853_1 | n6296 | n6297;
  assign n5851 = ~n6485_1 & (n5849 | n5850);
  assign n5852 = (n6293 | n6294_1) & (n6295 | n6296);
  assign n5853_1 = ~n4746 ^ ~n5046;
  assign n5854 = ~n5849 & (~n8478 | (n5852 & n5853_1));
  assign n5855 = n6301 & ~n6308_1 & ~n6488;
  assign n5856 = n5855 & (n4846_1 | ~n5926);
  assign n5857 = n4720_1 ^ ~n5926;
  assign n5858_1 = (n4876_1 & n5926) | (~n4846_1 & (~n4876_1 | n5926));
  assign n5859 = ~n5989 & ~n6483;
  assign n5860 = ~n4970 & n4980;
  assign n5861 = n5860 & n4976 & n5859;
  assign n5862 = ~n4643 & (n5861 | (~n5989 & ~n5990));
  assign n5863_1 = n5445_1 & ~n5862 & (n4970 | ~n6485_1);
  assign n5864 = n6219_1 & n5926;
  assign n5865 = n5863_1 & (n5864 | ~n6626);
  assign n5866 = (n6321_1 | ~n6322) & (n6323 | n6324);
  assign n5867 = n4804 ^ ~Ng1496;
  assign n5868_1 = ~n5869 & (~n8487 | (n5866 & n5867));
  assign n5869 = n4934 | ~Ng2257;
  assign n5870 = n6324 | n6492 | ~n6322 | n6323 | n5867 | n5873_1 | n6320 | n6321_1;
  assign n5871 = ~n6495_1 & (n5869 | n5870);
  assign n5872 = (n6317_1 | n6318) & (n6319 | n6320);
  assign n5873_1 = ~n4716_1 ^ ~n5042;
  assign n5874 = ~n5869 & (~n8484 | (n5872 & n5873_1));
  assign n5875 = n6325 & ~n6332 & ~n6498;
  assign n5876 = n5875 & (n4804 | ~n5933_1);
  assign n5877 = n4696_1 ^ ~n5933_1;
  assign n5878_1 = (n4834_1 & n5933_1) | (~n4804 & (~n4834_1 | n5933_1));
  assign n5879 = ~n5997 & ~n6493;
  assign n5880 = ~n4962 & n4974;
  assign n5881 = n5880 & n4968_1 & n5879;
  assign n5882 = ~n4639 & (n5881 | (~n5997 & ~n5998_1));
  assign n5883_1 = n5442 & ~n5882 & (n4962 | ~n6495_1);
  assign n5884 = n6223_1 & n5933_1;
  assign n5885 = n5883_1 & (n5884 | ~n6664);
  assign n5886 = (n6345_1 | ~n6346) & (n6347 | n6348);
  assign n5887 = n4762 ^ ~Ng805;
  assign n5888_1 = ~n5889 & (~n8493 | (n5886 & n5887));
  assign n5889 = n4914 | ~Ng2257;
  assign n5890 = n6348 | n6502 | ~n6346 | n6347 | n5887 | n5893_1 | n6344 | n6345_1;
  assign n5891 = ~n6505_1 & (n5889 | n5890);
  assign n5892 = (n6341_1 | n6342) & (n6343 | n6344);
  assign n5893_1 = ~n4692_1 ^ ~n5038_1;
  assign n5894 = ~n5889 & (~n8490 | (n5892 & n5893_1));
  assign n5895 = n6349_1 & ~n6356 & ~n6508;
  assign n5896 = n5895 & (n4762 | ~n5940);
  assign n5897 = n4676_1 ^ ~n5940;
  assign n5898_1 = (n4792_1 & n5940) | (~n4762 & (~n4792_1 | n5940));
  assign n5899 = ~n6005 & ~n6503;
  assign n5900 = ~n4956 & n4966;
  assign n5901 = n5900 & n4960 & n5899;
  assign n5902 = ~n4633 & (n5901 | (~n6005 & ~n6006));
  assign n5903_1 = n5439 & ~n5902 & (n4956 | ~n6505_1);
  assign n5904 = n6227_1 & n5940;
  assign n5905 = n5903_1 & (n5904 | ~n6702_1);
  assign n5906 = (n6369 | ~n6370) & (n6371 | n6372);
  assign n5907 = n4726 ^ ~Ng117;
  assign n5908_1 = ~n5909 & (~n8499 | (n5906 & n5907));
  assign n5909 = n4884_1 | ~Ng2257;
  assign n5910 = n6372 | n6512 | ~n6370 | n6371 | n5907 | n5913_1 | n6368_1 | n6369;
  assign n5911 = ~n6515_1 & (n5909 | n5910);
  assign n5912 = (n6365 | n6366) & (n6367 | n6368_1);
  assign n5913_1 = ~n4672_1 ^ ~n5030;
  assign n5914 = ~n5909 & (~n8496 | (n5912 & n5913_1));
  assign n5915 = n6373_1 & ~n6380 & ~n6518;
  assign n5916 = n5915 & (n4726 | ~n5947);
  assign n5917 = n4662 ^ ~n5947;
  assign n5918_1 = (n4750 & n5947) | (~n4726 & (~n4750 | n5947));
  assign n5919 = ~n6013_1 & ~n6513;
  assign n5920 = ~n4950 & n4958_1;
  assign n5921 = n5920 & n4954 & n5919;
  assign n5922 = ~n4625 & (n5921 | (~n6013_1 & ~n6014));
  assign n5923_1 = n5436 & ~n5922 & (n4950 | ~n6515_1);
  assign n5924 = n6231_1 & n5947;
  assign n5925 = n5923_1 & (n5924 | ~n6740);
  assign n5926 = ~n4970 | n4976 | ~n4980;
  assign n5927 = n5856 & (~n4846_1 | n5926);
  assign n5928_1 = n5927 & n5857;
  assign n5929 = Ng2200 & ~n5863_1;
  assign n5930 = Ng2195 & ~n5863_1;
  assign n5931 = Ng2185 & ~n5863_1;
  assign n5932 = Ng2165 & ~n5863_1;
  assign n5933_1 = ~n4962 | n4968_1 | ~n4974;
  assign n5934 = n5876 & (~n4804 | n5933_1);
  assign n5935 = n5934 & n5877;
  assign n5936 = Ng1506 & ~n5883_1;
  assign n5937 = Ng1501 & ~n5883_1;
  assign n5938_1 = Ng1491 & ~n5883_1;
  assign n5939 = Ng1471 & ~n5883_1;
  assign n5940 = ~n4956 | n4960 | ~n4966;
  assign n5941 = n5896 & (~n4762 | n5940);
  assign n5942 = n5941 & n5897;
  assign n5943_1 = Ng813 & ~n5903_1;
  assign n5944 = Ng809 & ~n5903_1;
  assign n5945 = Ng801 & ~n5903_1;
  assign n5946 = Ng785 & ~n5903_1;
  assign n5947 = ~n4950 | n4954 | ~n4958_1;
  assign n5948_1 = n5916 & (~n4726 | n5947);
  assign n5949 = n5948_1 & n5917;
  assign n5950 = Ng125 & ~n5923_1;
  assign n5951 = Ng121 & ~n5923_1;
  assign n5952 = Ng113 & ~n5923_1;
  assign n5953_1 = Ng97 & ~n5923_1;
  assign n5954 = n4916 & (~n8500 | (\[1603]  & ~Ng1425));
  assign n5955 = n5954 & n4892_1 & n4860 & n4710 & n4830 & ~n8501;
  assign n5956 = (~Ng1243 | n8612) & n8613;
  assign n5957 = n5631 ^ ~n5636;
  assign n5958_1 = n5067_1 | ~n5068;
  assign n5959 = ~n5549 | n5958_1;
  assign n5960 = (~Ng1315 | Ng1420) & (~\[1603]  | Ng1422);
  assign n5961 = n5926 & (n4970 | ~n5990 | ~n6483);
  assign n5962 = n6021 & Ng2133 & Ng2129;
  assign n5963_1 = n5962 & Ng2124;
  assign n5964 = n5933_1 & (n4962 | ~n5998_1 | ~n6493);
  assign n5965 = n6025 & Ng1439 & Ng1435;
  assign n5966 = n5965 & Ng1430;
  assign n5967 = n5940 & (n4956 | ~n6006 | ~n6503);
  assign n5968_1 = n6029 & Ng753 & Ng749;
  assign n5969 = n5968_1 & Ng744;
  assign n5970 = n5947 & (n4950 | ~n6014 | ~n6513);
  assign n5971 = n6033_1 & Ng65 & Ng61;
  assign n5972 = n5971 & Ng56;
  assign n5973_1 = n6522 | n5975;
  assign n5974 = ~Ng3135 | n6524;
  assign n5975 = ~Ng3147 | n6131;
  assign n5976 = n5973_1 & (n5974 | n5975);
  assign n5977 = n6531 & (Ng3120 | ~Ng3135 | ~n6977);
  assign n5978_1 = n5974 | Ng3147 | n6131;
  assign n5979 = \[1605]  & ~Ng8284;
  assign n5980 = n4886 & (~n8510 | (\[1603]  & ~Ng739));
  assign n5981 = n5980 & n4854 & n4818 & n4686 & n4788 & ~n8511;
  assign n5982 = (~Ng557 | n8619) & n8620;
  assign n5983_1 = n5619 ^ ~n5624;
  assign n5984 = ~n5034 | ~n5671 | ~Ng2257 | ~n6485_1;
  assign n5985 = n5034 & (n5060 | ~n5671);
  assign n5986 = ~n5034 & (n5060 | n5671);
  assign n5987 = n5026 | ~Ng2257;
  assign n5988_1 = n5984 & (n5985 | n5986 | n5987);
  assign n5989 = n5849 | n6291 | n6292 | n6479 | n6480_1 | n6481;
  assign n5990 = n4970 | ~n4976 | n4980;
  assign n5991 = (~n5859 | ~n5860) & (n5989 | n5990);
  assign n5992 = ~n5022 | ~n5668 | ~Ng2257 | ~n6495_1;
  assign n5993_1 = n5022 & (n5056 | ~n5668);
  assign n5994 = ~n5022 & (n5056 | n5668);
  assign n5995 = n5014 | ~Ng2257;
  assign n5996 = n5992 & (n5993_1 | n5994 | n5995);
  assign n5997 = n5869 | n6315 | n6316 | n6489 | n6490_1 | n6491;
  assign n5998_1 = n4962 | ~n4968_1 | n4974;
  assign n5999 = (~n5879 | ~n5880) & (n5997 | n5998_1);
  assign n6000 = ~n5010 | ~n5665_1 | ~Ng2257 | ~n6505_1;
  assign n6001 = n5010 & (n5052 | ~n5665_1);
  assign n6002 = ~n5010 & (n5052 | n5665_1);
  assign n6003_1 = n5002 | ~Ng2257;
  assign n6004 = n6000 & (n6001 | n6002 | n6003_1);
  assign n6005 = n5889 | n6339 | n6340 | n6499 | n6500_1 | n6501;
  assign n6006 = n4956 | ~n4960 | n4966;
  assign n6007 = (~n5899 | ~n5900) & (n6005 | n6006);
  assign n6008_1 = ~n4998_1 | ~n5662 | ~Ng2257 | ~n6515_1;
  assign n6009 = n4998_1 & (n5050 | ~n5662);
  assign n6010 = ~n4998_1 & (n5050 | n5662);
  assign n6011 = n4990 | ~Ng2257;
  assign n6012 = n6008_1 & (n6009 | n6010 | n6011);
  assign n6013_1 = n5909 | n6363_1 | n6364 | n6509 | n6510_1 | n6511;
  assign n6014 = n4950 | ~n4954 | n4958_1;
  assign n6015 = (~n5919 | ~n5920) & (n6013_1 | n6014);
  assign n6016 = n5065 | ~n5066;
  assign n6017 = ~n5523 | n6016;
  assign n6018_1 = (~Ng1315 | Ng734) & (~\[1603]  | Ng736);
  assign n6019 = n5034 | ~n5060 | n5671;
  assign n6020 = ~n5987 & (~n5060 | n5670_1) & n6019;
  assign n6021 = n6154 & Ng2142 & Ng2138;
  assign n6022 = n6021 & Ng2133;
  assign n6023_1 = n5022 | ~n5056 | n5668;
  assign n6024 = ~n5995 & (~n5056 | n5667) & n6023_1;
  assign n6025 = n6161 & Ng1448 & Ng1444;
  assign n6026 = n6025 & Ng1439;
  assign n6027 = n5010 | ~n5052 | n5665_1;
  assign n6028_1 = ~n6003_1 & (~n5052 | n5664) & n6027;
  assign n6029 = n6168 & Ng762 & Ng758;
  assign n6030 = n6029 & Ng753;
  assign n6031 = n4998_1 | ~n5050 | n5662;
  assign n6032 = ~n6011 & (~n5050 | n5661) & n6031;
  assign n6033_1 = n6175_1 & Ng74 & Ng70;
  assign n6034 = n6033_1 & Ng65;
  assign n6035 = ~n858_1 & n5976;
  assign n6036 = (~Ng3105 | n6549) & (n5978_1 | Ng3128);
  assign n6037 = (~Ng3103 | n6547) & (~Ng3104 | n6548);
  assign n6038_1 = (n6545_1 | ~Ng3101) & (n6546 | ~Ng3102);
  assign n6039 = (n6542 | ~Ng3099) & (n6543 | ~Ng3100);
  assign n6040 = (n6540_1 | ~Ng3097) & (n6541 | ~Ng3098);
  assign n6041 = (~Ng3107 | n6536) & (~Ng3108 | n6538);
  assign n6042 = (~Ng3106 | n6535_1) & (n6531 | ~n8756);
  assign n6043_1 = Ng2753 & n6550_1;
  assign n6044 = Ng2760 & n6043_1;
  assign n6045 = (~n4573_1 | ~n5028_1) & (n4567 | ~n5008_1);
  assign n6046 = n5008_1 & (~n8522 | (n4571 & ~n5028_1));
  assign n6047 = n4573_1 & (~n8521 | (n4567 & ~n5018_1));
  assign n6048_1 = n5028_1 & n5018_1;
  assign n6049 = ~n5008_1 & (n6047 | (n4561 & n6048_1));
  assign n6050 = ~n4573_1 & (n6046 | (~n5036 & ~n6057_1));
  assign n6051 = ~n5028_1 | n4561 | n4571;
  assign n6052 = n6051 & (~n4567 | (n4571 & ~n5028_1));
  assign n6053_1 = n5028_1 & (n4573_1 | ~n5036);
  assign n6054 = n4567 & (~n5036 | (~n4571 & n6048_1));
  assign n6055 = ~n6054 & (n4561 | n5008_1 | n5036);
  assign n6056 = (~n5018_1 & (n4573_1 | n5028_1)) | (~n4573_1 & n5028_1);
  assign n6057_1 = n4567 | n4571;
  assign n6058 = (~n4561 | n6053_1) & (n6056 | n6057_1);
  assign n6059 = n4573_1 | n5018_1 | n6052;
  assign n6060 = (~n5008_1 & ~n7061_1) | (n6058 & (n5008_1 | ~n7061_1));
  assign n6061 = n6059 & (~n4573_1 | n6055) & n6060;
  assign n6062_1 = n6395 | ~Ng185 | ~Ng2616;
  assign n6063 = (~\[1603]  | ~Ng2673) & (~\[1605]  | ~Ng2670);
  assign n6064 = n6062_1 & n6063 & (~Ng1315 | ~Ng2676);
  assign n6065 = Ng2059 & n6556;
  assign n6066_1 = Ng2066 & n6065;
  assign n6067 = (~n4569 | ~n5016) & (n4559_1 | ~n4996);
  assign n6068 = n4996 & (~n8525 | (n4565 & ~n5016));
  assign n6069 = n4569 & (~n8524 | (n4559_1 & ~n5006));
  assign n6070 = n5016 & n5006;
  assign n6071_1 = ~n4996 & (n6069 | (n4553 & n6070));
  assign n6072 = ~n4569 & (n6068 | (~n5024 & ~n6079));
  assign n6073 = ~n5016 | n4553 | n4565;
  assign n6074 = n6073 & (~n4559_1 | (n4565 & ~n5016));
  assign n6075_1 = n5016 & (n4569 | ~n5024);
  assign n6076 = n4559_1 & (~n5024 | (~n4565 & n6070));
  assign n6077 = ~n6076 & (n4553 | n4996 | n5024);
  assign n6078 = (~n5006 & (n4569 | n5016)) | (~n4569 & n5016);
  assign n6079 = n4559_1 | n4565;
  assign n6080_1 = (~n4553 | n6075_1) & (n6078 | n6079);
  assign n6081 = n4569 | n5006 | n6074;
  assign n6082 = (~n4996 & ~n7077) | (n6080_1 & (n4996 | ~n7077));
  assign n6083 = n6081 & (~n4569 | n6077) & n6082;
  assign n6084_1 = n4888 | ~Ng185 | ~Ng1922;
  assign n6085 = (~\[1603]  | ~Ng1979) & (~\[1605]  | ~Ng1976);
  assign n6086 = n6084_1 & n6085 & (~Ng1315 | ~Ng1982);
  assign n6087 = Ng1365 & n6560_1;
  assign n6088 = Ng1372 & n6087;
  assign n6089_1 = (~n4563 | ~n5004) & (n4551 | ~n4988_1);
  assign n6090 = n4988_1 & (~n8528 | (n4557 & ~n5004));
  assign n6091 = n4563 & (~n8527 | (n4551 & ~n4994));
  assign n6092 = n5004 & n4994;
  assign n6093_1 = ~n4988_1 & (n6091 | (n4547 & n6092));
  assign n6094 = ~n4563 & (n6090 | (~n5012 & ~n6101));
  assign n6095 = ~n5004 | n4547 | n4557;
  assign n6096 = n6095 & (~n4551 | (n4557 & ~n5004));
  assign n6097 = n5004 & (n4563 | ~n5012);
  assign n6098_1 = n4551 & (~n5012 | (~n4557 & n6092));
  assign n6099 = ~n6098_1 & (n4547 | n4988_1 | n5012);
  assign n6100 = (~n4994 & (n4563 | n5004)) | (~n4563 & n5004);
  assign n6101 = n4551 | n4557;
  assign n6102_1 = (~n4547 | n6097) & (n6100 | n6101);
  assign n6103 = n4563 | n4994 | n6096;
  assign n6104 = (~n4988_1 & ~n7093) | (n6102_1 & (n4988_1 | ~n7093));
  assign n6105 = n6103 & (~n4563 | n6099) & n6104;
  assign n6106 = n3381_1 | ~Ng185 | ~Ng1228;
  assign n6107_1 = (~\[1603]  | ~Ng1285) & (~\[1605]  | ~Ng1282);
  assign n6108 = n6106 & n6107_1 & (~Ng1315 | ~Ng1288);
  assign n6109 = Ng679 & n6564;
  assign n6110 = Ng686 & n6109;
  assign n6111_1 = (~n4555_1 | ~n4992) & (n4545 | ~n4984);
  assign n6112 = n4984 & (~n8531 | (n4549 & ~n4992));
  assign n6113 = n4555_1 & (~n8530 | (n4545 & ~n4986));
  assign n6114 = n4992 & n4986;
  assign n6115 = ~n4984 & (n6113 | (n4543 & n6114));
  assign n6116_1 = ~n4555_1 & (n6112 | (~n5000 & ~n6123));
  assign n6117 = ~n4992 | n4543 | n4549;
  assign n6118 = n6117 & (~n4545 | (n4549 & ~n4992));
  assign n6119 = n4992 & (n4555_1 | ~n5000);
  assign n6120_1 = n4545 & (~n5000 | (~n4549 & n6114));
  assign n6121 = ~n6120_1 & (n4543 | n4984 | n5000);
  assign n6122 = (~n4986 & (n4555_1 | n4992)) | (~n4555_1 & n4992);
  assign n6123 = n4545 | n4549;
  assign n6124_1 = (~n4543 | n6119) & (n6122 | n6123);
  assign n6125 = n4555_1 | n4986 | n6118;
  assign n6126 = (~n4984 & ~n7109) | (n6124_1 & (n4984 | ~n7109));
  assign n6127 = n6125 & (~n4555_1 | n6121) & n6126;
  assign n6128_1 = n1875_1 | ~Ng185 | ~Ng542;
  assign n6129 = (~\[1603]  | ~Ng599) & (~\[1605]  | ~Ng596);
  assign n6130 = n6128_1 & n6129 & (~Ng1315 | ~Ng602);
  assign n6131 = Ng3126 | Ng3191 | Ng3126 | Ng3110;
  assign n6132 = n5973_1 & n5978_1;
  assign n6133_1 = (n6542 | ~Ng3161) & (n6540_1 | ~Ng3155);
  assign n6134 = (n6543 | ~Ng3164) & (n6541 | ~Ng3158);
  assign n6135 = (n6545_1 | ~Ng3167) & (n6546 | ~Ng3170);
  assign n6136 = (n6548 | ~Ng3176) & (n6549 | ~Ng3179);
  assign n6137 = n6547 | ~Ng3173;
  assign n6138_1 = (n6536 | ~Ng3185) & (n6535_1 | ~Ng3182);
  assign n6139 = (n6132 | ~Ng3135) & (n6538 | ~Ng3088);
  assign n6140 = n6139 & n6138_1 & n6137 & n6136 & n6135 & ~n858_1 & n6133_1 & n6134;
  assign n6141 = (n6536 | ~Ng3095) & (n6538 | ~Ng3096);
  assign n6142 = (n6549 | ~Ng3093) & (n6535_1 | ~Ng3094);
  assign n6143_1 = (n6547 | ~Ng3091) & (n6548 | ~Ng3092);
  assign n6144 = (n6545_1 | ~Ng3086) & (n6546 | ~Ng3087);
  assign n6145 = (n6542 | ~Ng3084) & (n6543 | ~Ng3085);
  assign n6146 = (n6540_1 | ~Ng3210) & (n6541 | ~Ng3211);
  assign n6147_1 = n8532 & (~Ng3120 | (n5976 & n5978_1));
  assign n6148 = n6147_1 & n6146 & n6145 & n6144 & n6143_1 & ~n858_1 & n6141 & n6142;
  assign n6149 = Ng2175 & Ng2190 & Ng2185 & Ng2195 & Ng2200 & Ng2180 & Ng2165 & Ng2170;
  assign n6150 = n6149 & (~n8533 | (\[1594]  & ~Ng2255));
  assign n6151_1 = n4880_1 & (~n4908 | ~n6150);
  assign n6152 = ~n4880_1 & (n4908 | n6150);
  assign n6153 = ~Ng2257 | n6151_1 | n6152;
  assign n6154 = n6203_1 & Ng2151 & Ng2147;
  assign n6155_1 = n6154 & Ng2142;
  assign n6156 = Ng1481 & Ng1496 & Ng1491 & Ng1501 & Ng1506 & Ng1486 & Ng1471 & Ng1476;
  assign n6157 = n6156 & (~n8534 | (\[1594]  & ~Ng1561));
  assign n6158 = n4838_1 & (~n4870 | ~n6157);
  assign n6159_1 = ~n4838_1 & (n4870 | n6157);
  assign n6160 = ~Ng2257 | n6158 | n6159_1;
  assign n6161 = n6207_1 & Ng1457 & Ng1453;
  assign n6162 = n6161 & Ng1448;
  assign n6163_1 = Ng793 & Ng805 & Ng801 & Ng809 & Ng813 & Ng797 & Ng785 & Ng789;
  assign n6164 = n6163_1 & (~n8535 | (\[1594]  & ~Ng867));
  assign n6165 = n4796_1 & (~n4828 | ~n6164);
  assign n6166 = ~n4796_1 & (n4828 | n6164);
  assign n6167_1 = ~Ng2257 | n6165 | n6166;
  assign n6168 = n6211_1 & Ng771 & Ng767;
  assign n6169 = n6168 & Ng762;
  assign n6170 = Ng105 & Ng117 & Ng113 & Ng121 & Ng125 & Ng109 & Ng97 & Ng101;
  assign n6171_1 = n6170 & (~n8536 | (\[1594]  & ~Ng179));
  assign n6172 = n4754 & (~n4786 | ~n6171_1);
  assign n6173 = ~n4754 & (n4786 | n6171_1);
  assign n6174 = ~Ng2257 | n6172 | n6173;
  assign n6175_1 = n6215_1 & Ng83 & Ng79;
  assign n6176 = n6175_1 & Ng74;
  assign n6177 = ~n4581 | n4982 | ~Ng2584;
  assign n6178 = ~n5028_1 | Pg3229 | n5018_1;
  assign n6179_1 = n6178 & (~Pg3229 | n5036) & ~n8670;
  assign n6180 = ~n4926 | Pg3229 | n4906;
  assign n6181 = n6180 & (~Pg3229 | n4940) & ~n8675;
  assign n6182 = ~n4579 | n4978_1 | ~Ng1890;
  assign n6183_1 = ~n5016 | Pg3229 | n5006;
  assign n6184 = n6183_1 & (~Pg3229 | n5024) & ~n8681;
  assign n6185 = ~n4896 | Pg3229 | n4868;
  assign n6186 = n6185 & (~Pg3229 | n4920) & ~n8686;
  assign n6187_1 = ~n4577_1 | n4972 | ~Ng1196;
  assign n6188 = ~n5004 | Pg3229 | n4994;
  assign n6189 = n6188 & (~Pg3229 | n5012) & ~n8692;
  assign n6190 = ~n4858 | Pg3229 | n4826;
  assign n6191_1 = n6190 & (~Pg3229 | n4890) & ~n8697;
  assign n6192 = ~n4575 | n4964 | ~Ng510;
  assign n6193 = ~n4992 | Pg3229 | n4986;
  assign n6194 = n6193 & (~Pg3229 | n5000) & ~n8703;
  assign n6195_1 = ~n4816 | Pg3229 | n4784;
  assign n6196 = n6195_1 & (~Pg3229 | n4852) & ~n8708;
  assign n6197 = ~Ng3013 | n6573;
  assign n6198 = n6197 | ~Ng3010;
  assign n6199_1 = Ng2903 & n6574_1;
  assign n6200 = Ng2900 & n6199_1;
  assign n6201 = n6240 & Ng2734 & Ng2720;
  assign n6202 = n6201 & Ng2746;
  assign n6203_1 = ~n6242 & Ng2160 & Ng2156;
  assign n6204 = n6203_1 & Ng2151;
  assign n6205 = n6244_1 & Ng2040 & Ng2026;
  assign n6206 = n6205 & Ng2052;
  assign n6207_1 = ~n6242 & Ng1466 & Ng1462;
  assign n6208 = n6207_1 & Ng1457;
  assign n6209 = n6247 & Ng1346 & Ng1332;
  assign n6210 = n6209 & Ng1358;
  assign n6211_1 = ~n6242 & Ng780 & Ng776;
  assign n6212 = n6211_1 & Ng771;
  assign n6213 = n6250 & Ng660 & Ng646;
  assign n6214 = n6213 & Ng672;
  assign n6215_1 = ~n6242 & Ng92 & Ng88;
  assign n6216 = n6215_1 & Ng83;
  assign n6217 = n6395_1 | ~n5127 | ~n5137 | n6396 | n6397 | n6398;
  assign n6218 = n6404 | n6402 | n6403_1 | n6399_1 | n6400 | n6401;
  assign n6219_1 = ~n4980 | ~n4970 | ~n4976;
  assign n6143 = (n6217 | n6218) & (n6219_1 | ~n6487);
  assign n6221 = n6405 | ~n5127 | ~n5135_1 | n6406 | n6407 | n6408_1;
  assign n6222 = n6414 | n6412_1 | n6413 | n6409 | n6410 | n6411;
  assign n6223_1 = ~n4974 | ~n4962 | ~n4968_1;
  assign n4636 = (n6221 | n6222) & (n6223_1 | ~n6497);
  assign n6225 = n6415 | ~n5127 | ~n5131 | n6416 | n6417_1 | n6418;
  assign n6226 = n6424 | n6422_1 | n6423 | n6419 | n6420 | n6421;
  assign n6227_1 = ~n4966 | ~n4956 | ~n4960;
  assign n3129_1 = (n6225 | n6226) & (n6227_1 | ~n6507);
  assign n6229 = n6425 | ~n5126 | ~n5127 | n6426_1 | n6427 | n6428;
  assign n6230 = n6434 | n6432 | n6433 | n6429 | n6430 | n6431_1;
  assign n6231_1 = ~n4958_1 | ~n4950 | ~n4954;
  assign n1623_1 = (n6229 | n6230) & (n6231_1 | ~n6517);
  assign n6233 = ~Ng3028 & ~Ng3036 & Ng3032 & Ng3018;
  assign n6234 = n6256 | Pg3234;
  assign n6235_1 = n6256 & Ng3028 & Ng3018;
  assign n6236 = n6235_1 & Ng3036;
  assign n6237 = ~Ng2917 & ~Ng2924 & Ng2912 & Ng2920;
  assign n6238 = n6258 & Ng2912 & Ng2917;
  assign n6239_1 = n6238 & Ng2924;
  assign n6240 = n6260 & Ng2727 & Ng2707;
  assign n6241 = n6240 & Ng2720;
  assign n6242 = ~Ng853 | ~n5127;
  assign n6243 = n6242 | ~Ng2160;
  assign n6244_1 = n6262 & Ng2033 & Ng2013;
  assign n6245 = n6244_1 & Ng2026;
  assign n6246 = n6242 | ~Ng1466;
  assign n6247 = n6264 & Ng1339 & Ng1319;
  assign n6248 = n6247 & Ng1332;
  assign n6249_1 = n6242 | ~Ng780;
  assign n6250 = n6266 & Ng653 & Ng633;
  assign n6251 = n6250 & Ng646;
  assign n6252 = n6242 | ~Ng92;
  assign n6253 = ~n6572 | ~Ng3006;
  assign n6254_1 = Ng2883 & Ng13457 & Ng2888;
  assign n6255 = n6254_1 & Ng2896;
  assign n6256 = n6551 & Ng13475;
  assign n6257 = n6256 & Ng3018;
  assign n6258 = Ng2888 & Ng2908 & Ng2903 & Ng2892 & ~Ng2883 & Ng13457 & ~Ng2900 & ~Ng2896;
  assign n6259_1 = n6258 & Ng2912;
  assign n6260 = Ng1315 & ~Ng2733 & Ng2714;
  assign n6261 = n6260 & Ng2707;
  assign n6262 = Ng1315 & ~Ng2039 & Ng2020;
  assign n6263_1 = n6262 & Ng2013;
  assign n6264 = Ng1315 & ~Ng1345 & Ng1326;
  assign n6265 = n6264 & Ng1319;
  assign n6266 = Ng1315 & ~Ng659 & Ng640;
  assign n6267_1 = n6266 & Ng633;
  assign n6268 = Ng2883 & Ng13457;
  assign n6269 = ~Ng1315 | Ng2733;
  assign n6270 = ~Ng1315 | n6271;
  assign n6271 = Ng1315 & n6555_1;
  assign n6272_1 = ~Ng1315 | Ng2039;
  assign n6273 = ~Ng1315 | Ng1345;
  assign n6274 = ~Ng1315 | Ng659;
  assign n6275 = ~Ng1315 | n6276_1;
  assign n6276_1 = n8750 & Ng1315;
  assign n6277 = ~n5848_1 & n5851 & (n4643 | ~n5859);
  assign n6278 = ~n5868_1 & n5871 & (n4639 | ~n5879);
  assign n6279 = ~n5888_1 & n5891 & (n4633 | ~n5899);
  assign n6280 = ~n5908_1 & n5911 & (n4625 | ~n5919);
  assign n6281_1 = ~Ng185 | ~Ng3139;
  assign n6282 = n6281_1 & ~n6523 & (Ng3139 | ~n8756);
  assign n6283 = ~Pg3234 & (n6234 | ~n6394);
  assign n7111 = ~n6283;
  assign n6285_1 = n4744 ^ ~Ng2195;
  assign n6286 = n4874 ^ ~Ng2170;
  assign n6287 = n4680_1 ^ ~Ng2180;
  assign n6288 = n4668_1 ^ ~Ng2175;
  assign n6289 = n4772 ^ ~Ng2200;
  assign n6290_1 = n4718 ^ ~Ng2190;
  assign n6291 = n4698 ^ ~Ng2185;
  assign n6292 = n4842_1 ^ ~Ng2165;
  assign n6293 = n4924_1 ^ ~Ng2175;
  assign n6294_1 = n4902 ^ ~Ng2165;
  assign n6295 = n4720_1 ^ ~Ng2195;
  assign n6296 = n4938_1 ^ ~Ng2185;
  assign n6297 = n4810_1 ^ ~Ng2180;
  assign n6298 = n4904 ^ ~n5044;
  assign n6299_1 = n4876_1 ^ ~Ng2200;
  assign n6300 = n4774_1 ^ ~Ng2170;
  assign n6301 = n4938_1 ^ ~n5926;
  assign n6302 = ~n4902 ^ ~n5926;
  assign n6303_1 = ~n4774_1 ^ ~n5926;
  assign n6304 = ~n4924_1 ^ ~n5926;
  assign n6305 = ~n4810_1 ^ ~n5926;
  assign n6306 = n6304 | n6308_1;
  assign n6307 = n5864 | n6302;
  assign n6308_1 = n6303_1 | n6307;
  assign n6309 = n4658 ^ ~Ng1481;
  assign n6310 = n4666 ^ ~Ng1486;
  assign n6311 = n4800 ^ ~Ng1471;
  assign n6312_1 = n4678 ^ ~Ng1491;
  assign n6313 = n4832 ^ ~Ng1476;
  assign n6314 = n4694 ^ ~Ng1496;
  assign n6315 = n4736 ^ ~Ng1506;
  assign n6316 = n4714 ^ ~Ng1501;
  assign n6317_1 = n4894 ^ ~Ng1481;
  assign n6318 = n4864 ^ ~Ng1471;
  assign n6319 = n4696_1 ^ ~Ng1501;
  assign n6320 = n4918 ^ ~Ng1491;
  assign n6321_1 = n4768 ^ ~Ng1486;
  assign n6322 = n4866_1 ^ ~n5040;
  assign n6323 = n4834_1 ^ ~Ng1506;
  assign n6324 = n4738 ^ ~Ng1476;
  assign n6325 = n4918 ^ ~n5933_1;
  assign n6326_1 = ~n4864 ^ ~n5933_1;
  assign n6327 = ~n4738 ^ ~n5933_1;
  assign n6328 = ~n4894 ^ ~n5933_1;
  assign n6329 = ~n4768 ^ ~n5933_1;
  assign n6330 = n6328 | n6332;
  assign n6331_1 = n5884 | n6326_1;
  assign n6332 = n6327 | n6331_1;
  assign n6333 = n4651 ^ ~Ng793;
  assign n6334 = n4790 ^ ~Ng789;
  assign n6335 = n4706 ^ ~Ng813;
  assign n6336_1 = n4656_1 ^ ~Ng797;
  assign n6337 = n4690 ^ ~Ng809;
  assign n6338 = n4674 ^ ~Ng805;
  assign n6339 = n4664_1 ^ ~Ng801;
  assign n6340 = n4758 ^ ~Ng785;
  assign n6341_1 = n4856_1 ^ ~Ng793;
  assign n6342 = n4822 ^ ~Ng785;
  assign n6343 = n4676_1 ^ ~Ng809;
  assign n6344 = n4888_1 ^ ~Ng801;
  assign n6345_1 = n4732_1 ^ ~Ng797;
  assign n6346 = n4824_1 ^ ~n5032;
  assign n6347 = n4792_1 ^ ~Ng813;
  assign n6348 = n4708_1 ^ ~Ng789;
  assign n6349_1 = n4888_1 ^ ~n5940;
  assign n6350 = ~n4822 ^ ~n5940;
  assign n6351 = ~n4708_1 ^ ~n5940;
  assign n6352 = ~n4856_1 ^ ~n5940;
  assign n6353_1 = ~n4732_1 ^ ~n5940;
  assign n6354 = n6352 | n6356;
  assign n6355 = n5904 | n6350;
  assign n6356 = n6351 | n6355;
  assign n6357 = n4647 ^ ~Ng105;
  assign n6358_1 = n4748 ^ ~Ng101;
  assign n6359 = n4682 ^ ~Ng125;
  assign n6360 = n4649 ^ ~Ng109;
  assign n6361 = n4670 ^ ~Ng121;
  assign n6362 = n4660_1 ^ ~Ng117;
  assign n6363_1 = n4654 ^ ~Ng113;
  assign n6364 = n4722 ^ ~Ng97;
  assign n6365 = n4814_1 ^ ~Ng105;
  assign n6366 = n4780 ^ ~Ng97;
  assign n6367 = n4662 ^ ~Ng121;
  assign n6368_1 = n4850 ^ ~Ng113;
  assign n6369 = n4702 ^ ~Ng109;
  assign n6370 = n4782 ^ ~n5020;
  assign n6371 = n4750 ^ ~Ng125;
  assign n6372 = n4684_1 ^ ~Ng101;
  assign n6373_1 = n4850 ^ ~n5947;
  assign n6374 = ~n4780 ^ ~n5947;
  assign n6375 = ~n4684_1 ^ ~n5947;
  assign n6376 = ~n4814_1 ^ ~n5947;
  assign n6377 = ~n4702 ^ ~n5947;
  assign n6378_1 = n6376 | n6380;
  assign n6379 = n5924 | n6374;
  assign n6380 = n6375 | n6379;
  assign n6381 = ~n4846_1 ^ ~n5855;
  assign n6382 = (~Ng2190 | n5863_1) & (~n5865 | n6381);
  assign n6383_1 = ~n4804 ^ ~n5875;
  assign n6384 = (~Ng1496 | n5883_1) & (~n5885 | n6383_1);
  assign n6385 = ~n4762 ^ ~n5895;
  assign n6386 = (~Ng805 | n5903_1) & (~n5905 | n6385);
  assign n6387_1 = ~n4726 ^ ~n5915;
  assign n6388 = (~Ng117 | n5923_1) & (~n5925 | n6387_1);
  assign n6389 = Pg3229 ^ ~n4878;
  assign n6390 = Pg3229 ^ ~n4836;
  assign n6391_1 = Pg3229 ^ ~n4794;
  assign n6392 = Pg3229 ^ ~n4752_1;
  assign n6393 = Ng13475 & Ng2993;
  assign n6394 = ~n6393 ^ ~Ng2998;
  assign n6395_1 = n4904 ^ ~Ng2120;
  assign n6396 = n4876_1 ^ ~Ng2129;
  assign n6397 = n4746 ^ ~Ng2124;
  assign n6398 = n4720_1 ^ ~Ng2133;
  assign n6399_1 = n4924_1 ^ ~Ng2151;
  assign n6400 = n4938_1 ^ ~Ng2142;
  assign n6401 = n4846_1 ^ ~Ng2138;
  assign n6402 = n4902 ^ ~Ng2160;
  assign n6403_1 = n4810_1 ^ ~Ng2147;
  assign n6404 = n4774_1 ^ ~Ng2156;
  assign n6405 = n4866_1 ^ ~Ng1426;
  assign n6406 = n4834_1 ^ ~Ng1435;
  assign n6407 = n4716_1 ^ ~Ng1430;
  assign n6408_1 = n4696_1 ^ ~Ng1439;
  assign n6409 = n4894 ^ ~Ng1457;
  assign n6410 = n4918 ^ ~Ng1448;
  assign n6411 = n4804 ^ ~Ng1444;
  assign n6412_1 = n4864 ^ ~Ng1466;
  assign n6413 = n4768 ^ ~Ng1453;
  assign n6414 = n4738 ^ ~Ng1462;
  assign n6415 = n4824_1 ^ ~Ng740;
  assign n6416 = n4792_1 ^ ~Ng749;
  assign n6417_1 = n4692_1 ^ ~Ng744;
  assign n6418 = n4676_1 ^ ~Ng753;
  assign n6419 = n4856_1 ^ ~Ng771;
  assign n6420 = n4888_1 ^ ~Ng762;
  assign n6421 = n4762 ^ ~Ng758;
  assign n6422_1 = n4822 ^ ~Ng780;
  assign n6423 = n4732_1 ^ ~Ng767;
  assign n6424 = n4708_1 ^ ~Ng776;
  assign n6425 = n4782 ^ ~Ng52;
  assign n6426_1 = n4750 ^ ~Ng61;
  assign n6427 = n4672_1 ^ ~Ng56;
  assign n6428 = n4662 ^ ~Ng65;
  assign n6429 = n4814_1 ^ ~Ng83;
  assign n6430 = n4850 ^ ~Ng74;
  assign n6431_1 = n4726 ^ ~Ng70;
  assign n6432 = n4780 ^ ~Ng92;
  assign n6433 = n4702 ^ ~Ng79;
  assign n6434 = n4684_1 ^ ~Ng88;
  assign n6435_1 = n4952 ^ ~Ng2760;
  assign n6436 = n4942 ^ ~Ng2740;
  assign n6437 = n4948_1 ^ ~Ng2753;
  assign n6438 = n4778_1 ^ ~Ng2766;
  assign n6439 = n4812 ^ ~Ng2707;
  assign n6440_1 = n4910_1 ^ ~Ng2734;
  assign n6441 = n4848 ^ ~Ng2727;
  assign n6442 = n4882 ^ ~Ng2720;
  assign n6443 = n4928_1 ^ ~Ng2746;
  assign n6444 = n4776 ^ ~Ng2714;
  assign n6445_1 = n4944 ^ ~Ng2066;
  assign n6446 = n4922 ^ ~Ng2046;
  assign n6447 = n4936 ^ ~Ng2059;
  assign n6448 = n4742_1 ^ ~Ng2072;
  assign n6449 = n4770 ^ ~Ng2013;
  assign n6450_1 = n4872 ^ ~Ng2040;
  assign n6451 = n4806 ^ ~Ng2033;
  assign n6452 = n4840 ^ ~Ng2026;
  assign n6453 = n4898 ^ ~Ng2052;
  assign n6454 = n4740 ^ ~Ng2020;
  assign n6455_1 = n4932 ^ ~Ng1372;
  assign n6456 = n4892_1 ^ ~Ng1352;
  assign n6457 = n4916 ^ ~Ng1365;
  assign n6458 = n4712_1 ^ ~Ng1378;
  assign n6459 = n4734 ^ ~Ng1319;
  assign n6460_1 = n4830 ^ ~Ng1346;
  assign n6461 = n4764 ^ ~Ng1339;
  assign n6462 = n4798 ^ ~Ng1332;
  assign n6463 = n4860 ^ ~Ng1358;
  assign n6464 = n4710 ^ ~Ng1326;
  assign n6465_1 = n4912 ^ ~Ng686;
  assign n6466 = n4854 ^ ~Ng666;
  assign n6467 = n4886 ^ ~Ng679;
  assign n6468 = n4688_1 ^ ~Ng692;
  assign n6469 = n4704_1 ^ ~Ng633;
  assign n6470_1 = n4788 ^ ~Ng660;
  assign n6471 = n4728_1 ^ ~Ng653;
  assign n6472 = n4756_1 ^ ~Ng646;
  assign n6473 = n4818 ^ ~Ng672;
  assign n6474 = n4686 ^ ~Ng640;
  assign n6417 = ~n6603;
  assign n6476 = ~n5072_1 | n5591;
  assign n4910 = ~n6602_1;
  assign n6478 = ~n5070 | n5574;
  assign n6479 = ~n4808 ^ ~n5046;
  assign n6480_1 = ~n4844 ^ ~n5044;
  assign n6481 = n6290_1 | n6288 | n6289 | n6285_1 | n6286 | n6287;
  assign n6482 = n6295 | n6293 | n6294_1;
  assign n6483 = n5848_1 | n5854;
  assign n6484 = ~n5849 & n5850;
  assign n6485_1 = Ng2257 & n4946;
  assign n6486 = n4938_1 & n4720_1 & n4902 & n4846_1 & n4876_1;
  assign n6487 = n4904 & n4810_1 & n6486 & n4746 & n4924_1 & n4774_1;
  assign n6488 = n6304 | n6305;
  assign n6489 = ~n4766 ^ ~n5042;
  assign n6490_1 = ~n4802 ^ ~n5040;
  assign n6491 = n6314 | n6312_1 | n6313 | n6309 | n6310 | n6311;
  assign n6492 = n6319 | n6317_1 | n6318;
  assign n6493 = n5868_1 | n5874;
  assign n6494 = ~n5869 & n5870;
  assign n6495_1 = Ng2257 & n4934;
  assign n6496 = n4918 & n4696_1 & n4864 & n4804 & n4834_1;
  assign n6497 = n4866_1 & n4768 & n6496 & n4716_1 & n4894 & n4738;
  assign n6498 = n6328 | n6329;
  assign n6499 = ~n4730 ^ ~n5038_1;
  assign n6500_1 = ~n4760_1 ^ ~n5032;
  assign n6501 = n6338 | n6336_1 | n6337 | n6333 | n6334 | n6335;
  assign n6502 = n6343 | n6341_1 | n6342;
  assign n6503 = n5888_1 | n5894;
  assign n6504 = ~n5889 & n5890;
  assign n6505_1 = Ng2257 & n4914;
  assign n6506 = n4888_1 & n4676_1 & n4822 & n4762 & n4792_1;
  assign n6507 = n4824_1 & n4732_1 & n6506 & n4692_1 & n4856_1 & n4708_1;
  assign n6508 = n6352 | n6353_1;
  assign n6509 = ~n4700_1 ^ ~n5030;
  assign n6510_1 = ~n4724_1 ^ ~n5020;
  assign n6511 = n6362 | n6360 | n6361 | n6357 | n6358_1 | n6359;
  assign n6512 = n6367 | n6365 | n6366;
  assign n6513 = n5908_1 | n5914;
  assign n6514 = ~n5909 & n5910;
  assign n6515_1 = Ng2257 & n4884_1;
  assign n6516 = n4850 & n4662 & n4780 & n4726 & n4750;
  assign n6517 = n4782 & n4702 & n6516 & n4672_1 & n4814_1 & n4684_1;
  assign n6518 = n6376 | n6377;
  assign n3403_1 = ~n6601;
  assign n6520_1 = ~n5068 | n5549;
  assign n6521 = ~Ng853 | ~Ng2257;
  assign n6522 = Ng3139 | Ng3120;
  assign n6523 = Ng3126 | Ng3191 | Ng3126 | ~Ng3110;
  assign n6524 = Ng3139 | ~Ng3120;
  assign n1897_1 = ~n6600;
  assign n6526 = ~n5066 | n5523;
  assign n6527 = ~n5060 | n5672 | n5987;
  assign n6528 = ~n5056 | n5669 | n5995;
  assign n6529 = ~n5052 | n5666 | n6003_1;
  assign n6530_1 = ~n5050 | n5663 | n6011;
  assign n6531 = n6522 | n6131 | Ng3135 | Ng3147;
  assign n6532 = Ng3147 | n6523;
  assign n6533 = ~Ng3139 | Ng3120;
  assign n6534 = ~Ng3135 | n6532;
  assign n6535_1 = n6533 | n6534;
  assign n6536 = n5974 | n6532;
  assign n6537 = ~Ng3139 | ~Ng3120;
  assign n6538 = n6534 | n6537;
  assign n6539 = Ng3135 | n6532;
  assign n6540_1 = n6522 | n6539;
  assign n6541 = n6533 | n6539;
  assign n6542 = n6524 | n6539;
  assign n6543 = n6537 | n6539;
  assign n6544 = ~Ng3147 | n6523 | Ng3135;
  assign n6545_1 = n6522 | n6544;
  assign n6546 = n6533 | n6544;
  assign n6547 = n6524 | n6544;
  assign n6548 = n6537 | n6544;
  assign n6549 = n6522 | n6534;
  assign n6550_1 = n6201 & Ng2740 & Ng2746;
  assign n6551 = ~Ng3010 & ~Ng3006 & ~Ng2993 & Ng3002 & Ng3013 & Ng2998 & Ng3024;
  assign n6552 = ~n5018_1 | ~n5036;
  assign n6553 = n4571 & ~n5018_1 & ~n6045;
  assign n6554 = n6050 | n6553 | n6049;
  assign n6555_1 = Ng3028 & n6551 & ~Ng3032 & Ng3018 & ~Ng3036;
  assign n6556 = n6205 & Ng2046 & Ng2052;
  assign n6557 = ~n5006 | ~n5024;
  assign n6558 = n4565 & ~n5006 & ~n6067;
  assign n6559 = n6072 | n6558 | n6071_1;
  assign n6560_1 = n6209 & Ng1352 & Ng1358;
  assign n6561 = ~n4994 | ~n5012;
  assign n6562 = n4557 & ~n4994 & ~n6089_1;
  assign n6563 = n6094 | n6562 | n6093_1;
  assign n6564 = n6213 & Ng666 & Ng672;
  assign n6565_1 = ~n4986 | ~n5000;
  assign n6566 = n4549 & ~n4986 & ~n6111_1;
  assign n6567 = n6116_1 | n6566 | n6115;
  assign n6568 = n8661 & (n4880_1 | ~n4908 | ~n6150);
  assign n6569 = n8662 & (n4838_1 | ~n4870 | ~n6157);
  assign n6570_1 = n8663 & (n4796_1 | ~n4828 | ~n6164);
  assign n6571 = n8664 & (n4754 | ~n4786 | ~n6171_1);
  assign n6572 = Ng2998 & n6393;
  assign n6573 = ~Ng3006 | ~Ng3002 | ~n6572;
  assign n6574_1 = n6254_1 & Ng2892 & Ng2896;
  assign n6575 = Ng2599 & ~Ng2733 & Ng2612;
  assign n6576 = n5127 | Ng2912 | Ng2920 | ~Ng2924 | Ng2917 | ~Ng2883 | Ng2888;
  assign n6577 = Ng1905 & ~Ng2039 & Ng1918;
  assign n6578 = Ng1211 & ~Ng1345 & Ng1224;
  assign n6579_1 = Ng525 & ~Ng659 & Ng538;
  assign n6580 = ~n4902 ^ ~n5864;
  assign n6581 = ~n4864 ^ ~n5884;
  assign n6582 = ~n4822 ^ ~n5904;
  assign n6583 = ~n4780 ^ ~n5924;
  assign n6584_1 = ~Ng3024 ^ ~n6198;
  assign n6585 = ~n4880_1 ^ ~n6150;
  assign n6586 = ~n4838_1 ^ ~n6157;
  assign n6587_1 = ~n4796_1 ^ ~n6164;
  assign n6588 = ~n4754 ^ ~n6171_1;
  assign n6589 = ~n4532 ^ ~n4541_1;
  assign n7213 = ~Ng3083 ^ ~n6589;
  assign n6591 = ~n4535 ^ ~n4538;
  assign n7255 = ~Ng2990 ^ ~n6591;
  assign n7209 = n6589 ^ ~n8762;
  assign n7260 = n6591 ^ ~n8762;
  assign n6595 = ~n5607 ^ ~n5612;
  assign n344 = ~Ng2934 ^ ~n6595;
  assign n6597_1 = ~n5597 ^ ~n5602;
  assign n349_1 = ~Ng2962 ^ ~n6597_1;
  assign n6599 = (~n4952 & ~n8454) | (~n4982 & (n4952 | ~n8454));
  assign n6600 = n8550 & (~Ng8284 | ~Ng544);
  assign n6601 = (n8551 & (~Ng8293 | ~Ng1230)) | (Ng8293 & ~Ng1230);
  assign n6602_1 = (n8552 & (~Ng8302 | ~Ng1924)) | (Ng8302 & ~Ng1924);
  assign n6603 = (n8553 & (~Ng8311 | ~Ng2618)) | (Ng8311 & ~Ng2618);
  assign n6604 = (~n5064 & (n4778_1 | n8455)) | (~n4778_1 & n8455);
  assign n6605 = (~n5064 & (n4812 | n8455)) | (~n4812 & n8455);
  assign n6606 = (~n5064 & (n4882 | n8455)) | (~n4882 & n8455);
  assign n6607_1 = (~n4848 & ~n8454) | (~n4982 & (n4848 | ~n8454));
  assign n6608 = (Ng1315 & n6603) | (~Ng3108 & (~Ng1315 | n6603));
  assign n784_1 = ~n6608;
  assign n6610 = (\[1603]  & n6603) | (~Ng3107 & (~\[1603]  | n6603));
  assign n779 = ~n6610;
  assign n6612_1 = (\[1605]  & n6603) | (~Ng3106 & (~\[1605]  | n6603));
  assign n774 = ~n6612_1;
  assign n6614 = (~n4944 & ~n8452) | (~n4978_1 & (n4944 | ~n8452));
  assign n6615 = (~n5062 & (n4742_1 | n8453)) | (~n4742_1 & n8453);
  assign n6616 = (~n5062 & (n4770 | n8453)) | (~n4770 & n8453);
  assign n6617_1 = (~n5062 & (n4840 | n8453)) | (~n4840 & n8453);
  assign n6618 = (~n4806 & ~n8452) | (~n4978_1 & (n4806 | ~n8452));
  assign n6619 = (Ng853 & n8565) | (~Ng2392 & (~Ng853 | n8565));
  assign n6003 = ~n6619;
  assign n6621 = (\[1594]  & n8565) | (~Ng2391 & (~\[1594]  | n8565));
  assign n5998 = ~n6621;
  assign n6623 = (\[1612]  & n8565) | (~Ng2390 & (~\[1612]  | n8565));
  assign n5993 = ~n6623;
  assign n6625 = n6486 & ~n4924_1 & ~n4904 & ~n4810_1 & ~n4746 & ~n4774_1;
  assign n6626 = (~n5926 & n6625) | (n6487 & (n5926 | n6625));
  assign n6627_1 = (~Ng853 & ~Ng2348) | (~n5503 & (Ng853 | ~Ng2348));
  assign n5760 = ~n6627_1;
  assign n6629 = (~\[1594]  & ~Ng2345) | (~n5503 & (\[1594]  | ~Ng2345));
  assign n5755 = ~n6629;
  assign n6631 = (~\[1612]  & ~Ng2342) | (~n5503 & (\[1612]  | ~Ng2342));
  assign n5750 = ~n6631;
  assign n6633 = (~Ng853 & ~Ng2321) | (~n5485_1 & (Ng853 | ~Ng2321));
  assign n5670 = ~n6633;
  assign n6635 = (~\[1594]  & ~Ng2318) | (~n5485_1 & (\[1594]  | ~Ng2318));
  assign n5665 = ~n6635;
  assign n6637_1 = (~\[1612]  & ~Ng2315) | (~n5485_1 & (\[1612]  | ~Ng2315));
  assign n5660 = ~n6637_1;
  assign n6639 = (~Ng853 & ~Ng2312) | (~n5479 & (Ng853 | ~Ng2312));
  assign n5640 = ~n6639;
  assign n6641 = (~\[1594]  & ~Ng2309) | (~n5479 & (\[1594]  | ~Ng2309));
  assign n5635 = ~n6641;
  assign n6643 = (~\[1612]  & ~Ng2306) | (~n5479 & (\[1612]  | ~Ng2306));
  assign n5630 = ~n6643;
  assign n6645 = (~Ng853 & ~Ng2303) | (~n5473 & (Ng853 | ~Ng2303));
  assign n5745 = ~n6645;
  assign n6647_1 = (~\[1594]  & ~Ng2300) | (~n5473 & (\[1594]  | ~Ng2300));
  assign n5740 = ~n6647_1;
  assign n6649 = (~\[1612]  & ~Ng2297) | (~n5473 & (\[1612]  | ~Ng2297));
  assign n5735 = ~n6649;
  assign n6651 = (~Ng853 & ~Ng2276) | (~n5506 & (Ng853 | ~Ng2276));
  assign n5655 = ~n6651;
  assign n6653 = (~\[1594]  & ~Ng2273) | (~n5506 & (\[1594]  | ~Ng2273));
  assign n5650 = ~n6653;
  assign n6655 = (~\[1612]  & ~Ng2270) | (~n5506 & (\[1612]  | ~Ng2270));
  assign n5645 = ~n6655;
  assign n6657_1 = (Ng853 & n8570) | (~Ng1698 & (~Ng853 | n8570));
  assign n4496 = ~n6657_1;
  assign n6659 = (\[1594]  & n8570) | (~Ng1697 & (~\[1594]  | n8570));
  assign n4491 = ~n6659;
  assign n6661 = (\[1612]  & n8570) | (~Ng1696 & (~\[1612]  | n8570));
  assign n4486 = ~n6661;
  assign n6663 = n6496 & ~n4894 & ~n4866_1 & ~n4768 & ~n4716_1 & ~n4738;
  assign n6664 = (~n5933_1 & n6663) | (n6497 & (n5933_1 | n6663));
  assign n6665 = (~Ng853 & ~Ng1654) | (~n5497 & (Ng853 | ~Ng1654));
  assign n4266 = ~n6665;
  assign n6667_1 = (~\[1594]  & ~Ng1651) | (~n5497 & (\[1594]  | ~Ng1651));
  assign n4261_1 = ~n6667_1;
  assign n6669 = (~\[1612]  & ~Ng1648) | (~n5497 & (\[1612]  | ~Ng1648));
  assign n4256 = ~n6669;
  assign n6671 = (~Ng853 & ~Ng1627) | (~n5476 & (Ng853 | ~Ng1627));
  assign n4176 = ~n6671;
  assign n6673 = (~\[1594]  & ~Ng1624) | (~n5476 & (\[1594]  | ~Ng1624));
  assign n4171 = ~n6673;
  assign n6675 = (~\[1612]  & ~Ng1621) | (~n5476 & (\[1612]  | ~Ng1621));
  assign n4166 = ~n6675;
  assign n6677_1 = (~Ng853 & ~Ng1618) | (~n5470_1 & (Ng853 | ~Ng1618));
  assign n4146 = ~n6677_1;
  assign n6679 = (~\[1594]  & ~Ng1615) | (~n5470_1 & (\[1594]  | ~Ng1615));
  assign n4141 = ~n6679;
  assign n6681 = (~\[1612]  & ~Ng1612) | (~n5470_1 & (\[1612]  | ~Ng1612));
  assign n4136_1 = ~n6681;
  assign n6683 = (~Ng853 & ~Ng1609) | (~n5464 & (Ng853 | ~Ng1609));
  assign n4251 = ~n6683;
  assign n6685 = (~\[1594]  & ~Ng1606) | (~n5464 & (\[1594]  | ~Ng1606));
  assign n4246 = ~n6685;
  assign n6687_1 = (~\[1612]  & ~Ng1603) | (~n5464 & (\[1612]  | ~Ng1603));
  assign n4241_1 = ~n6687_1;
  assign n6689 = (~Ng853 & ~Ng1582) | (~n5500_1 & (Ng853 | ~Ng1582));
  assign n4161 = ~n6689;
  assign n6691 = (~\[1594]  & ~Ng1579) | (~n5500_1 & (\[1594]  | ~Ng1579));
  assign n4156 = ~n6691;
  assign n6693 = (~\[1612]  & ~Ng1576) | (~n5500_1 & (\[1612]  | ~Ng1576));
  assign n4151 = ~n6693;
  assign n6695 = (Ng853 & n8575) | (~Ng1004 & (~Ng853 | n8575));
  assign n2989_1 = ~n6695;
  assign n6697_1 = (\[1594]  & n8575) | (~Ng1003 & (~\[1594]  | n8575));
  assign n2984_1 = ~n6697_1;
  assign n6699 = (\[1612]  & n8575) | (~Ng1002 & (~\[1612]  | n8575));
  assign n2979_1 = ~n6699;
  assign n6701 = n6506 & ~n4856_1 & ~n4824_1 & ~n4732_1 & ~n4692_1 & ~n4708_1;
  assign n6702_1 = (~n5940 & n6701) | (n6507 & (n5940 | n6701));
  assign n6703 = (~Ng853 & ~Ng960) | (~n5491 & (Ng853 | ~Ng960));
  assign n2759_1 = ~n6703;
  assign n6705 = (~\[1594]  & ~Ng957) | (~n5491 & (\[1594]  | ~Ng957));
  assign n2754_1 = ~n6705;
  assign n6707_1 = (~\[1612]  & ~Ng954) | (~n5491 & (\[1612]  | ~Ng954));
  assign n2749_1 = ~n6707_1;
  assign n6709 = (~Ng853 & ~Ng933) | (~n5467 & (Ng853 | ~Ng933));
  assign n2669 = ~n6709;
  assign n6711 = (~\[1594]  & ~Ng930) | (~n5467 & (\[1594]  | ~Ng930));
  assign n2664 = ~n6711;
  assign n6713 = (~\[1612]  & ~Ng927) | (~n5467 & (\[1612]  | ~Ng927));
  assign n2659 = ~n6713;
  assign n6715 = (~Ng853 & ~Ng924) | (~n5461 & (Ng853 | ~Ng924));
  assign n2639 = ~n6715;
  assign n6717_1 = (~\[1594]  & ~Ng921) | (~n5461 & (\[1594]  | ~Ng921));
  assign n2634 = ~n6717_1;
  assign n6719 = (~\[1612]  & ~Ng918) | (~n5461 & (\[1612]  | ~Ng918));
  assign n2629 = ~n6719;
  assign n6721 = (~Ng853 & ~Ng915) | (~n5455_1 & (Ng853 | ~Ng915));
  assign n2744_1 = ~n6721;
  assign n6723 = (~\[1594]  & ~Ng912) | (~n5455_1 & (\[1594]  | ~Ng912));
  assign n2739_1 = ~n6723;
  assign n6725 = (~\[1612]  & ~Ng909) | (~n5455_1 & (\[1612]  | ~Ng909));
  assign n2734_1 = ~n6725;
  assign n6727_1 = (~Ng853 & ~Ng888) | (~n5494 & (Ng853 | ~Ng888));
  assign n2654 = ~n6727_1;
  assign n6729 = (~\[1594]  & ~Ng885) | (~n5494 & (\[1594]  | ~Ng885));
  assign n2649 = ~n6729;
  assign n6731 = (~\[1612]  & ~Ng882) | (~n5494 & (\[1612]  | ~Ng882));
  assign n2644 = ~n6731;
  assign n6733 = (Ng853 & n8580) | (~Ng317 & (~Ng853 | n8580));
  assign n1483_1 = ~n6733;
  assign n6735 = (\[1594]  & n8580) | (~Ng316 & (~\[1594]  | n8580));
  assign n1478_1 = ~n6735;
  assign n6737_1 = (\[1612]  & n8580) | (~Ng315 & (~\[1612]  | n8580));
  assign n1473_1 = ~n6737_1;
  assign n6739 = n6516 & ~n4814_1 & ~n4782 & ~n4702 & ~n4672_1 & ~n4684_1;
  assign n6740 = (~n5947 & n6739) | (n6517 & (n5947 | n6739));
  assign n6741 = (~Ng853 & ~Ng273) | (~n5482 & (Ng853 | ~Ng273));
  assign n1253_1 = ~n6741;
  assign n6743 = (~\[1594]  & ~Ng270) | (~n5482 & (\[1594]  | ~Ng270));
  assign n1248_1 = ~n6743;
  assign n6745 = (~\[1612]  & ~Ng267) | (~n5482 & (\[1612]  | ~Ng267));
  assign n1243_1 = ~n6745;
  assign n6747_1 = (~Ng853 & ~Ng246) | (~n5458 & (Ng853 | ~Ng246));
  assign n1163_1 = ~n6747_1;
  assign n6749 = (~\[1594]  & ~Ng243) | (~n5458 & (\[1594]  | ~Ng243));
  assign n1158_1 = ~n6749;
  assign n6751 = (~\[1612]  & ~Ng240) | (~n5458 & (\[1612]  | ~Ng240));
  assign n1153_1 = ~n6751;
  assign n6753 = (~Ng853 & ~Ng237) | (~n5452 & (Ng853 | ~Ng237));
  assign n1133_1 = ~n6753;
  assign n6755 = (~\[1594]  & ~Ng234) | (~n5452 & (\[1594]  | ~Ng234));
  assign n1128_1 = ~n6755;
  assign n6757_1 = (~\[1612]  & ~Ng231) | (~n5452 & (\[1612]  | ~Ng231));
  assign n1123_1 = ~n6757_1;
  assign n6759 = (~Ng853 & ~Ng228) | (~n5449 & (Ng853 | ~Ng228));
  assign n1238_1 = ~n6759;
  assign n6761 = (~\[1594]  & ~Ng225) | (~n5449 & (\[1594]  | ~Ng225));
  assign n1233_1 = ~n6761;
  assign n6763 = (~\[1612]  & ~Ng222) | (~n5449 & (\[1612]  | ~Ng222));
  assign n1228_1 = ~n6763;
  assign n6765 = (~Ng853 & ~Ng201) | (~n5488 & (Ng853 | ~Ng201));
  assign n1148_1 = ~n6765;
  assign n6767_1 = (~\[1594]  & ~Ng198) | (~n5488 & (\[1594]  | ~Ng198));
  assign n1143_1 = ~n6767_1;
  assign n6769 = (~\[1612]  & ~Ng195) | (~n5488 & (\[1612]  | ~Ng195));
  assign n1138_1 = ~n6769;
  assign n6771 = (~Ng853 & ~Ng2395) | (~n5446 & (Ng853 | ~Ng2395));
  assign n6018 = ~n6771;
  assign n6773 = (\[1594]  & ~n5446) | (~Ng2394 & (~\[1594]  | ~n5446));
  assign n6013 = ~n6773;
  assign n6775 = (~\[1612]  & ~Ng2393) | (~n5446 & (\[1612]  | ~Ng2393));
  assign n6008 = ~n6775;
  assign n6777_1 = (~Ng853 & ~Ng1701) | (~n5443 & (Ng853 | ~Ng1701));
  assign n4511 = ~n6777_1;
  assign n6779 = (\[1594]  & ~n5443) | (~Ng1700 & (~\[1594]  | ~n5443));
  assign n4506_1 = ~n6779;
  assign n6781 = (~\[1612]  & ~Ng1699) | (~n5443 & (\[1612]  | ~Ng1699));
  assign n4501 = ~n6781;
  assign n6783 = (~Ng853 & ~Ng1007) | (~n5440_1 & (Ng853 | ~Ng1007));
  assign n3004_1 = ~n6783;
  assign n6785 = (\[1594]  & ~n5440_1) | (~Ng1006 & (~\[1594]  | ~n5440_1));
  assign n2999 = ~n6785;
  assign n6787_1 = (~\[1612]  & ~Ng1005) | (~n5440_1 & (\[1612]  | ~Ng1005));
  assign n2994_1 = ~n6787_1;
  assign n6789 = (~Ng853 & ~Ng320) | (~n5437 & (Ng853 | ~Ng320));
  assign n1498 = ~n6789;
  assign n6791 = (\[1594]  & ~n5437) | (~Ng319 & (~\[1594]  | ~n5437));
  assign n1493 = ~n6791;
  assign n6793 = (~\[1612]  & ~Ng318) | (~n5437 & (\[1612]  | ~Ng318));
  assign n1488_1 = ~n6793;
  assign n6795 = (n5865 & n8585) | (n5929 & (~n5865 | n8585));
  assign n6796 = (Ng853 & ~n6795) | (~Ng2339 & (~Ng853 | ~n6795));
  assign n5730 = ~n6796;
  assign n6798 = (\[1594]  & ~n6795) | (~Ng2336 & (~\[1594]  | ~n6795));
  assign n5725 = ~n6798;
  assign n6800 = (\[1612]  & ~n6795) | (~Ng2333 & (~\[1612]  | ~n6795));
  assign n5720 = ~n6800;
  assign n6802_1 = (~Ng853 & ~Ng2330) | (n6382 & (Ng853 | ~Ng2330));
  assign n5700 = ~n6802_1;
  assign n6804 = (~\[1594]  & ~Ng2327) | (n6382 & (\[1594]  | ~Ng2327));
  assign n5695 = ~n6804;
  assign n6806 = (~\[1612]  & ~Ng2324) | (n6382 & (\[1612]  | ~Ng2324));
  assign n5690 = ~n6806;
  assign n6808 = (n5865 & n8586) | (n5930 & (~n5865 | n8586));
  assign n6809 = (Ng853 & ~n6808) | (~Ng2294 & (~Ng853 | ~n6808));
  assign n5715 = ~n6809;
  assign n6811 = (\[1594]  & ~n6808) | (~Ng2291 & (~\[1594]  | ~n6808));
  assign n5710 = ~n6811;
  assign n6813 = (\[1612]  & ~n6808) | (~Ng2288 & (~\[1612]  | ~n6808));
  assign n5705 = ~n6813;
  assign n6815 = (n5865 & n8588) | (n5931 & (~n5865 | n8588));
  assign n6816 = (Ng853 & ~n6815) | (~Ng2285 & (~Ng853 | ~n6815));
  assign n5685 = ~n6816;
  assign n6818 = (\[1594]  & ~n6815) | (~Ng2282 & (~\[1594]  | ~n6815));
  assign n5680 = ~n6818;
  assign n6820 = (\[1612]  & ~n6815) | (~Ng2279 & (~\[1612]  | ~n6815));
  assign n5675 = ~n6820;
  assign n6822_1 = (n5865 & n6580) | (n5932 & (~n5865 | n6580));
  assign n6823 = (Ng853 & ~n6822_1) | (~Ng2267 & (~Ng853 | ~n6822_1));
  assign n5625 = ~n6823;
  assign n6825 = (\[1594]  & ~n6822_1) | (~Ng2264 & (~\[1594]  | ~n6822_1));
  assign n5620 = ~n6825;
  assign n6827_1 = (\[1612]  & ~n6822_1) | (~Ng2261 & (~\[1612]  | ~n6822_1));
  assign n5615 = ~n6827_1;
  assign n6829 = (n5885 & n8589) | (n5936 & (~n5885 | n8589));
  assign n6830 = (Ng853 & ~n6829) | (~Ng1645 & (~Ng853 | ~n6829));
  assign n4236_1 = ~n6830;
  assign n6832_1 = (\[1594]  & ~n6829) | (~Ng1642 & (~\[1594]  | ~n6829));
  assign n4231 = ~n6832_1;
  assign n6834 = (\[1612]  & ~n6829) | (~Ng1639 & (~\[1612]  | ~n6829));
  assign n4226 = ~n6834;
  assign n6836 = (~Ng853 & ~Ng1636) | (n6384 & (Ng853 | ~Ng1636));
  assign n4206 = ~n6836;
  assign n6838 = (~\[1594]  & ~Ng1633) | (n6384 & (\[1594]  | ~Ng1633));
  assign n4201 = ~n6838;
  assign n6840 = (~\[1612]  & ~Ng1630) | (n6384 & (\[1612]  | ~Ng1630));
  assign n4196 = ~n6840;
  assign n6842_1 = (n5885 & n8590) | (n5937 & (~n5885 | n8590));
  assign n6843 = (Ng853 & ~n6842_1) | (~Ng1600 & (~Ng853 | ~n6842_1));
  assign n4221 = ~n6843;
  assign n6845 = (\[1594]  & ~n6842_1) | (~Ng1597 & (~\[1594]  | ~n6842_1));
  assign n4216 = ~n6845;
  assign n6847_1 = (\[1612]  & ~n6842_1) | (~Ng1594 & (~\[1612]  | ~n6842_1));
  assign n4211 = ~n6847_1;
  assign n6849 = (n5885 & n8592) | (n5938_1 & (~n5885 | n8592));
  assign n6850 = (Ng853 & ~n6849) | (~Ng1591 & (~Ng853 | ~n6849));
  assign n4191_1 = ~n6850;
  assign n6852_1 = (\[1594]  & ~n6849) | (~Ng1588 & (~\[1594]  | ~n6849));
  assign n4186 = ~n6852_1;
  assign n6854 = (\[1612]  & ~n6849) | (~Ng1585 & (~\[1612]  | ~n6849));
  assign n4181_1 = ~n6854;
  assign n6856 = (n5885 & n6581) | (n5939 & (~n5885 | n6581));
  assign n6857_1 = (Ng853 & ~n6856) | (~Ng1573 & (~Ng853 | ~n6856));
  assign n4131 = ~n6857_1;
  assign n6859 = (\[1594]  & ~n6856) | (~Ng1570 & (~\[1594]  | ~n6856));
  assign n4126 = ~n6859;
  assign n6861 = (\[1612]  & ~n6856) | (~Ng1567 & (~\[1612]  | ~n6856));
  assign n4121 = ~n6861;
  assign n6863 = (n5905 & n8593) | (n5943_1 & (~n5905 | n8593));
  assign n6864 = (Ng853 & ~n6863) | (~Ng951 & (~Ng853 | ~n6863));
  assign n2729_1 = ~n6864;
  assign n6866 = (\[1594]  & ~n6863) | (~Ng948 & (~\[1594]  | ~n6863));
  assign n2724_1 = ~n6866;
  assign n6868 = (\[1612]  & ~n6863) | (~Ng945 & (~\[1612]  | ~n6863));
  assign n2719 = ~n6868;
  assign n6870 = (~Ng853 & ~Ng942) | (n6386 & (Ng853 | ~Ng942));
  assign n2699_1 = ~n6870;
  assign n6872_1 = (~\[1594]  & ~Ng939) | (n6386 & (\[1594]  | ~Ng939));
  assign n2694_1 = ~n6872_1;
  assign n6874 = (~\[1612]  & ~Ng936) | (n6386 & (\[1612]  | ~Ng936));
  assign n2689 = ~n6874;
  assign n6876 = (n5905 & n8594) | (n5944 & (~n5905 | n8594));
  assign n6877_1 = (Ng853 & ~n6876) | (~Ng906 & (~Ng853 | ~n6876));
  assign n2714_1 = ~n6877_1;
  assign n6879 = (\[1594]  & ~n6876) | (~Ng903 & (~\[1594]  | ~n6876));
  assign n2709 = ~n6879;
  assign n6881 = (\[1612]  & ~n6876) | (~Ng900 & (~\[1612]  | ~n6876));
  assign n2704_1 = ~n6881;
  assign n6883 = (n5905 & n8596) | (n5945 & (~n5905 | n8596));
  assign n6884 = (Ng853 & ~n6883) | (~Ng897 & (~Ng853 | ~n6883));
  assign n2684 = ~n6884;
  assign n6886 = (\[1594]  & ~n6883) | (~Ng894 & (~\[1594]  | ~n6883));
  assign n2679 = ~n6886;
  assign n6888 = (\[1612]  & ~n6883) | (~Ng891 & (~\[1612]  | ~n6883));
  assign n2674 = ~n6888;
  assign n6890 = (n5905 & n6582) | (n5946 & (~n5905 | n6582));
  assign n6891 = (Ng853 & ~n6890) | (~Ng879 & (~Ng853 | ~n6890));
  assign n2624 = ~n6891;
  assign n6893 = (\[1594]  & ~n6890) | (~Ng876 & (~\[1594]  | ~n6890));
  assign n2619_1 = ~n6893;
  assign n6895 = (\[1612]  & ~n6890) | (~Ng873 & (~\[1612]  | ~n6890));
  assign n2614 = ~n6895;
  assign n6897_1 = (n5925 & n8597) | (n5950 & (~n5925 | n8597));
  assign n6898 = (Ng853 & ~n6897_1) | (~Ng264 & (~Ng853 | ~n6897_1));
  assign n1223_1 = ~n6898;
  assign n6900 = (\[1594]  & ~n6897_1) | (~Ng261 & (~\[1594]  | ~n6897_1));
  assign n1218_1 = ~n6900;
  assign n6902_1 = (\[1612]  & ~n6897_1) | (~Ng258 & (~\[1612]  | ~n6897_1));
  assign n1213_1 = ~n6902_1;
  assign n6904 = (~Ng853 & ~Ng255) | (n6388 & (Ng853 | ~Ng255));
  assign n1193_1 = ~n6904;
  assign n6906 = (~\[1594]  & ~Ng252) | (n6388 & (\[1594]  | ~Ng252));
  assign n1188_1 = ~n6906;
  assign n6908 = (~\[1612]  & ~Ng249) | (n6388 & (\[1612]  | ~Ng249));
  assign n1183_1 = ~n6908;
  assign n6910 = (n5925 & n8598) | (n5951 & (~n5925 | n8598));
  assign n6911 = (Ng853 & ~n6910) | (~Ng219 & (~Ng853 | ~n6910));
  assign n1208_1 = ~n6911;
  assign n6913 = (\[1594]  & ~n6910) | (~Ng216 & (~\[1594]  | ~n6910));
  assign n1203_1 = ~n6913;
  assign n6915 = (\[1612]  & ~n6910) | (~Ng213 & (~\[1612]  | ~n6910));
  assign n1198_1 = ~n6915;
  assign n6917_1 = (n5925 & n8600) | (n5952 & (~n5925 | n8600));
  assign n6918 = (Ng853 & ~n6917_1) | (~Ng210 & (~Ng853 | ~n6917_1));
  assign n1178 = ~n6918;
  assign n6920 = (\[1594]  & ~n6917_1) | (~Ng207 & (~\[1594]  | ~n6917_1));
  assign n1173_1 = ~n6920;
  assign n6922_1 = (\[1612]  & ~n6917_1) | (~Ng204 & (~\[1612]  | ~n6917_1));
  assign n1168_1 = ~n6922_1;
  assign n6924 = (n5925 & n6583) | (n5953_1 & (~n5925 | n6583));
  assign n6925 = (Ng853 & ~n6924) | (~Ng192 & (~Ng853 | ~n6924));
  assign n1118_1 = ~n6925;
  assign n6927 = (\[1594]  & ~n6924) | (~Ng189 & (~\[1594]  | ~n6924));
  assign n1113_1 = ~n6927;
  assign n6929 = (\[1612]  & ~n6924) | (~Ng186 & (~\[1612]  | ~n6924));
  assign n1108 = ~n6929;
  assign n5077 = (Ng1886 & Ng1887) | (n8605 & (~Ng1886 | Ng1887));
  assign n6932 = (Ng2580 & ~Ng2581) | (n8606 & (~Ng2580 | ~Ng2581));
  assign n6584 = ~n6932;
  assign n6934 = n8607 & (\[1594]  | ~Ng305 | ~Ng299);
  assign n1618_1 = ~n6934;
  assign n6936_1 = (~Ng986 & Ng985) | (n8608 & (Ng986 | Ng985));
  assign n3124_1 = ~n6936_1;
  assign n6938 = (~Ng1680 & Ng1679) | (n8609 & (Ng1680 | Ng1679));
  assign n4631 = ~n6938;
  assign n6940 = (~Ng2374 & Ng2373) | (n8610 & (Ng2374 | Ng2373));
  assign n6138 = ~n6940;
  assign n6942 = (Ng1315 & n6602_1) | (~Ng3105 & (~Ng1315 | n6602_1));
  assign n769_1 = ~n6942;
  assign n6944 = (\[1603]  & n6602_1) | (~Ng3104 & (~\[1603]  | n6602_1));
  assign n764_1 = ~n6944;
  assign n6946_1 = (\[1605]  & n6602_1) | (~Ng3103 & (~\[1605]  | n6602_1));
  assign n759_1 = ~n6946_1;
  assign n6948 = (~n4932 & ~n5528) | (~n4972 & (n4932 | ~n5528));
  assign n6949 = (~n5058_1 & (n4712_1 | n8451)) | (~n4712_1 & n8451);
  assign n6950 = (~n5058_1 & (n4734 | n8451)) | (~n4734 & n8451);
  assign n6951_1 = (~n5058_1 & (n4798 | n8451)) | (~n4798 & n8451);
  assign n6952 = (~n4764 & ~n5528) | (~n4972 & (n4764 | ~n5528));
  assign n6953 = (Ng853 & n8614) | (~Ng2389 & (~Ng853 | n8614));
  assign n5988 = ~n6953;
  assign n6955 = (\[1594]  & n8614) | (~Ng2388 & (~\[1594]  | n8614));
  assign n5983 = ~n6955;
  assign n6957 = (\[1612]  & n8614) | (~Ng2387 & (~\[1612]  | n8614));
  assign n5978 = ~n6957;
  assign n6959 = (Ng853 & n8615) | (~Ng1695 & (~Ng853 | n8615));
  assign n4481 = ~n6959;
  assign n6961_1 = (\[1594]  & n8615) | (~Ng1694 & (~\[1594]  | n8615));
  assign n4476 = ~n6961_1;
  assign n6963 = (\[1612]  & n8615) | (~Ng1693 & (~\[1612]  | n8615));
  assign n4471 = ~n6963;
  assign n6965 = (Ng853 & n8616) | (~Ng1001 & (~Ng853 | n8616));
  assign n2974_1 = ~n6965;
  assign n6967 = (\[1594]  & n8616) | (~Ng1000 & (~\[1594]  | n8616));
  assign n2969_1 = ~n6967;
  assign n6969 = (\[1612]  & n8616) | (~Ng999 & (~\[1612]  | n8616));
  assign n2964_1 = ~n6969;
  assign n6971_1 = (Ng853 & n8617) | (~Ng314 & (~Ng853 | n8617));
  assign n1468_1 = ~n6971_1;
  assign n6973 = (\[1594]  & n8617) | (~Ng313 & (~\[1594]  | n8617));
  assign n1463_1 = ~n6973;
  assign n6975 = (\[1612]  & n8617) | (~Ng312 & (~\[1612]  | n8617));
  assign n1458_1 = ~n6975;
  assign n6977 = (Ng3147 & n6282) | (~n6131 & (~Ng3147 | n6282));
  assign n6978 = (~n4912 & ~n5508) | (~n4964 & (n4912 | ~n5508));
  assign n6979 = (~n5054 & (n4688_1 | n8450)) | (~n4688_1 & n8450);
  assign n6980 = (~n5054 & (n4704_1 | n8450)) | (~n4704_1 & n8450);
  assign n6981_1 = (~n5054 & (n4756_1 | n8450)) | (~n4756_1 & n8450);
  assign n6982 = (~n4728_1 & ~n5508) | (~n4964 & (n4728_1 | ~n5508));
  assign n6983 = (Ng853 & n8621) | (~Ng2498 & (~Ng853 | n8621));
  assign n5913 = ~n6983;
  assign n6985 = (\[1594]  & n8621) | (~Ng2495 & (~\[1594]  | n8621));
  assign n5908 = ~n6985;
  assign n6987 = (\[1612]  & n8621) | (~Ng2492 & (~\[1612]  | n8621));
  assign n5903 = ~n6987;
  assign n6989 = (~Ng2396 & ~n8623) | (~n5991 & (~Ng2396 | n8623));
  assign n6033 = ~n6989;
  assign n6991_1 = (~n5991 & n8624) | (~Ng2398 & (~n5991 | ~n8624));
  assign n6028 = ~n6991_1;
  assign n6993 = (~Ng2397 & ~n8625) | (~n5991 & (~Ng2397 | n8625));
  assign n6023 = ~n6993;
  assign n6995 = (Ng853 & n8626) | (~Ng1804 & (~Ng853 | n8626));
  assign n4406 = ~n6995;
  assign n6997 = (\[1594]  & n8626) | (~Ng1801 & (~\[1594]  | n8626));
  assign n4401 = ~n6997;
  assign n6999 = (\[1612]  & n8626) | (~Ng1798 & (~\[1612]  | n8626));
  assign n4396 = ~n6999;
  assign n7001_1 = (~Ng1702 & ~n8628) | (~n5999 & (~Ng1702 | n8628));
  assign n4526 = ~n7001_1;
  assign n7003 = (~n5999 & n8629) | (~Ng1704 & (~n5999 | ~n8629));
  assign n4521 = ~n7003;
  assign n7005 = (~Ng1703 & ~n8630) | (~n5999 & (~Ng1703 | n8630));
  assign n4516 = ~n7005;
  assign n7007 = (Ng853 & n8631) | (~Ng1110 & (~Ng853 | n8631));
  assign n2899 = ~n7007;
  assign n7009 = (\[1594]  & n8631) | (~Ng1107 & (~\[1594]  | n8631));
  assign n2894 = ~n7009;
  assign n7011_1 = (\[1612]  & n8631) | (~Ng1104 & (~\[1612]  | n8631));
  assign n2889 = ~n7011_1;
  assign n7013 = (~Ng1008 & ~n8633) | (~n6007 & (~Ng1008 | n8633));
  assign n3019_1 = ~n7013;
  assign n7015 = (~n6007 & n8634) | (~Ng1010 & (~n6007 | ~n8634));
  assign n3014 = ~n7015;
  assign n7017 = (~Ng1009 & ~n8635) | (~n6007 & (~Ng1009 | n8635));
  assign n3009_1 = ~n7017;
  assign n7019 = (Ng853 & n8636) | (~Ng423 & (~Ng853 | n8636));
  assign n1393 = ~n7019;
  assign n7021_1 = (\[1594]  & n8636) | (~Ng420 & (~\[1594]  | n8636));
  assign n1388 = ~n7021_1;
  assign n7023 = (\[1612]  & n8636) | (~Ng417 & (~\[1612]  | n8636));
  assign n1383 = ~n7023;
  assign n7025 = (~Ng321 & ~n8638) | (~n6015 & (~Ng321 | n8638));
  assign n1513_1 = ~n7025;
  assign n7027 = (~n6015 & n8639) | (~Ng323 & (~n6015 | ~n8639));
  assign n1508 = ~n7027;
  assign n7029 = (~Ng322 & ~n8640) | (~n6015 & (~Ng322 | n8640));
  assign n1503 = ~n7029;
  assign n7031_1 = (Ng853 & n8642) | (~Ng2489 & (~Ng853 | n8642));
  assign n5898 = ~n7031_1;
  assign n7033 = (\[1594]  & n8642) | (~Ng2486 & (~\[1594]  | n8642));
  assign n5893 = ~n7033;
  assign n7035 = (\[1612]  & n8642) | (~Ng2483 & (~\[1612]  | n8642));
  assign n5888 = ~n7035;
  assign n7037 = (Ng853 & n8644) | (~Ng1795 & (~Ng853 | n8644));
  assign n4391 = ~n7037;
  assign n7039 = (\[1594]  & n8644) | (~Ng1792 & (~\[1594]  | n8644));
  assign n4386 = ~n7039;
  assign n7041_1 = (\[1612]  & n8644) | (~Ng1789 & (~\[1612]  | n8644));
  assign n4381 = ~n7041_1;
  assign n7043 = (Ng853 & n8646) | (~Ng1101 & (~Ng853 | n8646));
  assign n2884_1 = ~n7043;
  assign n7045 = (\[1594]  & n8646) | (~Ng1098 & (~\[1594]  | n8646));
  assign n2879_1 = ~n7045;
  assign n7047 = (\[1612]  & n8646) | (~Ng1095 & (~\[1612]  | n8646));
  assign n2874_1 = ~n7047;
  assign n7049 = (Ng853 & n8648) | (~Ng414 & (~Ng853 | n8648));
  assign n1378_1 = ~n7049;
  assign n7051_1 = (\[1594]  & n8648) | (~Ng411 & (~\[1594]  | n8648));
  assign n1373_1 = ~n7051_1;
  assign n7053 = (\[1612]  & n8648) | (~Ng408 & (~\[1612]  | n8648));
  assign n1368 = ~n7053;
  assign n7055 = (Ng1315 & n6601) | (~Ng3102 & (~Ng1315 | n6601));
  assign n754_1 = ~n7055;
  assign n7057 = (\[1603]  & n6601) | (~Ng3101 & (~\[1603]  | n6601));
  assign n749_1 = ~n7057;
  assign n7059 = (\[1605]  & n6601) | (~Ng3100 & (~\[1605]  | n6601));
  assign n744_1 = ~n7059;
  assign n7061_1 = n4571 & (~n6056 | (~n4567 & ~n6053_1));
  assign n7062 = (~n6061 & n6064) | (n5084 & (~n6061 | ~n6064));
  assign n7063 = (Ng1315 & n8650) | (~Ng2694 & (~Ng1315 | n8650));
  assign n6540 = ~n7063;
  assign n7065 = (\[1603]  & n8650) | (~Ng2691 & (~\[1603]  | n8650));
  assign n6535 = ~n7065;
  assign n7067 = (\[1605]  & n8650) | (~Ng2688 & (~\[1605]  | n8650));
  assign n6530 = ~n7067;
  assign n7069 = n5084 | n6064;
  assign n7070 = n6061 & n7069 & (~n5084 | n6554);
  assign n7071_1 = (Ng1315 & n8651) | (~Ng2685 & (~Ng1315 | n8651));
  assign n6555 = ~n7071_1;
  assign n7073 = (\[1603]  & n8651) | (~Ng2682 & (~\[1603]  | n8651));
  assign n6550 = ~n7073;
  assign n7075 = (\[1605]  & n8651) | (~Ng2679 & (~\[1605]  | n8651));
  assign n6545 = ~n7075;
  assign n7077 = n4565 & (~n6078 | (~n4559_1 & ~n6075_1));
  assign n7078 = (~n6083 & n6086) | (n5081 & (~n6083 | ~n6086));
  assign n7079 = (Ng1315 & n8653) | (~Ng2000 & (~Ng1315 | n8653));
  assign n5033 = ~n7079;
  assign n7081_1 = (\[1603]  & n8653) | (~Ng1997 & (~\[1603]  | n8653));
  assign n5028 = ~n7081_1;
  assign n7083 = (\[1605]  & n8653) | (~Ng1994 & (~\[1605]  | n8653));
  assign n5023 = ~n7083;
  assign n7085 = n5081 | n6086;
  assign n7086_1 = n6083 & n7085 & (~n5081 | n6559);
  assign n7087 = (Ng1315 & n8654) | (~Ng1991 & (~Ng1315 | n8654));
  assign n5048 = ~n7087;
  assign n7089 = (\[1603]  & n8654) | (~Ng1988 & (~\[1603]  | n8654));
  assign n5043 = ~n7089;
  assign n7091_1 = (\[1605]  & n8654) | (~Ng1985 & (~\[1605]  | n8654));
  assign n5038 = ~n7091_1;
  assign n7093 = n4557 & (~n6100 | (~n4551 & ~n6097));
  assign n7094 = (~n6105 & n6108) | (n5078 & (~n6105 | ~n6108));
  assign n7095 = (Ng1315 & n8656) | (~Ng1306 & (~Ng1315 | n8656));
  assign n3526_1 = ~n7095;
  assign n7097 = (\[1603]  & n8656) | (~Ng1303 & (~\[1603]  | n8656));
  assign n3521_1 = ~n7097;
  assign n7099 = (\[1605]  & n8656) | (~Ng1300 & (~\[1605]  | n8656));
  assign n3516_1 = ~n7099;
  assign n7101_1 = n5078 | n6108;
  assign n7102 = n6105 & n7101_1 & (~n5078 | n6563);
  assign n7103 = (Ng1315 & n8657) | (~Ng1297 & (~Ng1315 | n8657));
  assign n3541_1 = ~n7103;
  assign n7105 = (\[1603]  & n8657) | (~Ng1294 & (~\[1603]  | n8657));
  assign n3536_1 = ~n7105;
  assign n7107 = (\[1605]  & n8657) | (~Ng1291 & (~\[1605]  | n8657));
  assign n3531_1 = ~n7107;
  assign n7109 = n4549 & (~n6122 | (~n4545 & ~n6119));
  assign n7110 = (~n6127 & n6130) | (n5075 & (~n6127 | ~n6130));
  assign n7111_1 = (Ng1315 & n8659) | (~Ng620 & (~Ng1315 | n8659));
  assign n2020_1 = ~n7111_1;
  assign n7113 = (\[1603]  & n8659) | (~Ng617 & (~\[1603]  | n8659));
  assign n2015_1 = ~n7113;
  assign n7115 = (\[1605]  & n8659) | (~Ng614 & (~\[1605]  | n8659));
  assign n2010 = ~n7115;
  assign n7117 = n5075 | n6130;
  assign n7118 = n6127 & n7117 & (~n5075 | n6567);
  assign n7119 = (Ng1315 & n8660) | (~Ng611 & (~Ng1315 | n8660));
  assign n2035_1 = ~n7119;
  assign n7121_1 = (\[1603]  & n8660) | (~Ng608 & (~\[1603]  | n8660));
  assign n2030 = ~n7121_1;
  assign n7123 = (\[1605]  & n8660) | (~Ng605 & (~\[1605]  | n8660));
  assign n2025_1 = ~n7123;
  assign n7125 = (~n8665 & n8666) | (~Ng2658 & (n8665 | n8666));
  assign n6495 = ~n7125;
  assign n7127 = (n8666 & ~n8667) | (~Ng2660 & (n8666 | n8667));
  assign n6490 = ~n7127;
  assign n7129 = (n8666 & ~n8668) | (~Ng2659 & (n8666 | n8668));
  assign n6485 = ~n7129;
  assign n7131_1 = (n6552 & ~n8669) | (n5018_1 & (n6552 | n8669));
  assign n7132 = (~Ng2655 & n8665) | (~n7131_1 & (~Ng2655 | ~n8665));
  assign n6480 = ~n7132;
  assign n7134 = (~n7131_1 & ~n8667) | (~Ng2657 & (~n7131_1 | n8667));
  assign n6475 = ~n7134;
  assign n7136_1 = (~Ng2656 & n8668) | (~n7131_1 & (~Ng2656 | ~n8668));
  assign n6470 = ~n7136_1;
  assign n7138 = (~n5028_1 & n8669) | (n5018_1 & (n5028_1 | n8669));
  assign n7139 = (~Ng2652 & n8665) | (~n7138 & (~Ng2652 | ~n8665));
  assign n6465 = ~n7139;
  assign n7141_1 = (~n7138 & ~n8667) | (~Ng2654 & (~n7138 | n8667));
  assign n6460 = ~n7141_1;
  assign n7143 = (~Ng2653 & n8668) | (~n7138 & (~Ng2653 | ~n8668));
  assign n6455 = ~n7143;
  assign n7145 = (~Ng2649 & n8665) | (~n6179_1 & (~Ng2649 | ~n8665));
  assign n6450 = ~n7145;
  assign n7147 = (~n6179_1 & ~n8667) | (~Ng2651 & (~n6179_1 | n8667));
  assign n6445 = ~n7147;
  assign n7149 = (~Ng2650 & n8668) | (~n6179_1 & (~Ng2650 | ~n8668));
  assign n6440 = ~n7149;
  assign n7151_1 = (n8671 & n8672) | (~Ng11589 & (~n8671 | n8672));
  assign n5883 = ~n7151_1;
  assign n7153 = (n8672 & n8673) | (~Ng11588 & (n8672 | ~n8673));
  assign n5878 = ~n7153;
  assign n7155 = (n8672 & n8674) | (~Ng11587 & (n8672 | ~n8674));
  assign n5873 = ~n7155;
  assign n7157 = (n4906 | ~n6389) & ~n8764;
  assign n7158 = (~Ng11586 & ~n8671) | (~n7157 & (~Ng11586 | n8671));
  assign n5868 = ~n7158;
  assign n7160_1 = (~n7157 & n8673) | (~Ng11585 & (~n7157 | ~n8673));
  assign n5863 = ~n7160_1;
  assign n7162 = (~Ng11584 & ~n8674) | (~n7157 & (~Ng11584 | n8674));
  assign n5858 = ~n7162;
  assign n7164 = (~n4926 & n6389) | (n4906 & (n4926 | n6389));
  assign n7165 = (~Ng11583 & ~n8671) | (~n7164 & (~Ng11583 | n8671));
  assign n5853 = ~n7165;
  assign n7167_1 = (~n7164 & n8673) | (~Ng11582 & (~n7164 | ~n8673));
  assign n5848 = ~n7167_1;
  assign n7169 = (~Ng11581 & ~n8674) | (~n7164 & (~Ng11581 | n8674));
  assign n5843 = ~n7169;
  assign n7171 = (~Ng11580 & ~n8671) | (~n6181 & (~Ng11580 | n8671));
  assign n5838 = ~n7171;
  assign n7173 = (~n6181 & n8673) | (~Ng11579 & (~n6181 | ~n8673));
  assign n5833 = ~n7173;
  assign n7175 = (~Ng11578 & ~n8674) | (~n6181 & (~Ng11578 | n8674));
  assign n5828 = ~n7175;
  assign n7177 = (~n8676 & n8677) | (~Ng1964 & (n8676 | n8677));
  assign n4988 = ~n7177;
  assign n7179 = (n8677 & ~n8678) | (~Ng1966 & (n8677 | n8678));
  assign n4983 = ~n7179;
  assign n7181 = (n8677 & ~n8679) | (~Ng1965 & (n8677 | n8679));
  assign n4978 = ~n7181;
  assign n7183 = (n6557 & ~n8680) | (n5006 & (n6557 | n8680));
  assign n7184_1 = (~Ng1961 & n8676) | (~n7183 & (~Ng1961 | ~n8676));
  assign n4973 = ~n7184_1;
  assign n7186 = (~n7183 & ~n8678) | (~Ng1963 & (~n7183 | n8678));
  assign n4968 = ~n7186;
  assign n7188_1 = (~Ng1962 & n8679) | (~n7183 & (~Ng1962 | ~n8679));
  assign n4963 = ~n7188_1;
  assign n7190 = (~n5016 & n8680) | (n5006 & (n5016 | n8680));
  assign n7191 = (~Ng1958 & n8676) | (~n7190 & (~Ng1958 | ~n8676));
  assign n4958 = ~n7191;
  assign n7193 = (~n7190 & ~n8678) | (~Ng1960 & (~n7190 | n8678));
  assign n4953 = ~n7193;
  assign n7195 = (~Ng1959 & n8679) | (~n7190 & (~Ng1959 | ~n8679));
  assign n4948 = ~n7195;
  assign n7197 = (~Ng1955 & n8676) | (~n6184 & (~Ng1955 | ~n8676));
  assign n4943 = ~n7197;
  assign n7199 = (~n6184 & ~n8678) | (~Ng1957 & (~n6184 | n8678));
  assign n4938 = ~n7199;
  assign n7201 = (~Ng1956 & n8679) | (~n6184 & (~Ng1956 | ~n8679));
  assign n4933 = ~n7201;
  assign n7203 = (n8682 & n8683) | (~Ng11562 & (~n8682 | n8683));
  assign n4376 = ~n7203;
  assign n7205 = (n8683 & n8684) | (~Ng11561 & (n8683 | ~n8684));
  assign n4371 = ~n7205;
  assign n7207 = (n8683 & n8685) | (~Ng11560 & (n8683 | ~n8685));
  assign n4366 = ~n7207;
  assign n7209_1 = (n4868 | ~n6390) & ~n8765;
  assign n7210 = (~Ng11559 & ~n8682) | (~n7209_1 & (~Ng11559 | n8682));
  assign n4361 = ~n7210;
  assign n7212 = (~n7209_1 & n8684) | (~Ng11558 & (~n7209_1 | ~n8684));
  assign n4356 = ~n7212;
  assign n7214 = (~Ng11557 & ~n8685) | (~n7209_1 & (~Ng11557 | n8685));
  assign n4351 = ~n7214;
  assign n7216 = (~n4896 & n6390) | (n4868 & (n4896 | n6390));
  assign n7217 = (~Ng11556 & ~n8682) | (~n7216 & (~Ng11556 | n8682));
  assign n4346 = ~n7217;
  assign n7219 = (~n7216 & n8684) | (~Ng11555 & (~n7216 | ~n8684));
  assign n4341_1 = ~n7219;
  assign n7221 = (~Ng11554 & ~n8685) | (~n7216 & (~Ng11554 | n8685));
  assign n4336_1 = ~n7221;
  assign n7223 = (~Ng11553 & ~n8682) | (~n6186 & (~Ng11553 | n8682));
  assign n4331_1 = ~n7223;
  assign n7225 = (~n6186 & n8684) | (~Ng11552 & (~n6186 | ~n8684));
  assign n4326 = ~n7225;
  assign n7227 = (~Ng11551 & ~n8685) | (~n6186 & (~Ng11551 | n8685));
  assign n4321 = ~n7227;
  assign n7229 = (~n8687 & n8688) | (~Ng1270 & (n8687 | n8688));
  assign n3481_1 = ~n7229;
  assign n7231 = (n8688 & ~n8689) | (~Ng1272 & (n8688 | n8689));
  assign n3476_1 = ~n7231;
  assign n7233 = (n8688 & ~n8690) | (~Ng1271 & (n8688 | n8690));
  assign n3471_1 = ~n7233;
  assign n7235 = (n6561 & ~n8691) | (n4994 & (n6561 | n8691));
  assign n7236 = (~Ng1267 & n8687) | (~n7235 & (~Ng1267 | ~n8687));
  assign n3466_1 = ~n7236;
  assign n7238_1 = (~n7235 & ~n8689) | (~Ng1269 & (~n7235 | n8689));
  assign n3461_1 = ~n7238_1;
  assign n7240 = (~Ng1268 & n8690) | (~n7235 & (~Ng1268 | ~n8690));
  assign n3456_1 = ~n7240;
  assign n7242_1 = (~n5004 & n8691) | (n4994 & (n5004 | n8691));
  assign n7243 = (~Ng1264 & n8687) | (~n7242_1 & (~Ng1264 | ~n8687));
  assign n3451_1 = ~n7243;
  assign n7245 = (~n7242_1 & ~n8689) | (~Ng1266 & (~n7242_1 | n8689));
  assign n3446_1 = ~n7245;
  assign n7247 = (~Ng1265 & n8690) | (~n7242_1 & (~Ng1265 | ~n8690));
  assign n3441_1 = ~n7247;
  assign n7249 = (~Ng1261 & n8687) | (~n6189 & (~Ng1261 | ~n8687));
  assign n3436_1 = ~n7249;
  assign n7251 = (~n6189 & ~n8689) | (~Ng1263 & (~n6189 | n8689));
  assign n3431_1 = ~n7251;
  assign n7253 = (~Ng1262 & n8690) | (~n6189 & (~Ng1262 | ~n8690));
  assign n3426_1 = ~n7253;
  assign n7255_1 = (n8693 & n8694) | (~Ng11535 & (~n8693 | n8694));
  assign n2869_1 = ~n7255_1;
  assign n7257 = (n8694 & n8695) | (~Ng11534 & (n8694 | ~n8695));
  assign n2864_1 = ~n7257;
  assign n7259 = (n8694 & n8696) | (~Ng11533 & (n8694 | ~n8696));
  assign n2859_1 = ~n7259;
  assign n7261 = (n4826 | ~n6391_1) & ~n8766;
  assign n7262 = (~Ng11532 & ~n8693) | (~n7261 & (~Ng11532 | n8693));
  assign n2854_1 = ~n7262;
  assign n7264 = (~n7261 & n8695) | (~Ng11531 & (~n7261 | ~n8695));
  assign n2849_1 = ~n7264;
  assign n7266 = (~Ng11530 & ~n8696) | (~n7261 & (~Ng11530 | n8696));
  assign n2844_1 = ~n7266;
  assign n7268 = (~n4858 & n6391_1) | (n4826 & (n4858 | n6391_1));
  assign n7269 = (~Ng11529 & ~n8693) | (~n7268 & (~Ng11529 | n8693));
  assign n2839_1 = ~n7269;
  assign n7271 = (~n7268 & n8695) | (~Ng11528 & (~n7268 | ~n8695));
  assign n2834_1 = ~n7271;
  assign n7273 = (~Ng11527 & ~n8696) | (~n7268 & (~Ng11527 | n8696));
  assign n2829_1 = ~n7273;
  assign n7275 = (~Ng11526 & ~n8693) | (~n6191_1 & (~Ng11526 | n8693));
  assign n2824_1 = ~n7275;
  assign n7277 = (~n6191_1 & n8695) | (~Ng11525 & (~n6191_1 | ~n8695));
  assign n2819_1 = ~n7277;
  assign n7279 = (~Ng11524 & ~n8696) | (~n6191_1 & (~Ng11524 | n8696));
  assign n2814_1 = ~n7279;
  assign n7281 = (~n8698 & n8699) | (~Ng584 & (n8698 | n8699));
  assign n1975 = ~n7281;
  assign n7283 = (n8699 & ~n8700) | (~Ng586 & (n8699 | n8700));
  assign n1970_1 = ~n7283;
  assign n7285 = (n8699 & ~n8701) | (~Ng585 & (n8699 | n8701));
  assign n1965 = ~n7285;
  assign n7287 = (n6565_1 & ~n8702) | (n4986 & (n6565_1 | n8702));
  assign n7288 = (~Ng581 & n8698) | (~n7287 & (~Ng581 | ~n8698));
  assign n1960_1 = ~n7288;
  assign n7290 = (~n7287 & ~n8700) | (~Ng583 & (~n7287 | n8700));
  assign n1955 = ~n7290;
  assign n7292 = (~Ng582 & n8701) | (~n7287 & (~Ng582 | ~n8701));
  assign n1950 = ~n7292;
  assign n7294 = (~n4992 & n8702) | (n4986 & (n4992 | n8702));
  assign n7295 = (~Ng578 & n8698) | (~n7294 & (~Ng578 | ~n8698));
  assign n1945_1 = ~n7295;
  assign n7297 = (~n7294 & ~n8700) | (~Ng580 & (~n7294 | n8700));
  assign n1940_1 = ~n7297;
  assign n7299 = (~Ng579 & n8701) | (~n7294 & (~Ng579 | ~n8701));
  assign n1935_1 = ~n7299;
  assign n7301 = (~Ng575 & n8698) | (~n6194 & (~Ng575 | ~n8698));
  assign n1930_1 = ~n7301;
  assign n7303 = (~n6194 & ~n8700) | (~Ng577 & (~n6194 | n8700));
  assign n1925 = ~n7303;
  assign n7305 = (~Ng576 & n8701) | (~n6194 & (~Ng576 | ~n8701));
  assign n1920_1 = ~n7305;
  assign n7307 = (n8704 & n8705) | (~Ng11508 & (~n8704 | n8705));
  assign n1363_1 = ~n7307;
  assign n7309 = (n8705 & n8706) | (~Ng11507 & (n8705 | ~n8706));
  assign n1358_1 = ~n7309;
  assign n7311 = (n8705 & n8707) | (~Ng11506 & (n8705 | ~n8707));
  assign n1353 = ~n7311;
  assign n7313 = (n4784 | ~n6392) & ~n8767;
  assign n7314 = (~Ng11505 & ~n8704) | (~n7313 & (~Ng11505 | n8704));
  assign n1348 = ~n7314;
  assign n7316 = (~n7313 & n8706) | (~Ng11504 & (~n7313 | ~n8706));
  assign n1343_1 = ~n7316;
  assign n7318 = (~Ng11503 & ~n8707) | (~n7313 & (~Ng11503 | n8707));
  assign n1338_1 = ~n7318;
  assign n7320 = (~n4816 & n6392) | (n4784 & (n4816 | n6392));
  assign n7321 = (~Ng11502 & ~n8704) | (~n7320 & (~Ng11502 | n8704));
  assign n1333_1 = ~n7321;
  assign n7323 = (~n7320 & n8706) | (~Ng11501 & (~n7320 | ~n8706));
  assign n1328_1 = ~n7323;
  assign n7325 = (~Ng11500 & ~n8707) | (~n7320 & (~Ng11500 | n8707));
  assign n1323_1 = ~n7325;
  assign n7327 = (~Ng11499 & ~n8704) | (~n6196 & (~Ng11499 | n8704));
  assign n1318 = ~n7327;
  assign n7329 = (~n6196 & n8706) | (~Ng11498 & (~n6196 | ~n8706));
  assign n1313 = ~n7329;
  assign n7331 = (~Ng11497 & ~n8707) | (~n6196 & (~Ng11497 | n8707));
  assign n1308_1 = ~n7331;
  assign n7333 = (Ng853 & n8709) | (~Ng2519 & (~Ng853 | n8709));
  assign n5958 = ~n7333;
  assign n7335 = (\[1594]  & n8709) | (~Ng2516 & (~\[1594]  | n8709));
  assign n5953 = ~n7335;
  assign n7337 = (\[1612]  & n8709) | (~Ng2513 & (~\[1612]  | n8709));
  assign n5948 = ~n7337;
  assign n7339 = (Ng853 & n8710) | (~Ng2510 & (~Ng853 | n8710));
  assign n5943 = ~n7339;
  assign n7341 = (\[1594]  & n8710) | (~Ng2507 & (~\[1594]  | n8710));
  assign n5938 = ~n7341;
  assign n7343 = (\[1612]  & n8710) | (~Ng2504 & (~\[1612]  | n8710));
  assign n5933 = ~n7343;
  assign n7345 = (Ng853 & n8711) | (~Ng1825 & (~Ng853 | n8711));
  assign n4451_1 = ~n7345;
  assign n7347 = (\[1594]  & n8711) | (~Ng1822 & (~\[1594]  | n8711));
  assign n4446_1 = ~n7347;
  assign n7349 = (\[1612]  & n8711) | (~Ng1819 & (~\[1612]  | n8711));
  assign n4441 = ~n7349;
  assign n7351 = (Ng853 & n8712) | (~Ng1816 & (~Ng853 | n8712));
  assign n4436 = ~n7351;
  assign n7353 = (\[1594]  & n8712) | (~Ng1813 & (~\[1594]  | n8712));
  assign n4431 = ~n7353;
  assign n7355 = (\[1612]  & n8712) | (~Ng1810 & (~\[1612]  | n8712));
  assign n4426 = ~n7355;
  assign n7357 = (Ng853 & n8713) | (~Ng1131 & (~Ng853 | n8713));
  assign n2944_1 = ~n7357;
  assign n7359 = (\[1594]  & n8713) | (~Ng1128 & (~\[1594]  | n8713));
  assign n2939_1 = ~n7359;
  assign n7361 = (\[1612]  & n8713) | (~Ng1125 & (~\[1612]  | n8713));
  assign n2934_1 = ~n7361;
  assign n7363 = (Ng853 & n8714) | (~Ng1122 & (~Ng853 | n8714));
  assign n2929_1 = ~n7363;
  assign n7365 = (\[1594]  & n8714) | (~Ng1119 & (~\[1594]  | n8714));
  assign n2924_1 = ~n7365;
  assign n7367 = (\[1612]  & n8714) | (~Ng1116 & (~\[1612]  | n8714));
  assign n2919_1 = ~n7367;
  assign n7369 = (Ng853 & n8715) | (~Ng444 & (~Ng853 | n8715));
  assign n1438_1 = ~n7369;
  assign n7371 = (\[1594]  & n8715) | (~Ng441 & (~\[1594]  | n8715));
  assign n1433_1 = ~n7371;
  assign n7373 = (\[1612]  & n8715) | (~Ng438 & (~\[1612]  | n8715));
  assign n1428_1 = ~n7373;
  assign n7375 = (Ng853 & n8716) | (~Ng435 & (~Ng853 | n8716));
  assign n1423_1 = ~n7375;
  assign n7377 = (\[1594]  & n8716) | (~Ng432 & (~\[1594]  | n8716));
  assign n1418_1 = ~n7377;
  assign n7379 = (\[1612]  & n8716) | (~Ng429 & (~\[1612]  | n8716));
  assign n1413 = ~n7379;
  assign n7381 = (Ng1315 & n8717) | (~Ng2571 & (~Ng1315 | n8717));
  assign n6570 = ~n7381;
  assign n7383 = (\[1603]  & n8717) | (~Ng2568 & (~\[1603]  | n8717));
  assign n6565 = ~n7383;
  assign n7385 = (\[1605]  & n8717) | (~Ng2565 & (~\[1605]  | n8717));
  assign n6560 = ~n7385;
  assign n7387 = (~n8718 & n8719) | (~Ng2477 & (n8718 | n8719));
  assign n6048 = ~n7387;
  assign n7389 = (n8719 & ~n8720) | (~Ng2479 & (n8719 | n8720));
  assign n6043 = ~n7389;
  assign n7391 = (n8719 & ~n8721) | (~Ng2478 & (n8719 | n8721));
  assign n6038 = ~n7391;
  assign n7393 = (Ng1315 & n8722) | (~Ng1877 & (~Ng1315 | n8722));
  assign n5063 = ~n7393;
  assign n7395 = (\[1603]  & n8722) | (~Ng1874 & (~\[1603]  | n8722));
  assign n5058 = ~n7395;
  assign n7397 = (\[1605]  & n8722) | (~Ng1871 & (~\[1605]  | n8722));
  assign n5053 = ~n7397;
  assign n7399 = (~n8718 & n8723) | (~Ng1783 & (n8718 | n8723));
  assign n4541 = ~n7399;
  assign n7401 = (~n8720 & n8723) | (~Ng1785 & (n8720 | n8723));
  assign n4536 = ~n7401;
  assign n7403 = (~n8721 & n8723) | (~Ng1784 & (n8721 | n8723));
  assign n4531 = ~n7403;
  assign n7405 = (Ng1315 & n8724) | (~Ng1183 & (~Ng1315 | n8724));
  assign n3556_1 = ~n7405;
  assign n7407 = (\[1603]  & n8724) | (~Ng1180 & (~\[1603]  | n8724));
  assign n3551_1 = ~n7407;
  assign n7409 = (\[1605]  & n8724) | (~Ng1177 & (~\[1605]  | n8724));
  assign n3546_1 = ~n7409;
  assign n7411 = (~n8718 & n8725) | (~Ng1089 & (n8718 | n8725));
  assign n3034_1 = ~n7411;
  assign n7413 = (~n8720 & n8725) | (~Ng1091 & (n8720 | n8725));
  assign n3029_1 = ~n7413;
  assign n7415 = (~n8721 & n8725) | (~Ng1090 & (n8721 | n8725));
  assign n3024_1 = ~n7415;
  assign n7417 = (Ng1315 & n8726) | (~Ng496 & (~Ng1315 | n8726));
  assign n2050_1 = ~n7417;
  assign n7419 = (\[1603]  & n8726) | (~Ng493 & (~\[1603]  | n8726));
  assign n2045_1 = ~n7419;
  assign n7421 = (\[1605]  & n8726) | (~Ng490 & (~\[1605]  | n8726));
  assign n2040 = ~n7421;
  assign n7423 = (~n8718 & n8727) | (~Ng402 & (n8718 | n8727));
  assign n1528 = ~n7423;
  assign n7425 = (~n8720 & n8727) | (~Ng404 & (n8720 | n8727));
  assign n1523_1 = ~n7425;
  assign n7427 = (~n8721 & n8727) | (~Ng403 & (n8721 | n8727));
  assign n1518_1 = ~n7427;
  assign n7429 = (Ng1315 & n6600) | (~Ng3099 & (~Ng1315 | n6600));
  assign n739_1 = ~n7429;
  assign n7431 = (\[1603]  & n6600) | (~Ng3098 & (~\[1603]  | n6600));
  assign n734_1 = ~n7431;
  assign n7433 = (\[1605]  & n6600) | (~Ng3097 & (~\[1605]  | n6600));
  assign n729 = ~n7433;
  assign n7435 = (~n6234 & n8728) | (Pg3234 & (n6234 | n8728));
  assign n7106 = ~n7435;
  assign n7437 = (~n5193 & ~Ng2808) | (~n5191 & (n5193 | ~Ng2808));
  assign n6892 = ~n7437;
  assign n7439 = (~n5188 & ~Ng2810) | (~n5191 & (n5188 | ~Ng2810));
  assign n6887 = ~n7439;
  assign n7441 = (~n5181 & ~Ng2809) | (~n5191 & (n5181 | ~Ng2809));
  assign n6882 = ~n7441;
  assign n7443 = (~Ng2253 & n8729) | (n6149 & (~Ng2253 | ~n8729));
  assign n5610 = ~n7443;
  assign n7445 = (n8730 & ~Ng2255) | (n6149 & (~n8730 | ~Ng2255));
  assign n5605 = ~n7445;
  assign n7447 = (~Ng2254 & n8731) | (n6149 & (~Ng2254 | ~n8731));
  assign n5600 = ~n7447;
  assign n7449 = (~Ng2250 & n8729) | (Ng2165 & (~Ng2250 | ~n8729));
  assign n5595 = ~n7449;
  assign n7451 = (Ng2165 & ~n8730) | (~Ng2252 & (Ng2165 | n8730));
  assign n5590 = ~n7451;
  assign n7453 = (~Ng2251 & n8731) | (Ng2165 & (~Ng2251 | ~n8731));
  assign n5585 = ~n7453;
  assign n7455 = (~Ng2247 & n8729) | (Ng2170 & (~Ng2247 | ~n8729));
  assign n5580 = ~n7455;
  assign n7457 = (Ng2170 & ~n8730) | (~Ng2249 & (Ng2170 | n8730));
  assign n5575 = ~n7457;
  assign n7459 = (~Ng2248 & n8731) | (Ng2170 & (~Ng2248 | ~n8731));
  assign n5570 = ~n7459;
  assign n7461 = (~n8729 & n8732) | (~Ng2244 & (n8729 | n8732));
  assign n5565 = ~n7461;
  assign n7463 = (~n8730 & n8732) | (~Ng2246 & (n8730 | n8732));
  assign n5560 = ~n7463;
  assign n7465 = (~n8731 & n8732) | (~Ng2245 & (n8731 | n8732));
  assign n5555 = ~n7465;
  assign n7467 = (~n5186 & ~Ng2114) | (~n5184 & (n5186 | ~Ng2114));
  assign n5385 = ~n7467;
  assign n7469 = (~n5178 & ~Ng2116) | (~n5184 & (n5178 | ~Ng2116));
  assign n5380 = ~n7469;
  assign n7471 = (~n5171 & ~Ng2115) | (~n5184 & (n5171 | ~Ng2115));
  assign n5375 = ~n7471;
  assign n7473 = (~Ng1559 & n8729) | (n6156 & (~Ng1559 | ~n8729));
  assign n4116_1 = ~n7473;
  assign n7475 = (n8730 & ~Ng1561) | (n6156 & (~n8730 | ~Ng1561));
  assign n4111_1 = ~n7475;
  assign n7477 = (~Ng1560 & n8731) | (n6156 & (~Ng1560 | ~n8731));
  assign n4106 = ~n7477;
  assign n7479 = (~Ng1556 & n8729) | (Ng1471 & (~Ng1556 | ~n8729));
  assign n4101 = ~n7479;
  assign n7481 = (Ng1471 & ~n8730) | (~Ng1558 & (Ng1471 | n8730));
  assign n4096_1 = ~n7481;
  assign n7483 = (~Ng1557 & n8731) | (Ng1471 & (~Ng1557 | ~n8731));
  assign n4091 = ~n7483;
  assign n7485 = (~Ng1553 & n8729) | (Ng1476 & (~Ng1553 | ~n8729));
  assign n4086_1 = ~n7485;
  assign n7487 = (Ng1476 & ~n8730) | (~Ng1555 & (Ng1476 | n8730));
  assign n4081_1 = ~n7487;
  assign n7489 = (~Ng1554 & n8731) | (Ng1476 & (~Ng1554 | ~n8731));
  assign n4076 = ~n7489;
  assign n7491 = (~n8729 & n8733) | (~Ng1550 & (n8729 | n8733));
  assign n4071_1 = ~n7491;
  assign n7493 = (~n8730 & n8733) | (~Ng1552 & (n8730 | n8733));
  assign n4066_1 = ~n7493;
  assign n7495 = (~n8731 & n8733) | (~Ng1551 & (n8731 | n8733));
  assign n4061 = ~n7495;
  assign n7497 = (~n5176 & ~Ng1420) | (~n5174 & (n5176 | ~Ng1420));
  assign n3891 = ~n7497;
  assign n7499 = (~n5168 & ~Ng1422) | (~n5174 & (n5168 | ~Ng1422));
  assign n3886_1 = ~n7499;
  assign n7501 = (~n5161 & ~Ng1421) | (~n5174 & (n5161 | ~Ng1421));
  assign n3881_1 = ~n7501;
  assign n7503 = (~Ng865 & n8729) | (n6163_1 & (~Ng865 | ~n8729));
  assign n2609 = ~n7503;
  assign n7505 = (n8730 & ~Ng867) | (n6163_1 & (~n8730 | ~Ng867));
  assign n2604 = ~n7505;
  assign n7507 = (~Ng866 & n8731) | (n6163_1 & (~Ng866 | ~n8731));
  assign n2599_1 = ~n7507;
  assign n7509 = (~Ng862 & n8729) | (Ng785 & (~Ng862 | ~n8729));
  assign n2594 = ~n7509;
  assign n7511 = (Ng785 & ~n8730) | (~Ng864 & (Ng785 | n8730));
  assign n2589 = ~n7511;
  assign n7513 = (~Ng863 & n8731) | (Ng785 & (~Ng863 | ~n8731));
  assign n2584_1 = ~n7513;
  assign n7515 = (~Ng859 & n8729) | (Ng789 & (~Ng859 | ~n8729));
  assign n2579 = ~n7515;
  assign n7517 = (Ng789 & ~n8730) | (~Ng861 & (Ng789 | n8730));
  assign n2574 = ~n7517;
  assign n7519 = (~Ng860 & n8731) | (Ng789 & (~Ng860 | ~n8731));
  assign n2569 = ~n7519;
  assign n7521 = (~n8729 & n8734) | (~Ng856 & (n8729 | n8734));
  assign n2564 = ~n7521;
  assign n7523 = (~n8730 & n8734) | (~Ng858 & (n8730 | n8734));
  assign n2559 = ~n7523;
  assign n7525 = (~n8731 & n8734) | (~Ng857 & (n8731 | n8734));
  assign n2554 = ~n7525;
  assign n7527 = (~n5166 & ~Ng734) | (~n5164 & (n5166 | ~Ng734));
  assign n2372 = ~n7527;
  assign n7529 = (~n5158 & ~Ng736) | (~n5164 & (n5158 | ~Ng736));
  assign n2367_1 = ~n7529;
  assign n7531 = (~n5154 & ~Ng735) | (~n5164 & (n5154 | ~Ng735));
  assign n2362_1 = ~n7531;
  assign n7533 = (~Ng177 & n8729) | (n6170 & (~Ng177 | ~n8729));
  assign n1103_1 = ~n7533;
  assign n7535 = (n8730 & ~Ng179) | (n6170 & (~n8730 | ~Ng179));
  assign n1098_1 = ~n7535;
  assign n7537 = (~Ng178 & n8731) | (n6170 & (~Ng178 | ~n8731));
  assign n1093_1 = ~n7537;
  assign n7539 = (~Ng174 & n8729) | (Ng97 & (~Ng174 | ~n8729));
  assign n1088_1 = ~n7539;
  assign n7541 = (Ng97 & ~n8730) | (~Ng176 & (Ng97 | n8730));
  assign n1083_1 = ~n7541;
  assign n7543 = (~Ng175 & n8731) | (Ng97 & (~Ng175 | ~n8731));
  assign n1078_1 = ~n7543;
  assign n7545 = (~Ng171 & n8729) | (Ng101 & (~Ng171 | ~n8729));
  assign n1073_1 = ~n7545;
  assign n7547 = (~Ng173 & n8730) | (Ng101 & (~Ng173 | ~n8730));
  assign n1068_1 = ~n7547;
  assign n7549 = (Ng101 & ~n8731) | (~Ng172 & (Ng101 | n8731));
  assign n1063 = ~n7549;
  assign n7551 = (~n8729 & n8735) | (~Ng168 & (n8729 | n8735));
  assign n1058_1 = ~n7551;
  assign n7553 = (~n8730 & n8735) | (~Ng170 & (n8730 | n8735));
  assign n1053 = ~n7553;
  assign n7555 = (~n8731 & n8735) | (~Ng169 & (n8731 | n8735));
  assign n1048 = ~n7555;
  assign n7557 = (Ng1315 & n8736) | (~Ng2676 & (~Ng1315 | n8736));
  assign n6525 = ~n7557;
  assign n7559 = (\[1603]  & n8736) | (~Ng2673 & (~\[1603]  | n8736));
  assign n6520 = ~n7559;
  assign n7561 = (\[1605]  & n8736) | (~Ng2670 & (~\[1605]  | n8736));
  assign n6515 = ~n7561;
  assign n7563 = (Ng1315 & n8737) | (~Ng2667 & (~Ng1315 | n8737));
  assign n6510 = ~n7563;
  assign n7565 = (\[1603]  & n8737) | (~Ng2664 & (~\[1603]  | n8737));
  assign n6505 = ~n7565;
  assign n7567 = (\[1605]  & n8737) | (~Ng2661 & (~\[1605]  | n8737));
  assign n6500 = ~n7567;
  assign n7569 = (~Pg3229 & ~Ng2380) | (Ng2366 & (Pg3229 | ~Ng2380));
  assign n6632 = ~n7569;
  assign n7571 = (Ng2160 & ~n8738) | (n6242 & (~Ng2160 | ~n8738));
  assign n5765 = ~n7571;
  assign n7573 = (Ng1315 & n8739) | (~Ng1982 & (~Ng1315 | n8739));
  assign n5018 = ~n7573;
  assign n7575 = (\[1603]  & n8739) | (~Ng1979 & (~\[1603]  | n8739));
  assign n5013 = ~n7575;
  assign n7577 = (\[1605]  & n8739) | (~Ng1976 & (~\[1605]  | n8739));
  assign n5008 = ~n7577;
  assign n7579 = (Ng1315 & n8740) | (~Ng1973 & (~Ng1315 | n8740));
  assign n5003 = ~n7579;
  assign n7581 = (\[1603]  & n8740) | (~Ng1970 & (~\[1603]  | n8740));
  assign n4998 = ~n7581;
  assign n7583 = (\[1605]  & n8740) | (~Ng1967 & (~\[1605]  | n8740));
  assign n4993 = ~n7583;
  assign n7585 = (~Pg3229 & ~Ng1686) | (Ng1672 & (Pg3229 | ~Ng1686));
  assign n5125 = ~n7585;
  assign n7587 = (Ng1466 & ~n8738) | (n6242 & (~Ng1466 | ~n8738));
  assign n4271 = ~n7587;
  assign n7589 = (Ng1315 & n8741) | (~Ng1288 & (~Ng1315 | n8741));
  assign n3511_1 = ~n7589;
  assign n7591 = (\[1603]  & n8741) | (~Ng1285 & (~\[1603]  | n8741));
  assign n3506_1 = ~n7591;
  assign n7593 = (\[1605]  & n8741) | (~Ng1282 & (~\[1605]  | n8741));
  assign n3501_1 = ~n7593;
  assign n7595 = (Ng1315 & n8742) | (~Ng1279 & (~Ng1315 | n8742));
  assign n3496_1 = ~n7595;
  assign n7597 = (\[1603]  & n8742) | (~Ng1276 & (~\[1603]  | n8742));
  assign n3491_1 = ~n7597;
  assign n7599 = (\[1605]  & n8742) | (~Ng1273 & (~\[1605]  | n8742));
  assign n3486_1 = ~n7599;
  assign n7601 = (~Pg3229 & ~Ng992) | (Ng978 & (Pg3229 | ~Ng992));
  assign n3618_1 = ~n7601;
  assign n7603 = (Ng780 & ~n8738) | (n6242 & (~Ng780 | ~n8738));
  assign n2764_1 = ~n7603;
  assign n7605 = (Ng1315 & n8743) | (~Ng602 & (~Ng1315 | n8743));
  assign n2005_1 = ~n7605;
  assign n7607 = (\[1603]  & n8743) | (~Ng599 & (~\[1603]  | n8743));
  assign n2000_1 = ~n7607;
  assign n7609 = (\[1605]  & n8743) | (~Ng596 & (~\[1605]  | n8743));
  assign n1995_1 = ~n7609;
  assign n7611 = (Ng1315 & n8744) | (~Ng593 & (~Ng1315 | n8744));
  assign n1990_1 = ~n7611;
  assign n7613 = (\[1603]  & n8744) | (~Ng590 & (~\[1603]  | n8744));
  assign n1985 = ~n7613;
  assign n7615 = (\[1605]  & n8744) | (~Ng587 & (~\[1605]  | n8744));
  assign n1980 = ~n7615;
  assign n7617 = (~Pg3229 & ~Ng305) | (Ng291 & (Pg3229 | ~Ng305));
  assign n2112 = ~n7617;
  assign n7619 = (Ng92 & ~n8738) | (n6242 & (~Ng92 | ~n8738));
  assign n1258_1 = ~n7619;
  assign n7621 = ~n8746 & (~Ng3147 | n6537 | ~Ng3097);
  assign n7622 = (~\[1612]  & ~Ng11593) | (n5137 & (\[1612]  | ~Ng11593));
  assign n6341 = ~n7622;
  assign n7624 = (~Ng853 & ~Ng2554) | (n5990 & (Ng853 | ~Ng2554));
  assign n6363 = ~n7624;
  assign n7626 = (\[1594]  & n5990) | (~Ng2553 & (~\[1594]  | n5990));
  assign n6358 = ~n7626;
  assign n7628 = (~\[1612]  & ~Ng2552) | (n5990 & (\[1612]  | ~Ng2552));
  assign n6353 = ~n7628;
  assign n7630 = (~Ng853 & ~Ng11595) | (n6219_1 & (Ng853 | ~Ng11595));
  assign n6391 = ~n7630;
  assign n7632 = (~\[1594]  & ~Ng11594) | (n6219_1 & (\[1594]  | ~Ng11594));
  assign n6387 = ~n7632;
  assign n7634 = (~\[1612]  & ~Ng11598) | (n6219_1 & (\[1612]  | ~Ng11598));
  assign n6383 = ~n7634;
  assign n7636 = (~Ng853 & ~Ng11597) | (n5137 & (Ng853 | ~Ng11597));
  assign n6349 = ~n7636;
  assign n7638 = (~\[1594]  & ~Ng11596) | (n5137 & (\[1594]  | ~Ng11596));
  assign n6345 = ~n7638;
  assign n7640 = (~\[1612]  & ~Ng11566) | (n5135_1 & (\[1612]  | ~Ng11566));
  assign n4834 = ~n7640;
  assign n7642 = (~Ng853 & ~Ng1860) | (n5998_1 & (Ng853 | ~Ng1860));
  assign n4856 = ~n7642;
  assign n7644 = (\[1594]  & n5998_1) | (~Ng1859 & (~\[1594]  | n5998_1));
  assign n4851 = ~n7644;
  assign n7646 = (~\[1612]  & ~Ng1858) | (n5998_1 & (\[1612]  | ~Ng1858));
  assign n4846 = ~n7646;
  assign n7648 = (~Ng853 & ~Ng11568) | (n6223_1 & (Ng853 | ~Ng11568));
  assign n4884 = ~n7648;
  assign n7650 = (~\[1594]  & ~Ng11567) | (n6223_1 & (\[1594]  | ~Ng11567));
  assign n4880 = ~n7650;
  assign n7652 = (~\[1612]  & ~Ng11571) | (n6223_1 & (\[1612]  | ~Ng11571));
  assign n4876 = ~n7652;
  assign n7654 = (~Ng853 & ~Ng11570) | (n5135_1 & (Ng853 | ~Ng11570));
  assign n4842 = ~n7654;
  assign n7656 = (~\[1594]  & ~Ng11569) | (n5135_1 & (\[1594]  | ~Ng11569));
  assign n4838 = ~n7656;
  assign n7658 = (~\[1612]  & ~Ng11539) | (n5131 & (\[1612]  | ~Ng11539));
  assign n3327_1 = ~n7658;
  assign n7660 = (~Ng853 & ~Ng1166) | (n6006 & (Ng853 | ~Ng1166));
  assign n3349_1 = ~n7660;
  assign n7662 = (\[1594]  & n6006) | (~Ng1165 & (~\[1594]  | n6006));
  assign n3344_1 = ~n7662;
  assign n7664 = (~\[1612]  & ~Ng1164) | (n6006 & (\[1612]  | ~Ng1164));
  assign n3339_1 = ~n7664;
  assign n7666 = (~Ng853 & ~Ng11541) | (n6227_1 & (Ng853 | ~Ng11541));
  assign n3377_1 = ~n7666;
  assign n7668 = (~\[1594]  & ~Ng11540) | (n6227_1 & (\[1594]  | ~Ng11540));
  assign n3373_1 = ~n7668;
  assign n7670 = (~\[1612]  & ~Ng11544) | (n6227_1 & (\[1612]  | ~Ng11544));
  assign n3369_1 = ~n7670;
  assign n7672 = (~Ng853 & ~Ng11543) | (n5131 & (Ng853 | ~Ng11543));
  assign n3335_1 = ~n7672;
  assign n7674 = (~\[1594]  & ~Ng11542) | (n5131 & (\[1594]  | ~Ng11542));
  assign n3331_1 = ~n7674;
  assign n7676 = (~\[1612]  & ~Ng11512) | (n5126 & (\[1612]  | ~Ng11512));
  assign n1821_1 = ~n7676;
  assign n7678 = (~Ng853 & ~Ng479) | (n6014 & (Ng853 | ~Ng479));
  assign n1843_1 = ~n7678;
  assign n7680 = (\[1594]  & n6014) | (~Ng478 & (~\[1594]  | n6014));
  assign n1838 = ~n7680;
  assign n7682 = (~\[1612]  & ~Ng477) | (n6014 & (\[1612]  | ~Ng477));
  assign n1833 = ~n7682;
  assign n7684 = (~Ng853 & ~Ng11514) | (n6231_1 & (Ng853 | ~Ng11514));
  assign n1871_1 = ~n7684;
  assign n7686 = (~\[1594]  & ~Ng11513) | (n6231_1 & (\[1594]  | ~Ng11513));
  assign n1867_1 = ~n7686;
  assign n7688 = (~\[1612]  & ~Ng11517) | (n6231_1 & (\[1612]  | ~Ng11517));
  assign n1863 = ~n7688;
  assign n7690 = (~Ng853 & ~Ng11516) | (n5126 & (Ng853 | ~Ng11516));
  assign n1829 = ~n7690;
  assign n7692 = (~\[1594]  & ~Ng11515) | (n5126 & (\[1594]  | ~Ng11515));
  assign n1825_1 = ~n7692;
  assign n7694 = (~Ng853 & ~Ng2563) | (n4908 & (Ng853 | ~Ng2563));
  assign n6336 = ~n7694;
  assign n7696 = (\[1594]  & n4908) | (~Ng2562 & (~\[1594]  | n4908));
  assign n6331 = ~n7696;
  assign n7698 = (~\[1612]  & ~Ng2561) | (n4908 & (\[1612]  | ~Ng2561));
  assign n6326 = ~n7698;
  assign n7700 = (~Ng853 & ~Ng2539) | (~n5034 & (Ng853 | ~Ng2539));
  assign n6378 = ~n7700;
  assign n7702 = (\[1594]  & ~n5034) | (~Ng2559 & (~\[1594]  | ~n5034));
  assign n6373 = ~n7702;
  assign n7704 = (~\[1612]  & ~Ng2555) | (~n5034 & (\[1612]  | ~Ng2555));
  assign n6368 = ~n7704;
  assign n7706 = (n6521 & ~Ng2238) | (~n5044 & (~n6521 | ~Ng2238));
  assign n5550 = ~n7706;
  assign n7708 = (~n5044 & ~n8747) | (~Ng2240 & (~n5044 | n8747));
  assign n5545 = ~n7708;
  assign n7710 = (~Ng2239 & n8748) | (~n5044 & (~Ng2239 | ~n8748));
  assign n5540 = ~n7710;
  assign n7712 = (n6521 & ~Ng2235) | (~n5046 & (~n6521 | ~Ng2235));
  assign n5535 = ~n7712;
  assign n7714 = (~n5046 & ~n8747) | (~Ng2237 & (~n5046 | n8747));
  assign n5530 = ~n7714;
  assign n7716 = (~Ng2236 & n8748) | (~n5046 & (~Ng2236 | ~n8748));
  assign n5525 = ~n7716;
  assign n7718 = (n6521 & ~Ng2232) | (Ng2200 & (~n6521 | ~Ng2232));
  assign n5520 = ~n7718;
  assign n7720 = (Ng2200 & ~n8747) | (~Ng2234 & (Ng2200 | n8747));
  assign n5515 = ~n7720;
  assign n7722 = (~Ng2233 & n8748) | (Ng2200 & (~Ng2233 | ~n8748));
  assign n5510 = ~n7722;
  assign n7724 = (n6521 & ~Ng2229) | (Ng2195 & (~n6521 | ~Ng2229));
  assign n5505 = ~n7724;
  assign n7726 = (Ng2195 & ~n8747) | (~Ng2231 & (Ng2195 | n8747));
  assign n5500 = ~n7726;
  assign n7728 = (~Ng2230 & n8748) | (Ng2195 & (~Ng2230 | ~n8748));
  assign n5495 = ~n7728;
  assign n7730 = (n6521 & ~Ng2226) | (Ng2190 & (~n6521 | ~Ng2226));
  assign n5490 = ~n7730;
  assign n7732 = (Ng2190 & ~n8747) | (~Ng2228 & (Ng2190 | n8747));
  assign n5485 = ~n7732;
  assign n7734 = (~Ng2227 & n8748) | (Ng2190 & (~Ng2227 | ~n8748));
  assign n5480 = ~n7734;
  assign n7736 = (n6521 & ~Ng2223) | (Ng2185 & (~n6521 | ~Ng2223));
  assign n5475 = ~n7736;
  assign n7738 = (Ng2185 & ~n8747) | (~Ng2225 & (Ng2185 | n8747));
  assign n5470 = ~n7738;
  assign n7740 = (~Ng2224 & n8748) | (Ng2185 & (~Ng2224 | ~n8748));
  assign n5465 = ~n7740;
  assign n7742 = (n6521 & ~Ng2220) | (Ng2180 & (~n6521 | ~Ng2220));
  assign n5460 = ~n7742;
  assign n7744 = (Ng2180 & ~n8747) | (~Ng2222 & (Ng2180 | n8747));
  assign n5455 = ~n7744;
  assign n7746 = (~Ng2221 & n8748) | (Ng2180 & (~Ng2221 | ~n8748));
  assign n5450 = ~n7746;
  assign n7748 = (n6521 & ~Ng2217) | (Ng2175 & (~n6521 | ~Ng2217));
  assign n5445 = ~n7748;
  assign n7750 = (~Ng2219 & n8747) | (Ng2175 & (~Ng2219 | ~n8747));
  assign n5440 = ~n7750;
  assign n7752 = (Ng2175 & ~n8748) | (~Ng2218 & (Ng2175 | n8748));
  assign n5435 = ~n7752;
  assign n7754 = (n6521 & ~Ng2208) | (Ng2170 & (~n6521 | ~Ng2208));
  assign n5430 = ~n7754;
  assign n7756 = (Ng2170 & ~n8747) | (~Ng2210 & (Ng2170 | n8747));
  assign n5425 = ~n7756;
  assign n7758 = (~Ng2209 & n8748) | (Ng2170 & (~Ng2209 | ~n8748));
  assign n5420 = ~n7758;
  assign n7760 = (n6521 & ~Ng2205) | (Ng2165 & (~n6521 | ~Ng2205));
  assign n5415 = ~n7760;
  assign n7762 = (Ng2165 & ~n8747) | (~Ng2207 & (Ng2165 | n8747));
  assign n5410 = ~n7762;
  assign n7764 = (~Ng2206 & n8748) | (Ng2165 & (~Ng2206 | ~n8748));
  assign n5405 = ~n7764;
  assign n7766 = (~Ng853 & ~Ng1869) | (n4870 & (Ng853 | ~Ng1869));
  assign n4829 = ~n7766;
  assign n7768 = (\[1594]  & n4870) | (~Ng1868 & (~\[1594]  | n4870));
  assign n4824 = ~n7768;
  assign n7770 = (~\[1612]  & ~Ng1867) | (n4870 & (\[1612]  | ~Ng1867));
  assign n4819 = ~n7770;
  assign n7772 = (~Ng853 & ~Ng1845) | (~n5022 & (Ng853 | ~Ng1845));
  assign n4871_1 = ~n7772;
  assign n7774 = (\[1594]  & ~n5022) | (~Ng1865 & (~\[1594]  | ~n5022));
  assign n4866 = ~n7774;
  assign n7776 = (~\[1612]  & ~Ng1861) | (~n5022 & (\[1612]  | ~Ng1861));
  assign n4861 = ~n7776;
  assign n7778 = (n6521 & ~Ng1544) | (~n5040 & (~n6521 | ~Ng1544));
  assign n4056 = ~n7778;
  assign n7780 = (~n5040 & ~n8747) | (~Ng1546 & (~n5040 | n8747));
  assign n4051 = ~n7780;
  assign n7782 = (~Ng1545 & n8748) | (~n5040 & (~Ng1545 | ~n8748));
  assign n4046 = ~n7782;
  assign n7784 = (n6521 & ~Ng1541) | (~n5042 & (~n6521 | ~Ng1541));
  assign n4041_1 = ~n7784;
  assign n7786 = (~n5042 & ~n8747) | (~Ng1543 & (~n5042 | n8747));
  assign n4036 = ~n7786;
  assign n7788 = (~Ng1542 & n8748) | (~n5042 & (~Ng1542 | ~n8748));
  assign n4031_1 = ~n7788;
  assign n7790 = (n6521 & ~Ng1538) | (Ng1506 & (~n6521 | ~Ng1538));
  assign n4026 = ~n7790;
  assign n7792 = (Ng1506 & ~n8747) | (~Ng1540 & (Ng1506 | n8747));
  assign n4021 = ~n7792;
  assign n7794 = (~Ng1539 & n8748) | (Ng1506 & (~Ng1539 | ~n8748));
  assign n4016_1 = ~n7794;
  assign n7796 = (n6521 & ~Ng1535) | (Ng1501 & (~n6521 | ~Ng1535));
  assign n4011_1 = ~n7796;
  assign n7798 = (Ng1501 & ~n8747) | (~Ng1537 & (Ng1501 | n8747));
  assign n4006_1 = ~n7798;
  assign n7800 = (~Ng1536 & n8748) | (Ng1501 & (~Ng1536 | ~n8748));
  assign n4001_1 = ~n7800;
  assign n7802 = (n6521 & ~Ng1532) | (Ng1496 & (~n6521 | ~Ng1532));
  assign n3996_1 = ~n7802;
  assign n7804 = (Ng1496 & ~n8747) | (~Ng1534 & (Ng1496 | n8747));
  assign n3991 = ~n7804;
  assign n7806 = (~Ng1533 & n8748) | (Ng1496 & (~Ng1533 | ~n8748));
  assign n3986 = ~n7806;
  assign n7808 = (n6521 & ~Ng1529) | (Ng1491 & (~n6521 | ~Ng1529));
  assign n3981 = ~n7808;
  assign n7810 = (Ng1491 & ~n8747) | (~Ng1531 & (Ng1491 | n8747));
  assign n3976 = ~n7810;
  assign n7812 = (~Ng1530 & n8748) | (Ng1491 & (~Ng1530 | ~n8748));
  assign n3971 = ~n7812;
  assign n7814 = (n6521 & ~Ng1526) | (Ng1486 & (~n6521 | ~Ng1526));
  assign n3966 = ~n7814;
  assign n7816 = (~Ng1528 & n8747) | (Ng1486 & (~Ng1528 | ~n8747));
  assign n3961_1 = ~n7816;
  assign n7818 = (Ng1486 & ~n8748) | (~Ng1527 & (Ng1486 | n8748));
  assign n3956 = ~n7818;
  assign n7820 = (n6521 & ~Ng1523) | (Ng1481 & (~n6521 | ~Ng1523));
  assign n3951 = ~n7820;
  assign n7822 = (~Ng1525 & n8747) | (Ng1481 & (~Ng1525 | ~n8747));
  assign n3946 = ~n7822;
  assign n7824 = (Ng1481 & ~n8748) | (~Ng1524 & (Ng1481 | n8748));
  assign n3941_1 = ~n7824;
  assign n7826 = (n6521 & ~Ng1514) | (Ng1476 & (~n6521 | ~Ng1514));
  assign n3936 = ~n7826;
  assign n7828 = (Ng1476 & ~n8747) | (~Ng1516 & (Ng1476 | n8747));
  assign n3931 = ~n7828;
  assign n7830 = (~Ng1515 & n8748) | (Ng1476 & (~Ng1515 | ~n8748));
  assign n3926_1 = ~n7830;
  assign n7832 = (n6521 & ~Ng1511) | (Ng1471 & (~n6521 | ~Ng1511));
  assign n3921 = ~n7832;
  assign n7834 = (Ng1471 & ~n8747) | (~Ng1513 & (Ng1471 | n8747));
  assign n3916_1 = ~n7834;
  assign n7836 = (~Ng1512 & n8748) | (Ng1471 & (~Ng1512 | ~n8748));
  assign n3911 = ~n7836;
  assign n7838 = (~Ng853 & ~Ng1175) | (n4828 & (Ng853 | ~Ng1175));
  assign n3322_1 = ~n7838;
  assign n7840 = (\[1594]  & n4828) | (~Ng1174 & (~\[1594]  | n4828));
  assign n3317_1 = ~n7840;
  assign n7842 = (~\[1612]  & ~Ng1173) | (n4828 & (\[1612]  | ~Ng1173));
  assign n3312_1 = ~n7842;
  assign n7844 = (~Ng853 & ~Ng1151) | (~n5010 & (Ng853 | ~Ng1151));
  assign n3364_1 = ~n7844;
  assign n7846 = (\[1594]  & ~n5010) | (~Ng1171 & (~\[1594]  | ~n5010));
  assign n3359_1 = ~n7846;
  assign n7848 = (~\[1612]  & ~Ng1167) | (~n5010 & (\[1612]  | ~Ng1167));
  assign n3354_1 = ~n7848;
  assign n7850 = (n6521 & ~Ng850) | (~n5032 & (~n6521 | ~Ng850));
  assign n2549 = ~n7850;
  assign n7852 = (~n5032 & ~n8747) | (~Ng852 & (~n5032 | n8747));
  assign n2544 = ~n7852;
  assign n7854 = (~Ng851 & n8748) | (~n5032 & (~Ng851 | ~n8748));
  assign n2539 = ~n7854;
  assign n7856 = (n6521 & ~Ng847) | (~n5038_1 & (~n6521 | ~Ng847));
  assign n2534_1 = ~n7856;
  assign n7858 = (~n5038_1 & ~n8747) | (~Ng849 & (~n5038_1 | n8747));
  assign n2529 = ~n7858;
  assign n7860 = (~Ng848 & n8748) | (~n5038_1 & (~Ng848 | ~n8748));
  assign n2524_1 = ~n7860;
  assign n7862 = (n6521 & ~Ng844) | (Ng813 & (~n6521 | ~Ng844));
  assign n2519_1 = ~n7862;
  assign n7864 = (Ng813 & ~n8747) | (~Ng846 & (Ng813 | n8747));
  assign n2514_1 = ~n7864;
  assign n7866 = (~Ng845 & n8748) | (Ng813 & (~Ng845 | ~n8748));
  assign n2509 = ~n7866;
  assign n7868 = (n6521 & ~Ng841) | (Ng809 & (~n6521 | ~Ng841));
  assign n2504_1 = ~n7868;
  assign n7870 = (Ng809 & ~n8747) | (~Ng843 & (Ng809 | n8747));
  assign n2499_1 = ~n7870;
  assign n7872 = (~Ng842 & n8748) | (Ng809 & (~Ng842 | ~n8748));
  assign n2494 = ~n7872;
  assign n7874 = (n6521 & ~Ng838) | (Ng805 & (~n6521 | ~Ng838));
  assign n2489_1 = ~n7874;
  assign n7876 = (Ng805 & ~n8747) | (~Ng840 & (Ng805 | n8747));
  assign n2484 = ~n7876;
  assign n7878 = (~Ng839 & n8748) | (Ng805 & (~Ng839 | ~n8748));
  assign n2479 = ~n7878;
  assign n7880 = (n6521 & ~Ng835) | (Ng801 & (~n6521 | ~Ng835));
  assign n2474 = ~n7880;
  assign n7882 = (~Ng837 & n8747) | (Ng801 & (~Ng837 | ~n8747));
  assign n2469 = ~n7882;
  assign n7884 = (Ng801 & ~n8748) | (~Ng836 & (Ng801 | n8748));
  assign n2464 = ~n7884;
  assign n7886 = (n6521 & ~Ng832) | (Ng797 & (~n6521 | ~Ng832));
  assign n2459 = ~n7886;
  assign n7888 = (~Ng834 & n8747) | (Ng797 & (~Ng834 | ~n8747));
  assign n2454 = ~n7888;
  assign n7890 = (Ng797 & ~n8748) | (~Ng833 & (Ng797 | n8748));
  assign n2449 = ~n7890;
  assign n7892 = (n6521 & ~Ng829) | (Ng793 & (~n6521 | ~Ng829));
  assign n2444_1 = ~n7892;
  assign n7894 = (~Ng831 & n8747) | (Ng793 & (~Ng831 | ~n8747));
  assign n2439 = ~n7894;
  assign n7896 = (Ng793 & ~n8748) | (~Ng830 & (Ng793 | n8748));
  assign n2434 = ~n7896;
  assign n7898 = (n6521 & ~Ng820) | (Ng789 & (~n6521 | ~Ng820));
  assign n2429_1 = ~n7898;
  assign n7900 = (Ng789 & ~n8747) | (~Ng822 & (Ng789 | n8747));
  assign n2424_1 = ~n7900;
  assign n7902 = (~Ng821 & n8748) | (Ng789 & (~Ng821 | ~n8748));
  assign n2419 = ~n7902;
  assign n7904 = (n6521 & ~Ng817) | (Ng785 & (~n6521 | ~Ng817));
  assign n2414 = ~n7904;
  assign n7906 = (Ng785 & ~n8747) | (~Ng819 & (Ng785 | n8747));
  assign n2409 = ~n7906;
  assign n7908 = (~Ng818 & n8748) | (Ng785 & (~Ng818 | ~n8748));
  assign n2404 = ~n7908;
  assign n7910 = (~Ng853 & ~Ng488) | (n4786 & (Ng853 | ~Ng488));
  assign n1816_1 = ~n7910;
  assign n7912 = (\[1594]  & n4786) | (~Ng487 & (~\[1594]  | n4786));
  assign n1811_1 = ~n7912;
  assign n7914 = (~\[1612]  & ~Ng486) | (n4786 & (\[1612]  | ~Ng486));
  assign n1806_1 = ~n7914;
  assign n7916 = (~Ng853 & ~Ng464) | (~n4998_1 & (Ng853 | ~Ng464));
  assign n1858_1 = ~n7916;
  assign n7918 = (\[1594]  & ~n4998_1) | (~Ng484 & (~\[1594]  | ~n4998_1));
  assign n1853_1 = ~n7918;
  assign n7920 = (~\[1612]  & ~Ng480) | (~n4998_1 & (\[1612]  | ~Ng480));
  assign n1848 = ~n7920;
  assign n7922 = (n6521 & ~Ng162) | (~n5020 & (~n6521 | ~Ng162));
  assign n1043_1 = ~n7922;
  assign n7924 = (~n5020 & ~n8747) | (~Ng164 & (~n5020 | n8747));
  assign n1038_1 = ~n7924;
  assign n7926 = (~Ng163 & n8748) | (~n5020 & (~Ng163 | ~n8748));
  assign n1033 = ~n7926;
  assign n7928 = (n6521 & ~Ng159) | (~n5030 & (~n6521 | ~Ng159));
  assign n1028_1 = ~n7928;
  assign n7930 = (~n5030 & ~n8747) | (~Ng161 & (~n5030 | n8747));
  assign n1023_1 = ~n7930;
  assign n7932 = (~Ng160 & n8748) | (~n5030 & (~Ng160 | ~n8748));
  assign n1018 = ~n7932;
  assign n7934 = (n6521 & ~Ng156) | (Ng125 & (~n6521 | ~Ng156));
  assign n1013_1 = ~n7934;
  assign n7936 = (Ng125 & ~n8747) | (~Ng158 & (Ng125 | n8747));
  assign n1008_1 = ~n7936;
  assign n7938 = (~Ng157 & n8748) | (Ng125 & (~Ng157 | ~n8748));
  assign n1003 = ~n7938;
  assign n7940 = (n6521 & ~Ng153) | (Ng121 & (~n6521 | ~Ng153));
  assign n998 = ~n7940;
  assign n7942 = (Ng121 & ~n8747) | (~Ng155 & (Ng121 | n8747));
  assign n993_1 = ~n7942;
  assign n7944 = (~Ng154 & n8748) | (Ng121 & (~Ng154 | ~n8748));
  assign n988_1 = ~n7944;
  assign n7946 = (n6521 & ~Ng150) | (Ng117 & (~n6521 | ~Ng150));
  assign n983_1 = ~n7946;
  assign n7948 = (~Ng152 & n8747) | (Ng117 & (~Ng152 | ~n8747));
  assign n978_1 = ~n7948;
  assign n7950 = (Ng117 & ~n8748) | (~Ng151 & (Ng117 | n8748));
  assign n973_1 = ~n7950;
  assign n7952 = (n6521 & ~Ng147) | (Ng113 & (~n6521 | ~Ng147));
  assign n968_1 = ~n7952;
  assign n7954 = (~Ng149 & n8747) | (Ng113 & (~Ng149 | ~n8747));
  assign n963_1 = ~n7954;
  assign n7956 = (Ng113 & ~n8748) | (~Ng148 & (Ng113 | n8748));
  assign n958 = ~n7956;
  assign n7958 = (n6521 & ~Ng144) | (Ng109 & (~n6521 | ~Ng144));
  assign n953_1 = ~n7958;
  assign n7960 = (~Ng146 & n8747) | (Ng109 & (~Ng146 | ~n8747));
  assign n948_1 = ~n7960;
  assign n7962 = (Ng109 & ~n8748) | (~Ng145 & (Ng109 | n8748));
  assign n943_1 = ~n7962;
  assign n7964 = (n6521 & ~Ng141) | (Ng105 & (~n6521 | ~Ng141));
  assign n938_1 = ~n7964;
  assign n7966 = (~Ng143 & n8747) | (Ng105 & (~Ng143 | ~n8747));
  assign n933_1 = ~n7966;
  assign n7968 = (Ng105 & ~n8748) | (~Ng142 & (Ng105 | n8748));
  assign n928 = ~n7968;
  assign n7970 = (n6521 & ~Ng132) | (Ng101 & (~n6521 | ~Ng132));
  assign n923_1 = ~n7970;
  assign n7972 = (Ng101 & ~n8747) | (~Ng134 & (Ng101 | n8747));
  assign n918_1 = ~n7972;
  assign n7974 = (~Ng133 & n8748) | (Ng101 & (~Ng133 | ~n8748));
  assign n913_1 = ~n7974;
  assign n7976 = (n6521 & ~Ng129) | (Ng97 & (~n6521 | ~Ng129));
  assign n908_1 = ~n7976;
  assign n7978 = (Ng97 & ~n8747) | (~Ng131 & (Ng97 | n8747));
  assign n903_1 = ~n7978;
  assign n7980 = (~Ng130 & n8748) | (Ng97 & (~Ng130 | ~n8748));
  assign n898_1 = ~n7980;
  assign n7982 = (~Ng2879 & n8749) | (~Pg8096 & (Ng2879 | n8749));
  assign n616 = ~n7982;
  assign n7984 = (Ng2879 & ~n8763) | (~Ng13455 & (~Ng2879 | ~n8763));
  assign n664_1 = ~n7984;
  assign n7986 = (~Ng2879 & ~Ng13439) | (n8749 & (Ng2879 | ~Ng13439));
  assign n475_1 = ~n7986;
  assign n7988 = (~Ng2879 & ~n8763) | (~Pg7519 & (Ng2879 | ~n8763));
  assign n544_1 = ~n7988;
  assign n7990 = (n5192 & ~Ng2805) | (~n5064 & (~n5192 | ~Ng2805));
  assign n6877 = ~n7990;
  assign n7992 = (~n5064 & ~n5115_1) | (~Ng2807 & (~n5064 | n5115_1));
  assign n6872 = ~n7992;
  assign n7994 = (n5180_1 & ~Ng2806) | (~n5064 & (~n5180_1 | ~Ng2806));
  assign n6867 = ~n7994;
  assign n7996 = (n5192 & ~Ng2802) | (~n4982 & (~n5192 | ~Ng2802));
  assign n6862 = ~n7996;
  assign n7998 = (n5115_1 & ~Ng2804) | (~n4982 & (~n5115_1 | ~Ng2804));
  assign n6857 = ~n7998;
  assign n8000 = (n5180_1 & ~Ng2803) | (~n4982 & (~n5180_1 | ~Ng2803));
  assign n6852 = ~n8000;
  assign n8002 = (~n5193 & ~Ng2799) | (Ng2766 & (n5193 | ~Ng2799));
  assign n6847 = ~n8002;
  assign n8004 = (n5188 & Ng2766) | (~Ng2801 & (~n5188 | Ng2766));
  assign n6842 = ~n8004;
  assign n8006 = (~n5181 & ~Ng2800) | (Ng2766 & (n5181 | ~Ng2800));
  assign n6837 = ~n8006;
  assign n8008 = (~n5193 & ~Ng2796) | (Ng2760 & (n5193 | ~Ng2796));
  assign n6832 = ~n8008;
  assign n8010 = (n5188 & Ng2760) | (~Ng2798 & (~n5188 | Ng2760));
  assign n6827 = ~n8010;
  assign n8012 = (~n5181 & ~Ng2797) | (Ng2760 & (n5181 | ~Ng2797));
  assign n6822 = ~n8012;
  assign n8014 = (~n5193 & ~Ng2793) | (Ng2753 & (n5193 | ~Ng2793));
  assign n6817 = ~n8014;
  assign n8016 = (n5188 & Ng2753) | (~Ng2795 & (~n5188 | Ng2753));
  assign n6812 = ~n8016;
  assign n8018 = (~n5181 & ~Ng2794) | (Ng2753 & (n5181 | ~Ng2794));
  assign n6807 = ~n8018;
  assign n8020 = (~n5193 & ~Ng2790) | (Ng2740 & (n5193 | ~Ng2790));
  assign n6802 = ~n8020;
  assign n8022 = (n5188 & Ng2740) | (~Ng2792 & (~n5188 | Ng2740));
  assign n6797 = ~n8022;
  assign n8024 = (~n5181 & ~Ng2791) | (Ng2740 & (n5181 | ~Ng2791));
  assign n6792 = ~n8024;
  assign n8026 = (~n5193 & ~Ng2787) | (Ng2746 & (n5193 | ~Ng2787));
  assign n6787 = ~n8026;
  assign n8028 = (n5188 & Ng2746) | (~Ng2789 & (~n5188 | Ng2746));
  assign n6782 = ~n8028;
  assign n8030 = (~n5181 & ~Ng2788) | (Ng2746 & (n5181 | ~Ng2788));
  assign n6777 = ~n8030;
  assign n8032 = (~n5193 & ~Ng2784) | (Ng2734 & (n5193 | ~Ng2784));
  assign n6772 = ~n8032;
  assign n8034 = (n5188 & Ng2734) | (~Ng2786 & (~n5188 | Ng2734));
  assign n6767 = ~n8034;
  assign n8036 = (~n5181 & ~Ng2785) | (Ng2734 & (n5181 | ~Ng2785));
  assign n6762 = ~n8036;
  assign n8038 = (~n5193 & ~Ng2781) | (Ng2720 & (n5193 | ~Ng2781));
  assign n6757 = ~n8038;
  assign n8040 = (n5188 & Ng2720) | (~Ng2783 & (~n5188 | Ng2720));
  assign n6752 = ~n8040;
  assign n8042 = (~n5181 & ~Ng2782) | (Ng2720 & (n5181 | ~Ng2782));
  assign n6747 = ~n8042;
  assign n8044 = (~n5193 & ~Ng2778) | (Ng2727 & (n5193 | ~Ng2778));
  assign n6742 = ~n8044;
  assign n8046 = (n5188 & Ng2727) | (~Ng2780 & (~n5188 | Ng2727));
  assign n6737 = ~n8046;
  assign n8048 = (~n5181 & ~Ng2779) | (Ng2727 & (n5181 | ~Ng2779));
  assign n6732 = ~n8048;
  assign n8050 = (~n5193 & ~Ng2775) | (Ng2707 & (n5193 | ~Ng2775));
  assign n6727 = ~n8050;
  assign n8052 = (n5188 & Ng2707) | (~Ng2777 & (~n5188 | Ng2707));
  assign n6722 = ~n8052;
  assign n8054 = (~n5181 & ~Ng2776) | (Ng2707 & (n5181 | ~Ng2776));
  assign n6717 = ~n8054;
  assign n8056 = (~n5193 & ~Ng2772) | (Ng2714 & (n5193 | ~Ng2772));
  assign n6712 = ~n8056;
  assign n8058 = (n5188 & Ng2714) | (~Ng2774 & (~n5188 | Ng2714));
  assign n6707 = ~n8058;
  assign n8060 = (~n5181 & ~Ng2773) | (Ng2714 & (n5181 | ~Ng2773));
  assign n6702 = ~n8060;
  assign n8062 = (n5185_1 & ~Ng2111) | (~n5062 & (~n5185_1 | ~Ng2111));
  assign n5370 = ~n8062;
  assign n8064 = (~n5062 & ~n5112) | (~Ng2113 & (~n5062 | n5112));
  assign n5365 = ~n8064;
  assign n8066 = (n5170_1 & ~Ng2112) | (~n5062 & (~n5170_1 | ~Ng2112));
  assign n5360 = ~n8066;
  assign n8068 = (n5185_1 & ~Ng2108) | (~n4978_1 & (~n5185_1 | ~Ng2108));
  assign n5355 = ~n8068;
  assign n8070 = (n5112 & ~Ng2110) | (~n4978_1 & (~n5112 | ~Ng2110));
  assign n5350 = ~n8070;
  assign n8072 = (n5170_1 & ~Ng2109) | (~n4978_1 & (~n5170_1 | ~Ng2109));
  assign n5345 = ~n8072;
  assign n8074 = (~n5186 & ~Ng2105) | (Ng2072 & (n5186 | ~Ng2105));
  assign n5340 = ~n8074;
  assign n8076 = (n5178 & Ng2072) | (~Ng2107 & (~n5178 | Ng2072));
  assign n5335 = ~n8076;
  assign n8078 = (~n5171 & ~Ng2106) | (Ng2072 & (n5171 | ~Ng2106));
  assign n5330 = ~n8078;
  assign n8080 = (~n5186 & ~Ng2102) | (Ng2066 & (n5186 | ~Ng2102));
  assign n5325 = ~n8080;
  assign n8082 = (n5178 & Ng2066) | (~Ng2104 & (~n5178 | Ng2066));
  assign n5320 = ~n8082;
  assign n8084 = (~n5171 & ~Ng2103) | (Ng2066 & (n5171 | ~Ng2103));
  assign n5315 = ~n8084;
  assign n8086 = (~n5186 & ~Ng2099) | (Ng2059 & (n5186 | ~Ng2099));
  assign n5310 = ~n8086;
  assign n8088 = (n5178 & Ng2059) | (~Ng2101 & (~n5178 | Ng2059));
  assign n5305 = ~n8088;
  assign n8090 = (~n5171 & ~Ng2100) | (Ng2059 & (n5171 | ~Ng2100));
  assign n5300 = ~n8090;
  assign n8092 = (~n5186 & ~Ng2096) | (Ng2046 & (n5186 | ~Ng2096));
  assign n5295 = ~n8092;
  assign n8094 = (n5178 & Ng2046) | (~Ng2098 & (~n5178 | Ng2046));
  assign n5290 = ~n8094;
  assign n8096 = (~n5171 & ~Ng2097) | (Ng2046 & (n5171 | ~Ng2097));
  assign n5285 = ~n8096;
  assign n8098 = (~n5186 & ~Ng2093) | (Ng2052 & (n5186 | ~Ng2093));
  assign n5280 = ~n8098;
  assign n8100 = (n5178 & Ng2052) | (~Ng2095 & (~n5178 | Ng2052));
  assign n5275 = ~n8100;
  assign n8102 = (~n5171 & ~Ng2094) | (Ng2052 & (n5171 | ~Ng2094));
  assign n5270 = ~n8102;
  assign n8104 = (~n5186 & ~Ng2090) | (Ng2040 & (n5186 | ~Ng2090));
  assign n5265 = ~n8104;
  assign n8106 = (n5178 & Ng2040) | (~Ng2092 & (~n5178 | Ng2040));
  assign n5260 = ~n8106;
  assign n8108 = (~n5171 & ~Ng2091) | (Ng2040 & (n5171 | ~Ng2091));
  assign n5255 = ~n8108;
  assign n8110 = (~n5186 & ~Ng2087) | (Ng2026 & (n5186 | ~Ng2087));
  assign n5250 = ~n8110;
  assign n8112 = (n5178 & Ng2026) | (~Ng2089 & (~n5178 | Ng2026));
  assign n5245 = ~n8112;
  assign n8114 = (~n5171 & ~Ng2088) | (Ng2026 & (n5171 | ~Ng2088));
  assign n5240 = ~n8114;
  assign n8116 = (~n5186 & ~Ng2084) | (Ng2033 & (n5186 | ~Ng2084));
  assign n5235 = ~n8116;
  assign n8118 = (n5178 & Ng2033) | (~Ng2086 & (~n5178 | Ng2033));
  assign n5230 = ~n8118;
  assign n8120 = (~n5171 & ~Ng2085) | (Ng2033 & (n5171 | ~Ng2085));
  assign n5225 = ~n8120;
  assign n8122 = (~n5186 & ~Ng2081) | (Ng2013 & (n5186 | ~Ng2081));
  assign n5220 = ~n8122;
  assign n8124 = (n5178 & Ng2013) | (~Ng2083 & (~n5178 | Ng2013));
  assign n5215 = ~n8124;
  assign n8126 = (~n5171 & ~Ng2082) | (Ng2013 & (n5171 | ~Ng2082));
  assign n5210 = ~n8126;
  assign n8128 = (~n5186 & ~Ng2078) | (Ng2020 & (n5186 | ~Ng2078));
  assign n5205 = ~n8128;
  assign n8130 = (n5178 & Ng2020) | (~Ng2080 & (~n5178 | Ng2020));
  assign n5200 = ~n8130;
  assign n8132 = (~n5171 & ~Ng2079) | (Ng2020 & (n5171 | ~Ng2079));
  assign n5195 = ~n8132;
  assign n8134 = (n5175_1 & ~Ng1417) | (~n5058_1 & (~n5175_1 | ~Ng1417));
  assign n3876_1 = ~n8134;
  assign n8136 = (~n5058_1 & ~n5109) | (~Ng1419 & (~n5058_1 | n5109));
  assign n3871_1 = ~n8136;
  assign n8138 = (n5160_1 & ~Ng1418) | (~n5058_1 & (~n5160_1 | ~Ng1418));
  assign n3866 = ~n8138;
  assign n8140 = (n5175_1 & ~Ng1414) | (~n4972 & (~n5175_1 | ~Ng1414));
  assign n3861_1 = ~n8140;
  assign n8142 = (n5109 & ~Ng1416) | (~n4972 & (~n5109 | ~Ng1416));
  assign n3856_1 = ~n8142;
  assign n8144 = (n5160_1 & ~Ng1415) | (~n4972 & (~n5160_1 | ~Ng1415));
  assign n3851_1 = ~n8144;
  assign n8146 = (~n5176 & ~Ng1411) | (Ng1378 & (n5176 | ~Ng1411));
  assign n3846_1 = ~n8146;
  assign n8148 = (n5168 & Ng1378) | (~Ng1413 & (~n5168 | Ng1378));
  assign n3841_1 = ~n8148;
  assign n8150 = (~n5161 & ~Ng1412) | (Ng1378 & (n5161 | ~Ng1412));
  assign n3836_1 = ~n8150;
  assign n8152 = (~n5176 & ~Ng1408) | (Ng1372 & (n5176 | ~Ng1408));
  assign n3831_1 = ~n8152;
  assign n8154 = (n5168 & Ng1372) | (~Ng1410 & (~n5168 | Ng1372));
  assign n3826_1 = ~n8154;
  assign n8156 = (~n5161 & ~Ng1409) | (Ng1372 & (n5161 | ~Ng1409));
  assign n3821 = ~n8156;
  assign n8158 = (~n5176 & ~Ng1405) | (Ng1365 & (n5176 | ~Ng1405));
  assign n3816 = ~n8158;
  assign n8160 = (n5168 & Ng1365) | (~Ng1407 & (~n5168 | Ng1365));
  assign n3811_1 = ~n8160;
  assign n8162 = (~n5161 & ~Ng1406) | (Ng1365 & (n5161 | ~Ng1406));
  assign n3806 = ~n8162;
  assign n8164 = (~n5176 & ~Ng1402) | (Ng1352 & (n5176 | ~Ng1402));
  assign n3801 = ~n8164;
  assign n8166 = (n5168 & Ng1352) | (~Ng1404 & (~n5168 | Ng1352));
  assign n3796_1 = ~n8166;
  assign n8168 = (~n5161 & ~Ng1403) | (Ng1352 & (n5161 | ~Ng1403));
  assign n3791 = ~n8168;
  assign n8170 = (~n5176 & ~Ng1399) | (Ng1358 & (n5176 | ~Ng1399));
  assign n3786 = ~n8170;
  assign n8172 = (n5168 & Ng1358) | (~Ng1401 & (~n5168 | Ng1358));
  assign n3781_1 = ~n8172;
  assign n8174 = (~n5161 & ~Ng1400) | (Ng1358 & (n5161 | ~Ng1400));
  assign n3776_1 = ~n8174;
  assign n8176 = (~n5176 & ~Ng1396) | (Ng1346 & (n5176 | ~Ng1396));
  assign n3771 = ~n8176;
  assign n8178 = (n5168 & Ng1346) | (~Ng1398 & (~n5168 | Ng1346));
  assign n3766_1 = ~n8178;
  assign n8180 = (~n5161 & ~Ng1397) | (Ng1346 & (n5161 | ~Ng1397));
  assign n3761 = ~n8180;
  assign n8182 = (~n5176 & ~Ng1393) | (Ng1332 & (n5176 | ~Ng1393));
  assign n3756_1 = ~n8182;
  assign n8184 = (n5168 & Ng1332) | (~Ng1395 & (~n5168 | Ng1332));
  assign n3751_1 = ~n8184;
  assign n8186 = (~n5161 & ~Ng1394) | (Ng1332 & (n5161 | ~Ng1394));
  assign n3746_1 = ~n8186;
  assign n8188 = (~n5176 & ~Ng1390) | (Ng1339 & (n5176 | ~Ng1390));
  assign n3741_1 = ~n8188;
  assign n8190 = (n5168 & Ng1339) | (~Ng1392 & (~n5168 | Ng1339));
  assign n3736_1 = ~n8190;
  assign n8192 = (~n5161 & ~Ng1391) | (Ng1339 & (n5161 | ~Ng1391));
  assign n3731_1 = ~n8192;
  assign n8194 = (~n5176 & ~Ng1387) | (Ng1319 & (n5176 | ~Ng1387));
  assign n3726_1 = ~n8194;
  assign n8196 = (n5168 & Ng1319) | (~Ng1389 & (~n5168 | Ng1319));
  assign n3721_1 = ~n8196;
  assign n8198 = (~n5161 & ~Ng1388) | (Ng1319 & (n5161 | ~Ng1388));
  assign n3716_1 = ~n8198;
  assign n8200 = (~n5176 & ~Ng1384) | (Ng1326 & (n5176 | ~Ng1384));
  assign n3711_1 = ~n8200;
  assign n8202 = (n5168 & Ng1326) | (~Ng1386 & (~n5168 | Ng1326));
  assign n3706_1 = ~n8202;
  assign n8204 = (~n5161 & ~Ng1385) | (Ng1326 & (n5161 | ~Ng1385));
  assign n3701_1 = ~n8204;
  assign n8206 = (n5165_1 & ~Ng731) | (~n5054 & (~n5165_1 | ~Ng731));
  assign n2357 = ~n8206;
  assign n8208 = (~n5054 & ~n5106) | (~Ng733 & (~n5054 | n5106));
  assign n2352 = ~n8208;
  assign n8210 = (n5153 & ~Ng732) | (~n5054 & (~n5153 | ~Ng732));
  assign n2347 = ~n8210;
  assign n8212 = (n5165_1 & ~Ng728) | (~n4964 & (~n5165_1 | ~Ng728));
  assign n2342 = ~n8212;
  assign n8214 = (n5106 & ~Ng730) | (~n4964 & (~n5106 | ~Ng730));
  assign n2337 = ~n8214;
  assign n8216 = (n5153 & ~Ng729) | (~n4964 & (~n5153 | ~Ng729));
  assign n2332_1 = ~n8216;
  assign n8218 = (~n5166 & ~Ng725) | (Ng692 & (n5166 | ~Ng725));
  assign n2327_1 = ~n8218;
  assign n8220 = (n5158 & Ng692) | (~Ng727 & (~n5158 | Ng692));
  assign n2322 = ~n8220;
  assign n8222 = (~n5154 & ~Ng726) | (Ng692 & (n5154 | ~Ng726));
  assign n2317 = ~n8222;
  assign n8224 = (~n5166 & ~Ng722) | (Ng686 & (n5166 | ~Ng722));
  assign n2312 = ~n8224;
  assign n8226 = (n5158 & Ng686) | (~Ng724 & (~n5158 | Ng686));
  assign n2307 = ~n8226;
  assign n8228 = (~n5154 & ~Ng723) | (Ng686 & (n5154 | ~Ng723));
  assign n2302 = ~n8228;
  assign n8230 = (~n5166 & ~Ng719) | (Ng679 & (n5166 | ~Ng719));
  assign n2297_1 = ~n8230;
  assign n8232 = (n5158 & Ng679) | (~Ng721 & (~n5158 | Ng679));
  assign n2292 = ~n8232;
  assign n8234 = (~n5154 & ~Ng720) | (Ng679 & (n5154 | ~Ng720));
  assign n2287 = ~n8234;
  assign n8236 = (~n5166 & ~Ng716) | (Ng666 & (n5166 | ~Ng716));
  assign n2282 = ~n8236;
  assign n8238 = (n5158 & Ng666) | (~Ng718 & (~n5158 | Ng666));
  assign n2277 = ~n8238;
  assign n8240 = (~n5154 & ~Ng717) | (Ng666 & (n5154 | ~Ng717));
  assign n2272 = ~n8240;
  assign n8242 = (~n5166 & ~Ng713) | (Ng672 & (n5166 | ~Ng713));
  assign n2267 = ~n8242;
  assign n8244 = (n5158 & Ng672) | (~Ng715 & (~n5158 | Ng672));
  assign n2262 = ~n8244;
  assign n8246 = (~n5154 & ~Ng714) | (Ng672 & (n5154 | ~Ng714));
  assign n2257_1 = ~n8246;
  assign n8248 = (~n5166 & ~Ng710) | (Ng660 & (n5166 | ~Ng710));
  assign n2252 = ~n8248;
  assign n8250 = (n5158 & Ng660) | (~Ng712 & (~n5158 | Ng660));
  assign n2247_1 = ~n8250;
  assign n8252 = (~n5154 & ~Ng711) | (Ng660 & (n5154 | ~Ng711));
  assign n2242 = ~n8252;
  assign n8254 = (~n5166 & ~Ng707) | (Ng646 & (n5166 | ~Ng707));
  assign n2237_1 = ~n8254;
  assign n8256 = (n5158 & Ng646) | (~Ng709 & (~n5158 | Ng646));
  assign n2232 = ~n8256;
  assign n8258 = (~n5154 & ~Ng708) | (Ng646 & (n5154 | ~Ng708));
  assign n2227_1 = ~n8258;
  assign n8260 = (~n5166 & ~Ng704) | (Ng653 & (n5166 | ~Ng704));
  assign n2222 = ~n8260;
  assign n8262 = (n5158 & Ng653) | (~Ng706 & (~n5158 | Ng653));
  assign n2217_1 = ~n8262;
  assign n8264 = (~n5154 & ~Ng705) | (Ng653 & (n5154 | ~Ng705));
  assign n2212_1 = ~n8264;
  assign n8266 = (~n5166 & ~Ng701) | (Ng633 & (n5166 | ~Ng701));
  assign n2207_1 = ~n8266;
  assign n8268 = (n5158 & Ng633) | (~Ng703 & (~n5158 | Ng633));
  assign n2202 = ~n8268;
  assign n8270 = (~n5154 & ~Ng702) | (Ng633 & (n5154 | ~Ng702));
  assign n2197 = ~n8270;
  assign n8272 = (~n5166 & ~Ng698) | (Ng640 & (n5166 | ~Ng698));
  assign n2192_1 = ~n8272;
  assign n8274 = (n5158 & Ng640) | (~Ng700 & (~n5158 | Ng640));
  assign n2187_1 = ~n8274;
  assign n8276 = (~n5154 & ~Ng699) | (Ng640 & (n5154 | ~Ng699));
  assign n2182_1 = ~n8276;
  assign n8278 = (~Ng2879 & ~Ng2975) | (~Pg4590 & (Ng2879 | ~Ng2975));
  assign n504_1 = ~n8278;
  assign n8280 = (~Ng2879 & ~Ng2978) | (~Pg4323 & (Ng2879 | ~Ng2978));
  assign n496_1 = ~n8280;
  assign n8282 = (~Ng2879 & ~Ng2981) | (~Pg4090 & (Ng2879 | ~Ng2981));
  assign n488_1 = ~n8282;
  assign n8284 = (~Ng2879 & ~Ng2874) | (~Pg8251 & (Ng2879 | ~Ng2874));
  assign n480_1 = ~n8284;
  assign n8286 = (~Ng2879 & ~Ng2935) | (~Pg4450 & (Ng2879 | ~Ng2935));
  assign n608_1 = ~n8286;
  assign n8288 = (~Ng2879 & ~Ng2938) | (~Pg4200 & (Ng2879 | ~Ng2938));
  assign n600_1 = ~n8288;
  assign n8290 = (~Ng2879 & ~Ng2941) | (~Pg3993 & (Ng2879 | ~Ng2941));
  assign n592_1 = ~n8290;
  assign n8292 = (~Ng2879 & ~Ng2944) | (~Pg8175 & (Ng2879 | ~Ng2944));
  assign n584_1 = ~n8292;
  assign n8294 = (~Ng2879 & ~Ng2947) | (~Pg8023 & (Ng2879 | ~Ng2947));
  assign n576_1 = ~n8294;
  assign n8296 = (~Ng2879 & ~Ng2953) | (~Pg4321 & (Ng2879 | ~Ng2953));
  assign n568_1 = ~n8296;
  assign n8298 = (~Ng2879 & ~Ng2956) | (~Pg4088 & (Ng2879 | ~Ng2956));
  assign n560_1 = ~n8298;
  assign n8300 = (~Ng2879 & ~Ng2959) | (~Pg8249 & (Ng2879 | ~Ng2959));
  assign n552_1 = ~n8300;
  assign n8302 = (~Ng2879 & ~Ng2963) | (~Pg7334 & (Ng2879 | ~Ng2963));
  assign n536_1 = ~n8302;
  assign n8304 = (~Ng2879 & ~Ng2966) | (~Pg6895 & (Ng2879 | ~Ng2966));
  assign n528_1 = ~n8304;
  assign n8306 = (~Ng2879 & ~Ng2969) | (~Pg6442 & (Ng2879 | ~Ng2969));
  assign n520_1 = ~n8306;
  assign n8308 = (~Ng2879 & ~Ng2972) | (~Pg6225 & (Ng2879 | ~Ng2972));
  assign n512_1 = ~n8308;
  assign n8310 = (~Ng1315 & ~Ng3084) | (~Ng559 & (Ng1315 | ~Ng3084));
  assign n679_1 = ~n8310;
  assign n8312 = (~\[1603]  & ~Ng3211) | (~Ng559 & (\[1603]  | ~Ng3211));
  assign n674 = ~n8312;
  assign n8314 = (~\[1605]  & ~Ng3210) | (~Ng559 & (\[1605]  | ~Ng3210));
  assign n669_1 = ~n8314;
  assign n8316 = (~Ng1315 & ~Ng3088) | (~Ng8311 & (Ng1315 | ~Ng3088));
  assign n844_1 = ~n8316;
  assign n8318 = (~\[1603]  & ~Ng3185) | (~Ng8311 & (\[1603]  | ~Ng3185));
  assign n839_1 = ~n8318;
  assign n8320 = (~\[1605]  & ~Ng3182) | (~Ng8311 & (\[1605]  | ~Ng3182));
  assign n834_1 = ~n8320;
  assign n8322 = (~Ng1315 & ~Ng3179) | (~Ng8302 & (Ng1315 | ~Ng3179));
  assign n829_1 = ~n8322;
  assign n8324 = (~\[1603]  & ~Ng3176) | (~Ng8302 & (\[1603]  | ~Ng3176));
  assign n824_1 = ~n8324;
  assign n8326 = (~\[1605]  & ~Ng3173) | (~Ng8302 & (\[1605]  | ~Ng3173));
  assign n819_1 = ~n8326;
  assign n8328 = (~Ng1315 & ~Ng3170) | (~Ng8293 & (Ng1315 | ~Ng3170));
  assign n814_1 = ~n8328;
  assign n8330 = (~\[1603]  & ~Ng3167) | (~Ng8293 & (\[1603]  | ~Ng3167));
  assign n809_1 = ~n8330;
  assign n8332 = (~\[1605]  & ~Ng3164) | (~Ng8293 & (\[1605]  | ~Ng3164));
  assign n804_1 = ~n8332;
  assign n8334 = (~Ng1315 & ~Ng3161) | (~Ng8284 & (Ng1315 | ~Ng3161));
  assign n799_1 = ~n8334;
  assign n8336 = (~\[1603]  & ~Ng3158) | (~Ng8284 & (\[1603]  | ~Ng3158));
  assign n794_1 = ~n8336;
  assign n8338 = (~\[1605]  & ~Ng3155) | (~Ng8284 & (\[1605]  | ~Ng3155));
  assign n789_1 = ~n8338;
  assign n8340 = (~Ng1315 & ~Ng3096) | (~Ng2633 & (Ng1315 | ~Ng3096));
  assign n724_1 = ~n8340;
  assign n8342 = (~\[1603]  & ~Ng3095) | (~Ng2633 & (\[1603]  | ~Ng3095));
  assign n719_1 = ~n8342;
  assign n8344 = (~\[1605]  & ~Ng3094) | (~Ng2633 & (\[1605]  | ~Ng3094));
  assign n714_1 = ~n8344;
  assign n8346 = (~Ng1315 & ~Ng3093) | (~Ng1939 & (Ng1315 | ~Ng3093));
  assign n709_1 = ~n8346;
  assign n8348 = (~\[1603]  & ~Ng3092) | (~Ng1939 & (\[1603]  | ~Ng3092));
  assign n704_1 = ~n8348;
  assign n8350 = (~\[1605]  & ~Ng3091) | (~Ng1939 & (\[1605]  | ~Ng3091));
  assign n699_1 = ~n8350;
  assign n8352 = (~Ng1315 & ~Ng3087) | (~Ng1245 & (Ng1315 | ~Ng3087));
  assign n694 = ~n8352;
  assign n8354 = (~\[1603]  & ~Ng3086) | (~Ng1245 & (\[1603]  | ~Ng3086));
  assign n689_1 = ~n8354;
  assign n8356 = (~\[1605]  & ~Ng3085) | (~Ng1245 & (\[1605]  | ~Ng3085));
  assign n684_1 = ~n8356;
  assign n8358 = (Ng2987 & ~Ng3074) | (~Ng3056 & (~Ng2987 | ~Ng3074));
  assign n7230 = ~n8358;
  assign n8360 = (Ng2987 & ~Ng3073) | (~Ng3055 & (~Ng2987 | ~Ng3073));
  assign n7226 = ~n8360;
  assign n8362 = (Ng2987 & ~Ng3072) | (~Ng3053 & (~Ng2987 | ~Ng3072));
  assign n7222 = ~n8362;
  assign n8364 = (Ng2987 & ~Ng3071) | (~Ng3052 & (~Ng2987 | ~Ng3071));
  assign n7218 = ~n8364;
  assign n8366 = (Ng2987 & ~Ng3070) | (~Ng3051 & (~Ng2987 | ~Ng3070));
  assign n7204 = ~n8366;
  assign n8368 = (Ng2987 & ~Ng3069) | (~Ng3050 & (~Ng2987 | ~Ng3069));
  assign n7200 = ~n8368;
  assign n8370 = (Ng2987 & ~Ng3068) | (~Ng3049 & (~Ng2987 | ~Ng3068));
  assign n7196 = ~n8370;
  assign n8372 = (Ng2987 & ~Ng3067) | (~Ng3048 & (~Ng2987 | ~Ng3067));
  assign n7192 = ~n8372;
  assign n8374 = (Ng2987 & ~Ng3066) | (~Ng3047 & (~Ng2987 | ~Ng3066));
  assign n7188 = ~n8374;
  assign n8376 = (Ng2987 & ~Ng3065) | (~Ng3046 & (~Ng2987 | ~Ng3065));
  assign n7184 = ~n8376;
  assign n8378 = (Ng2987 & ~Ng3064) | (~Ng3045 & (~Ng2987 | ~Ng3064));
  assign n7180 = ~n8378;
  assign n8380 = (Ng2987 & ~Ng3063) | (~Ng3044 & (~Ng2987 | ~Ng3063));
  assign n7176 = ~n8380;
  assign n8382 = (Ng2987 & ~Ng3062) | (~Ng3043 & (~Ng2987 | ~Ng3062));
  assign n7172 = ~n8382;
  assign n8384 = (Ng2987 & ~Ng2997) | (~Ng3061 & (~Ng2987 | ~Ng2997));
  assign n7250 = ~n8384;
  assign n8386 = (Ng2987 & ~Ng3078) | (~Ng3060 & (~Ng2987 | ~Ng3078));
  assign n7246 = ~n8386;
  assign n8388 = (Ng2987 & ~Ng3077) | (~Ng3059 & (~Ng2987 | ~Ng3077));
  assign n7242 = ~n8388;
  assign n8390 = (Ng2987 & ~Ng3076) | (~Ng3058 & (~Ng2987 | ~Ng3076));
  assign n7238 = ~n8390;
  assign n8392 = (Ng2987 & ~Ng3075) | (~Ng3057 & (~Ng2987 | ~Ng3075));
  assign n7234 = ~n8392;
  assign n8394 = (Ng2879 & ~Ng2874) | (~Ng2200 & (~Ng2879 | ~Ng2874));
  assign n624_1 = ~n8394;
  assign n8396 = (Ng2879 & ~Ng2978) | (~Ng2190 & (~Ng2879 | ~Ng2978));
  assign n634_1 = ~n8396;
  assign n8398 = (Ng2879 & ~Ng2981) | (~Ng2195 & (~Ng2879 | ~Ng2981));
  assign n629_1 = ~n8398;
  assign n8400 = (Ng2879 & ~Ng2975) | (~Ng2185 & (~Ng2879 | ~Ng2975));
  assign n639_1 = ~n8400;
  assign n8402 = (Ng2879 & ~Ng2972) | (~Ng2180 & (~Ng2879 | ~Ng2972));
  assign n644_1 = ~n8402;
  assign n8404 = (Ng2879 & ~Ng2969) | (~Ng2175 & (~Ng2879 | ~Ng2969));
  assign n649_1 = ~n8404;
  assign n8406 = (Ng2879 & ~Ng2966) | (~Ng2170 & (~Ng2879 | ~Ng2966));
  assign n654_1 = ~n8406;
  assign n8408 = (Ng2879 & ~Ng2963) | (~Ng2165 & (~Ng2879 | ~Ng2963));
  assign n659_1 = ~n8408;
  assign n8410 = (Ng2879 & ~Ng2935) | (~Ng1471 & (~Ng2879 | ~Ng2935));
  assign n470_1 = ~n8410;
  assign n8412 = (Ng2879 & ~Ng2938) | (~Ng1476 & (~Ng2879 | ~Ng2938));
  assign n465 = ~n8412;
  assign n8414 = (Ng2879 & ~Ng2941) | (~Ng1481 & (~Ng2879 | ~Ng2941));
  assign n460_1 = ~n8414;
  assign n8416 = (Ng2879 & ~Ng2944) | (~Ng1486 & (~Ng2879 | ~Ng2944));
  assign n455_1 = ~n8416;
  assign n8418 = (Ng2879 & ~Ng2947) | (~Ng1491 & (~Ng2879 | ~Ng2947));
  assign n450_1 = ~n8418;
  assign n8420 = (Ng2879 & ~Ng2953) | (~Ng1496 & (~Ng2879 | ~Ng2953));
  assign n445_1 = ~n8420;
  assign n8422 = (Ng2879 & ~Ng2956) | (~Ng1501 & (~Ng2879 | ~Ng2956));
  assign n440_1 = ~n8422;
  assign n8424 = (Ng2879 & ~Ng2959) | (~Ng1506 & (~Ng2879 | ~Ng2959));
  assign n435_1 = ~n8424;
  assign n8426 = (~Ng1315 & ~Ng2704) | (~Ng2584 & (Ng1315 | ~Ng2704));
  assign n6642 = ~n8426;
  assign n8428 = (Ng1315 & ~Ng2631) | (~Ng2584 & (~Ng1315 | ~Ng2631));
  assign n6254 = ~n8428;
  assign n8430 = (Ng1315 & Ng2628) | (~Ng2631 & (~Ng1315 | Ng2628));
  assign n6249 = ~n8430;
  assign n8432 = (~Ng1315 & ~Ng2010) | (~Ng1890 & (Ng1315 | ~Ng2010));
  assign n5135 = ~n8432;
  assign n8434 = (Ng1315 & ~Ng1937) | (~Ng1890 & (~Ng1315 | ~Ng1937));
  assign n4747 = ~n8434;
  assign n8436 = (Ng1315 & Ng1934) | (~Ng1937 & (~Ng1315 | Ng1934));
  assign n4742 = ~n8436;
  assign n8438 = (~Ng1315 & ~Ng1316) | (~Ng1196 & (Ng1315 | ~Ng1316));
  assign n3641_1 = ~n8438;
  assign n8440 = (Ng1315 & ~Ng1243) | (~Ng1196 & (~Ng1315 | ~Ng1243));
  assign n3240_1 = ~n8440;
  assign n8442 = (Ng1315 & Ng1240) | (~Ng1243 & (~Ng1315 | Ng1240));
  assign n3235_1 = ~n8442;
  assign n8444 = (~Ng1315 & ~Ng630) | (~Ng510 & (Ng1315 | ~Ng630));
  assign n2122_1 = ~n8444;
  assign n8446 = (Ng1315 & ~Ng557) | (~Ng510 & (~Ng1315 | ~Ng557));
  assign n1734_1 = ~n8446;
  assign n8448 = (Ng1315 & Ng554) | (~Ng557 & (~Ng1315 | Ng554));
  assign n1729_1 = ~n8448;
  assign n8450 = n5054 | n5981;
  assign n8451 = n5058_1 | n5955;
  assign n8452 = ~n4978_1 & n5840;
  assign n8453 = n5062 | ~n5840;
  assign n8454 = ~n4982 & n5833_1;
  assign n8455 = n5064 | ~n5833_1;
  assign n8456 = (~Ng1315 | Ng2811) & (~\[1605]  | Ng2812);
  assign n8457 = n4948_1 & (~n8456 | (\[1603]  & ~Ng2813));
  assign n8458 = (Ng2611 | n6476) & (n5072_1 | n5577);
  assign n8459 = (n5072_1 | ~n5590_1) & (n6476 | Ng2610);
  assign n8460 = (n5072_1 | ~n5587) & (n6476 | Ng2608);
  assign n8461 = (n5072_1 | ~n5585_1) & (n6476 | Ng2607);
  assign n8462 = (n5072_1 | ~n5579) & (n6476 | Ng2606);
  assign n8463 = (n5072_1 | ~n5589) & (n6476 | Ng2605);
  assign n8464 = (n5072_1 | ~n5583) & (n6476 | Ng2604);
  assign n8465 = (n5072_1 | ~n5581) & (n6476 | Ng2603);
  assign n8466 = (~Ng1315 | Ng2117) & (~\[1605]  | Ng2118);
  assign n8467 = n4936 & (~n8466 | (\[1603]  & ~Ng2119));
  assign n8468 = (n5070 | ~n5573) & (n6478 | Ng1917);
  assign n8469 = (n5070 | ~n5571) & (n6478 | Ng1916);
  assign n8470 = (n5070 | ~n5568) & (n6478 | Ng1914);
  assign n8471 = (n5070 | ~n5566) & (n6478 | Ng1913);
  assign n8472 = (n5070 | ~n5560_1) & (n6478 | Ng1912);
  assign n8473 = (n5070 | ~n5570_1) & (n6478 | Ng1911);
  assign n8474 = (n5070 | ~n5564) & (n6478 | Ng1910);
  assign n8475 = (n5070 | ~n5562) & (n6478 | Ng1909);
  assign n8476 = (n6293 | n5853_1) & (n6294_1 | n6295);
  assign n8477 = (n6295 | n5853_1) & (n6293 | n6296);
  assign n8478 = (~n6296 | ~n8476) & (~n6294_1 | ~n8477);
  assign n8479 = (n5847 | n6297) & (~n6298 | n6299_1);
  assign n8480 = (n5847 | n6299_1) & (n6297 | n6300);
  assign n8481 = (~n6300 | ~n8479) & (n6298 | ~n8480);
  assign n8482 = (n6317_1 | n5873_1) & (n6318 | n6319);
  assign n8483 = (n6319 | n5873_1) & (n6317_1 | n6320);
  assign n8484 = (~n6320 | ~n8482) & (~n6318 | ~n8483);
  assign n8485 = (n5867 | n6321_1) & (~n6322 | n6323);
  assign n8486 = (n5867 | n6323) & (n6321_1 | n6324);
  assign n8487 = (~n6324 | ~n8485) & (n6322 | ~n8486);
  assign n8488 = (n6341_1 | n5893_1) & (n6342 | n6343);
  assign n8489 = (n6343 | n5893_1) & (n6341_1 | n6344);
  assign n8490 = (~n6344 | ~n8488) & (~n6342 | ~n8489);
  assign n8491 = (n5887 | n6345_1) & (~n6346 | n6347);
  assign n8492 = (n5887 | n6347) & (n6345_1 | n6348);
  assign n8493 = (~n6348 | ~n8491) & (n6346 | ~n8492);
  assign n8494 = (n6365 | n5913_1) & (n6366 | n6367);
  assign n8495 = (n6367 | n5913_1) & (n6365 | n6368_1);
  assign n8496 = (~n6368_1 | ~n8494) & (~n6366 | ~n8495);
  assign n8497 = (n5907 | n6369) & (~n6370 | n6371);
  assign n8498 = (n5907 | n6371) & (n6369 | n6372);
  assign n8499 = (~n6372 | ~n8497) & (n6370 | ~n8498);
  assign n8500 = (~Ng1315 | Ng1423) & (~\[1605]  | Ng1424);
  assign n8501 = n4932 | n4862 | n4798 | n4734 | n4712_1 | n4764;
  assign n8502 = (n5068 | ~n5538) & (n6520_1 | Ng1223);
  assign n8503 = (n5068 | ~n5536) & (n6520_1 | Ng1222);
  assign n8504 = (n5068 | ~n5533) & (n6520_1 | Ng1220);
  assign n8505 = (n5068 | ~n5531) & (n6520_1 | Ng1219);
  assign n8506 = (n5068 | ~n5540_1) & (n6520_1 | Ng1218);
  assign n8507 = (n5068 | ~n5535_1) & (n6520_1 | Ng1217);
  assign n8508 = (n5068 | ~n5529) & (n6520_1 | Ng1216);
  assign n8509 = (n5068 | ~n5526) & (n6520_1 | Ng1215);
  assign n8510 = (~Ng1315 | Ng737) & (~\[1605]  | Ng738);
  assign n8511 = n4912 | n4820 | n4756_1 | n4704_1 | n4688_1 | n4728_1;
  assign n8512 = (n5066 | ~n5518) & (n6526 | Ng537);
  assign n8513 = (n5066 | ~n5516) & (n6526 | Ng536);
  assign n8514 = (n5066 | ~n5513) & (n6526 | Ng534);
  assign n8515 = (n5066 | ~n5511) & (n6526 | Ng533);
  assign n8516 = (n5066 | ~n5520_1) & (n6526 | Ng532);
  assign n8517 = (n5066 | ~n5515_1) & (n6526 | Ng531);
  assign n8518 = (n5066 | ~n5509) & (n6526 | Ng530);
  assign n8519 = (n5066 | ~n5522) & (n6526 | Ng529);
  assign n8520 = n5028_1 | n4561 | n4571;
  assign n8521 = n8520 & (n6552 | n6057_1);
  assign n8522 = (~n5018_1 | n6051) & (~n4567 | n6552);
  assign n8523 = n5016 | n4553 | n4565;
  assign n8524 = n8523 & (n6557 | n6079);
  assign n8525 = (~n5006 | n6073) & (~n4559_1 | n6557);
  assign n8526 = n5004 | n4547 | n4557;
  assign n8527 = n8526 & (n6561 | n6101);
  assign n8528 = (~n4994 | n6095) & (~n4551 | n6561);
  assign n8529 = n4992 | n4543 | n4549;
  assign n8530 = n8529 & (n6565_1 | n6123);
  assign n8531 = (~n4986 | n6117) & (~n4545 | n6565_1);
  assign n8532 = n6531 | ~n8745;
  assign n8533 = (~Ng853 | Ng2253) & (~\[1612]  | Ng2254);
  assign n8534 = (~Ng853 | Ng1559) & (~\[1612]  | Ng1560);
  assign n8535 = (~Ng853 | Ng865) & (~\[1612]  | Ng866);
  assign n8536 = (~Ng853 | Ng177) & (~\[1612]  | Ng178);
  assign n8537 = n6437 | n6435_1 | n6436;
  assign n8538 = n6440_1 | n6441 | n6442 | n6443 | n6439 | n8537 | n6444 | n6438;
  assign n8539 = ~Ng1315 | Ng2802;
  assign n8540 = n6447 | n6445_1 | n6446;
  assign n8541 = n6450_1 | n6451 | n6452 | n6453 | n6449 | n8540 | n6454 | n6448;
  assign n8542 = ~Ng1315 | Ng2108;
  assign n8543 = n6457 | n6455_1 | n6456;
  assign n8544 = n6460_1 | n6461 | n6462 | n6463 | n6459 | n8543 | n6464 | n6458;
  assign n8545 = ~Ng1315 | Ng1414;
  assign n8546 = n6467 | n6465_1 | n6466;
  assign n8547 = n6470_1 | n6471 | n6472 | n6473 | n6469 | n8546 | n6474 | n6468;
  assign n8548 = ~Ng1315 | Ng728;
  assign n8549 = n6522 & (Ng3139 | ~n8756);
  assign n8550 = ~Ng548 | \[1605]  | Ng8284;
  assign n8551 = (~\[1605]  & ~Ng1234) | (n6600 & (\[1605]  | ~Ng1234));
  assign n8552 = (~\[1605]  & ~Ng1928) | (n6601 & (\[1605]  | ~Ng1928));
  assign n8553 = (~\[1605]  & ~Ng2622) | (n6602_1 & (\[1605]  | ~Ng2622));
  assign n8554 = (~n4776 & n8454) | (n4982 & (n4776 | n8454));
  assign n8555 = (~Pg3229 & Ng2615) | (Ng2612 & (Pg3229 | Ng2615));
  assign n8556 = n5649 ^ ~n5650_1;
  assign n8557 = ~n8555 | Ng2631 | n6476;
  assign n8558 = (~Pg3229 & Ng1921) | (Ng1918 & (Pg3229 | Ng1921));
  assign n8559 = n5637 ^ ~n5638;
  assign n8560 = ~n8558 | Ng1937 | n6478;
  assign n8561 = ~n4980 & (n6485_1 | (~n4643 & ~n5989));
  assign n8562 = n4976 & (n8561 | (n4980 & ~n6277));
  assign n8563 = ~n4976 & (n4970 | n5558);
  assign n8564 = n4976 & ~n5558 & (~n4970 | n4980);
  assign n8565 = ~n5445_1 | n8563 | n8564;
  assign n8566 = ~n4974 & (n6495_1 | (~n4639 & ~n5997));
  assign n8567 = n4968_1 & (n8566 | (n4974 & ~n6278));
  assign n8568 = ~n4968_1 & (n4962 | n5556);
  assign n8569 = n4968_1 & ~n5556 & (~n4962 | n4974);
  assign n8570 = ~n5442 | n8568 | n8569;
  assign n8571 = ~n4966 & (n6505_1 | (~n4633 & ~n6005));
  assign n8572 = n4960 & (n8571 | (n4966 & ~n6279));
  assign n8573 = ~n4960 & (n4956 | n5554);
  assign n8574 = n4960 & ~n5554 & (~n4956 | n4966);
  assign n8575 = ~n5439 | n8573 | n8574;
  assign n8576 = ~n4958_1 & (n6515_1 | (~n4625 & ~n6013_1));
  assign n8577 = n4954 & (n8576 | (n4958_1 & ~n6280));
  assign n8578 = ~n4954 & (n4950 | n5552);
  assign n8579 = n4954 & ~n5552 & (~n4950 | n4958_1);
  assign n8580 = ~n5436 | n8578 | n8579;
  assign n8581 = n4976 & (~n4980 | ~Ng2257 | n6483);
  assign n8582 = n4968_1 & (~n4974 | ~Ng2257 | n6493);
  assign n8583 = n4960 & (~n4966 | ~Ng2257 | n6503);
  assign n8584 = n4954 & (~n4958_1 | ~Ng2257 | n6513);
  assign n8585 = n4876_1 ^ ~n5928_1;
  assign n8586 = n4720_1 ^ ~n5927;
  assign n8587 = n4938_1 | n6488 | n6308_1;
  assign n8588 = n8587 & (~n4938_1 | (~n6308_1 & ~n6488));
  assign n8589 = n4834_1 ^ ~n5935;
  assign n8590 = n4696_1 ^ ~n5934;
  assign n8591 = n4918 | n6498 | n6332;
  assign n8592 = n8591 & (~n4918 | (~n6332 & ~n6498));
  assign n8593 = n4792_1 ^ ~n5942;
  assign n8594 = n4676_1 ^ ~n5941;
  assign n8595 = n4888_1 | n6508 | n6356;
  assign n8596 = n8595 & (~n4888_1 | (~n6356 & ~n6508));
  assign n8597 = n4750 ^ ~n5949;
  assign n8598 = n4662 ^ ~n5948_1;
  assign n8599 = n4850 | n6518 | n6380;
  assign n8600 = n8599 & (~n4850 | (~n6380 & ~n6518));
  assign n8601 = Ng506 | \[1603]  | Pg16297;
  assign n2064_1 = n8601 & (~Ng506 | Ng507);
  assign n8603 = (\[1603]  & n2064_1) | (Pg16355 & (~\[1603]  | n2064_1));
  assign n3570_1 = (Ng1192 & Ng1193) | (n8603 & (~Ng1192 | Ng1193));
  assign n8605 = (\[1603]  & n3570_1) | (Pg16399 & (~\[1603]  | n3570_1));
  assign n8606 = (\[1603]  & ~n5077) | (~Pg16437 & (~\[1603]  | ~n5077));
  assign n8607 = Ng298 | Ng299;
  assign n8608 = (~\[1594]  & ~Ng992) | (n6934 & (\[1594]  | ~Ng992));
  assign n8609 = (~\[1594]  & ~Ng1686) | (n6936_1 & (\[1594]  | ~Ng1686));
  assign n8610 = (~\[1594]  & ~Ng2380) | (n6938 & (\[1594]  | ~Ng2380));
  assign n8611 = (~Pg3229 & Ng1227) | (Ng1224 & (Pg3229 | Ng1227));
  assign n8612 = n5625_1 ^ ~n5626;
  assign n8613 = ~n8611 | Ng1243 | n6520_1;
  assign n8614 = ~n5445_1 | n5961;
  assign n8615 = ~n5442 | n5964;
  assign n8616 = ~n5439 | n5967;
  assign n8617 = ~n5436 | n5970;
  assign n8618 = (~Pg3229 & Ng541) | (Ng538 & (Pg3229 | Ng541));
  assign n8619 = n5613 ^ ~n5614;
  assign n8620 = ~n8618 | Ng557 | n6526;
  assign n8621 = n5034 ^ ~n5988_1;
  assign n8622 = (n5990 & n6484) | (Ng2257 & (~n5990 | n6484));
  assign n8623 = Ng853 & n8622;
  assign n8624 = \[1594]  & n8622;
  assign n8625 = \[1612]  & n8622;
  assign n8626 = n5022 ^ ~n5996;
  assign n8627 = (n5998_1 & n6494) | (Ng2257 & (~n5998_1 | n6494));
  assign n8628 = Ng853 & n8627;
  assign n8629 = \[1594]  & n8627;
  assign n8630 = \[1612]  & n8627;
  assign n8631 = n5010 ^ ~n6004;
  assign n8632 = (n6006 & n6504) | (Ng2257 & (~n6006 | n6504));
  assign n8633 = Ng853 & n8632;
  assign n8634 = \[1594]  & n8632;
  assign n8635 = \[1612]  & n8632;
  assign n8636 = n4998_1 ^ ~n6012;
  assign n8637 = (n6014 & n6514) | (Ng2257 & (~n6014 | n6514));
  assign n8638 = Ng853 & n8637;
  assign n8639 = \[1594]  & n8637;
  assign n8640 = \[1612]  & n8637;
  assign n8641 = n6020 | n5411;
  assign n8642 = ~n5026 ^ ~n8641;
  assign n8643 = n6024 | n5404;
  assign n8644 = ~n5014 ^ ~n8643;
  assign n8645 = n6028_1 | n5397;
  assign n8646 = ~n5002 ^ ~n8645;
  assign n8647 = n6032 | n5392;
  assign n8648 = ~n4990 ^ ~n8647;
  assign n8649 = n6555_1 | n4982;
  assign n8650 = n8649 & (n6554 | ~n6555_1 | ~n7062);
  assign n8651 = (n6555_1 & ~n7070) | (n5064 & (~n6555_1 | ~n7070));
  assign n8652 = n6555_1 | n4978_1;
  assign n8653 = n8652 & (~n6555_1 | n6559 | ~n7078);
  assign n8654 = (n6555_1 & ~n7086_1) | (n5062 & (~n6555_1 | ~n7086_1));
  assign n8655 = n6555_1 | n4972;
  assign n8656 = n8655 & (~n6555_1 | n6563 | ~n7094);
  assign n8657 = (n6555_1 & ~n7102) | (n5058_1 & (~n6555_1 | ~n7102));
  assign n8658 = n6555_1 | n4964;
  assign n8659 = n8658 & (~n6555_1 | n6567 | ~n7110);
  assign n8660 = (n6555_1 & ~n7118) | (n5054 & (~n6555_1 | ~n7118));
  assign n8661 = ~n4880_1 | n4908 | n6150;
  assign n8662 = ~n4838_1 | n4870 | n6157;
  assign n8663 = ~n4796_1 | n4828 | n6164;
  assign n8664 = ~n4754 | n4786 | n6171_1;
  assign n8665 = ~Ng1315 | n5156;
  assign n8666 = n6048_1 & n8669;
  assign n8667 = ~\[1603]  | n5156;
  assign n8668 = ~\[1605]  | n5156;
  assign n8669 = Pg3229 ^ ~n5008_1;
  assign n8670 = ~n5008_1 & n5036 & (n5018_1 | ~n5028_1);
  assign n8671 = Ng853 & n5138;
  assign n8672 = n4906 & n4926 & n6389;
  assign n8673 = \[1594]  & n5138;
  assign n8674 = \[1612]  & n5138;
  assign n8675 = ~n4878 & n4940 & (n4906 | ~n4926);
  assign n8676 = ~Ng1315 | n5149;
  assign n8677 = n6070 & n8680;
  assign n8678 = ~\[1603]  | n5149;
  assign n8679 = ~\[1605]  | n5149;
  assign n8680 = Pg3229 ^ ~n4996;
  assign n8681 = ~n4996 & n5024 & (n5006 | ~n5016);
  assign n8682 = Ng853 & n5136;
  assign n8683 = n4868 & n4896 & n6390;
  assign n8684 = \[1594]  & n5136;
  assign n8685 = \[1612]  & n5136;
  assign n8686 = ~n4836 & n4920 & (n4868 | ~n4896);
  assign n8687 = ~Ng1315 | n5147;
  assign n8688 = n6092 & n8691;
  assign n8689 = ~\[1603]  | n5147;
  assign n8690 = ~\[1605]  | n5147;
  assign n8691 = Pg3229 ^ ~n4988_1;
  assign n8692 = ~n4988_1 & n5012 & (n4994 | ~n5004);
  assign n8693 = Ng853 & n5132;
  assign n8694 = n4826 & n4858 & n6391_1;
  assign n8695 = \[1594]  & n5132;
  assign n8696 = \[1612]  & n5132;
  assign n8697 = ~n4794 & n4890 & (n4826 | ~n4858);
  assign n8698 = ~Ng1315 | n5142;
  assign n8699 = n6114 & n8702;
  assign n8700 = ~\[1603]  | n5142;
  assign n8701 = ~\[1605]  | n5142;
  assign n8702 = Pg3229 ^ ~n4984;
  assign n8703 = ~n4984 & n5000 & (n4986 | ~n4992);
  assign n8704 = Ng853 & n5128;
  assign n8705 = n4784 & n4816 & n6392;
  assign n8706 = \[1594]  & n5128;
  assign n8707 = \[1612]  & n5128;
  assign n8708 = ~n4752_1 & n4852 & (n4784 | ~n4816);
  assign n8709 = n4908 ^ ~n8755;
  assign n8710 = n4880_1 ^ ~n8757;
  assign n8711 = n4870 ^ ~n8754;
  assign n8712 = n4838_1 ^ ~n8758;
  assign n8713 = n4828 ^ ~n8753;
  assign n8714 = n4796_1 ^ ~n8759;
  assign n8715 = n4786 ^ ~n8752;
  assign n8716 = n4754 ^ ~n8760;
  assign n8717 = ~Ng2584 | ~n4581 | ~n4982;
  assign n8718 = ~Ng853 | ~Ng2257;
  assign n8719 = n4615 & ~n5989;
  assign n8720 = ~\[1594]  | ~Ng2257;
  assign n8721 = ~\[1612]  | ~Ng2257;
  assign n8722 = ~Ng1890 | ~n4579 | ~n4978_1;
  assign n8723 = n4603 & ~n5997;
  assign n8724 = ~Ng1196 | ~n4577_1 | ~n4972;
  assign n8725 = n4593 & ~n6005;
  assign n8726 = ~Ng510 | ~n4575 | ~n4964;
  assign n8727 = n4585 & ~n6013_1;
  assign n8728 = Ng13475 ^ ~Ng2993;
  assign n8729 = ~Ng853 | n6576;
  assign n8730 = ~\[1594]  | n6576;
  assign n8731 = ~\[1612]  | n6576;
  assign n8732 = ~Ng2185 | Ng2190 | Ng2195 | ~Ng2200;
  assign n8733 = ~Ng1491 | Ng1496 | Ng1501 | ~Ng1506;
  assign n8734 = ~Ng801 | Ng805 | Ng809 | ~Ng813;
  assign n8735 = ~Ng113 | Ng117 | Ng121 | ~Ng125;
  assign n8736 = n6555_1 | n6064;
  assign n8737 = n6555_1 | n5084;
  assign n8738 = n6242 & n5230_1;
  assign n8739 = n6555_1 | n6086;
  assign n8740 = n6555_1 | n5081;
  assign n8741 = n6555_1 | n6108;
  assign n8742 = n6555_1 | n5078;
  assign n8743 = n6555_1 | n6130;
  assign n8744 = n6555_1 | n5075;
  assign n8745 = Ng2985 | Ng2984;
  assign n8746 = ~Ng3147 & (~n8549 | (~Ng3120 & n8745));
  assign n8747 = ~\[1594]  | ~Ng2257;
  assign n8748 = ~\[1612]  | ~Ng2257;
  assign n8749 = n6595 ^ ~n8761;
  assign n8750 = Ng3006 | Ng3010 | Ng3024 | Ng3002 | Ng3013;
  assign n5815 = ~n6576;
  assign n8752 = n4583 | ~Ng2257 | n6571;
  assign n8753 = n4591_1 | ~Ng2257 | n6570_1;
  assign n8754 = n4601 | ~Ng2257 | n6569;
  assign n8755 = n4613_1 | ~Ng2257 | n6568;
  assign n8756 = Ng2991 | Ng2992;
  assign n8757 = ~Ng2257 | n6585;
  assign n8758 = ~Ng2257 | n6586;
  assign n8759 = ~Ng2257 | n6587_1;
  assign n8760 = ~Ng2257 | n6588;
  assign n8761 = Pg3231 | ~Ng3139;
  assign n8762 = Pg3231 | ~Ng3120;
  assign n8763 = ~n6597_1 ^ ~n8761;
  assign n8764 = ~n6389 & n4906 & n4940;
  assign n8765 = ~n6390 & n4868 & n4920;
  assign n8766 = ~n6391_1 & n4826 & n4890;
  assign n8767 = ~n6392 & n4784 & n4852;
  assign Pg25442 = n858_1;
  assign Pg25420 = n858_1;
  assign Pg8167 = \[1594] ;
  assign Pg8106 = \[1605] ;
  assign Pg8087 = \[1612] ;
  assign Pg8082 = \[1594] ;
  assign Pg8030 = \[1603] ;
  assign Pg8012 = \[1612] ;
  assign Pg8007 = \[1594] ;
  assign Pg7961 = \[1612] ;
  assign Pg7956 = \[1594] ;
  assign Pg7909 = \[1612] ;
  assign Pg7487 = \[1603] ;
  assign Pg7425 = \[1605] ;
  assign Pg7390 = \[1603] ;
  assign Pg7357 = \[1603] ;
  assign Pg7302 = \[1605] ;
  assign Pg7264 = \[1594] ;
  assign Pg7229 = \[1605] ;
  assign Pg7194 = \[1603] ;
  assign Pg7161 = \[1603] ;
  assign Pg7084 = \[1594] ;
  assign Pg7052 = \[1605] ;
  assign Pg7014 = \[1594] ;
  assign Pg6979 = \[1605] ;
  assign Pg6944 = \[1603] ;
  assign Pg6911 = \[1603] ;
  assign Pg6837 = \[1612] ;
  assign Pg6782 = \[1594] ;
  assign Pg6750 = \[1605] ;
  assign Pg6712 = \[1594] ;
  assign Pg6677 = \[1605] ;
  assign Pg6642 = \[1603] ;
  assign Pg6573 = \[1612] ;
  assign Pg6518 = \[1594] ;
  assign Pg6485 = \[1605] ;
  assign Pg6447 = \[1594] ;
  assign Pg6368 = \[1612] ;
  assign Pg6313 = \[1594] ;
  assign Pg6231 = \[1612] ;
  assign Pg5796 = \[1603] ;
  assign Pg5747 = \[1605] ;
  assign Pg5738 = \[1603] ;
  assign Pg5695 = \[1605] ;
  assign Pg5686 = \[1603] ;
  assign Pg5657 = \[1605] ;
  assign Pg5648 = \[1603] ;
  assign Pg5637 = \[1609] ;
  assign Pg5629 = \[1605] ;
  assign Pg5612 = \[1609] ;
  assign Pg5595 = \[1609] ;
  assign Pg5555 = \[1612] ;
  assign Pg5549 = \[1609] ;
  assign Pg5511 = \[1612] ;
  assign Pg5472 = \[1612] ;
  assign Pg5437 = \[1612] ;
  assign n270_1 = Pg51;
  assign n353_1 = Pg8021;
  assign n362_1 = Pg3212;
  assign n366_1 = Pg3228;
  assign n370_1 = Pg3227;
  assign n374_1 = Pg3226;
  assign n378_1 = Pg3225;
  assign n382_1 = Pg3224;
  assign n386 = Pg3223;
  assign n390_1 = Pg3222;
  assign n394 = Pg3221;
  assign n398_1 = Pg3232;
  assign n402_1 = Pg3220;
  assign n406 = Pg3219;
  assign n410_1 = Pg3218;
  assign n414_1 = Pg3217;
  assign n418_1 = Pg3216;
  assign n422_1 = Pg3215;
  assign n426_1 = Pg3214;
  assign n430_1 = Pg3213;
  assign n483_1 = Pg8251;
  assign n491_1 = Pg4090;
  assign n499_1 = Pg4323;
  assign n507 = Pg4590;
  assign n515_1 = Pg6225;
  assign n523_1 = Pg6442;
  assign n531_1 = Pg6895;
  assign n539_1 = Pg7334;
  assign n547_1 = Pg7519;
  assign n555_1 = Pg8249;
  assign n563_1 = Pg4088;
  assign n571_1 = Pg4321;
  assign n579 = Pg8023;
  assign n587_1 = Pg8175;
  assign n595_1 = Pg3993;
  assign n603_1 = Pg4200;
  assign n611_1 = Pg4450;
  assign n619_1 = Pg8096;
  assign n848_1 = Pg24734;
  assign n872_1 = Pg26104;
  assign n876_1 = Pg25435;
  assign n880_1 = Pg27380;
  assign n884_1 = Pg26149;
  assign n888_1 = Pg26135;
  assign n1537_1 = Ng450;
  assign n1546_1 = Ng452;
  assign n1555_1 = Ng454;
  assign n1564 = Ng280;
  assign n1573 = Ng282;
  assign n1582_1 = Ng284;
  assign n1591 = Ng286;
  assign n1600_1 = Ng288;
  assign n1604_1 = Ng13407;
  assign n1608 = Ng290;
  assign n1627_1 = Ng11497;
  assign n1631 = Ng342;
  assign n1635 = Ng11498;
  assign n1639_1 = Ng350;
  assign n1643 = Ng11499;
  assign n1647_1 = Ng352;
  assign n1651 = Ng11500;
  assign n1655 = Ng357;
  assign n1659_1 = Ng11501;
  assign n1663_1 = Ng365;
  assign n1667 = Ng11502;
  assign n1671_1 = Ng367;
  assign n1675_1 = Ng11503;
  assign n1679_1 = Ng372;
  assign n1683_1 = Ng11504;
  assign n1687_1 = Ng380;
  assign n1691_1 = Ng11505;
  assign n1695 = Ng382;
  assign n1699_1 = Ng11506;
  assign n1703 = Ng387;
  assign n1707 = Ng11507;
  assign n1711_1 = Ng395;
  assign n1715 = Ng11508;
  assign n1719 = Ng397;
  assign n1743 = Ng513;
  assign n1747 = Ng523;
  assign n1752_1 = Ng11512;
  assign n1756 = Ng564;
  assign n1761_1 = Ng11515;
  assign n1765 = Ng570;
  assign n1770_1 = Ng11516;
  assign n1774_1 = Ng572;
  assign n1779_1 = Ng11517;
  assign n1783_1 = Ng574;
  assign n1788 = Ng11513;
  assign n1792_1 = Ng566;
  assign n1797_1 = Ng11514;
  assign n1801_1 = Ng568;
  assign n1879_1 = Ng528;
  assign n1883_1 = Ng535;
  assign n1892 = Ng543;
  assign n1906_1 = Ng549;
  assign n1915_1 = Ng558;
  assign n2054_1 = Ng8284;
  assign n2067 = Pg16297;
  assign n2391 = Ng13457;
  assign n2395_1 = \[1612] ;
  assign n2399 = \[1594] ;
  assign n3043_1 = Ng1137;
  assign n3052_1 = Ng1139;
  assign n3061_1 = Ng1141;
  assign n3070 = Ng967;
  assign n3079_1 = Ng969;
  assign n3088_1 = Ng971;
  assign n3097_1 = Ng973;
  assign n3106_1 = Ng975;
  assign n3110_1 = Ng13423;
  assign n3114_1 = Ng977;
  assign n3133_1 = Ng11524;
  assign n3137_1 = Ng1029;
  assign n3141_1 = Ng11525;
  assign n3145_1 = Ng1037;
  assign n3149_1 = Ng11526;
  assign n3153_1 = Ng1039;
  assign n3157_1 = Ng11527;
  assign n3161_1 = Ng1044;
  assign n3165_1 = Ng11528;
  assign n3169_1 = Ng1052;
  assign n3173_1 = Ng11529;
  assign n3177_1 = Ng1054;
  assign n3181_1 = Ng11530;
  assign n3185_1 = Ng1059;
  assign n3189_1 = Ng11531;
  assign n3193_1 = Ng1067;
  assign n3197_1 = Ng11532;
  assign n3201_1 = Ng1069;
  assign n3205_1 = Ng11533;
  assign n3209_1 = Ng1074;
  assign n3213_1 = Ng11534;
  assign n3217_1 = Ng1082;
  assign n3221_1 = Ng11535;
  assign n3225_1 = Ng1084;
  assign n3249_1 = Ng1199;
  assign n3253_1 = Ng1209;
  assign n3258_1 = Ng11539;
  assign n3262_1 = Ng1250;
  assign n3267_1 = Ng11542;
  assign n3271_1 = Ng1256;
  assign n3276_1 = Ng11543;
  assign n3280_1 = Ng1258;
  assign n3285_1 = Ng11544;
  assign n3289_1 = Ng1260;
  assign n3294_1 = Ng11540;
  assign n3298_1 = Ng1252;
  assign n3303_1 = Ng11541;
  assign n3307_1 = Ng1254;
  assign n3385_1 = Ng1214;
  assign n3389_1 = Ng1221;
  assign n3398_1 = Ng1229;
  assign n3412_1 = Ng1235;
  assign n3421_1 = Ng1244;
  assign n3560_1 = Ng8293;
  assign n3573_1 = Pg16355;
  assign n3628_1 = Ng13475;
  assign n3632_1 = \[1605] ;
  assign n3636_1 = \[1603] ;
  assign n4550 = Ng1831;
  assign n4559 = Ng1833;
  assign n4568 = Ng1835;
  assign n4577 = Ng1661;
  assign n4586 = Ng1663;
  assign n4595 = Ng1665;
  assign n4604 = Ng1667;
  assign n4613 = Ng1669;
  assign n4617 = Ng13439;
  assign n4621 = Ng1671;
  assign n4640 = Ng11551;
  assign n4644_1 = Ng1723;
  assign n4648 = Ng11552;
  assign n4652 = Ng1731;
  assign n4656 = Ng11553;
  assign n4660 = Ng1733;
  assign n4664 = Ng11554;
  assign n4668 = Ng1738;
  assign n4672 = Ng11555;
  assign n4676 = Ng1746;
  assign n4680 = Ng11556;
  assign n4684 = Ng1748;
  assign n4688 = Ng11557;
  assign n4692 = Ng1753;
  assign n4696 = Ng11558;
  assign n4700 = Ng1761;
  assign n4704 = Ng11559;
  assign n4708 = Ng1763;
  assign n4712 = Ng11560;
  assign n4716 = Ng1768;
  assign n4720 = Ng11561;
  assign n4724 = Ng1776;
  assign n4728 = Ng11562;
  assign n4732 = Ng1778;
  assign n4756 = Ng1893;
  assign n4760 = Ng1903;
  assign n4765 = Ng11566;
  assign n4769 = Ng1944;
  assign n4774 = Ng11569;
  assign n4778 = Ng1950;
  assign n4783 = Ng11570;
  assign n4787 = Ng1952;
  assign n4792 = Ng11571;
  assign n4796 = Ng1954;
  assign n4801 = Ng11567;
  assign n4805 = Ng1946;
  assign n4810 = Ng11568;
  assign n4814 = Ng1948;
  assign n4892 = Ng1908;
  assign n4896_1 = Ng1915;
  assign n4905_1 = Ng1923;
  assign n4919 = Ng1929;
  assign n4928 = Ng1938;
  assign n5067 = Ng8302;
  assign n5080 = Pg16399;
  assign n5819 = Ng2256;
  assign n5823 = \[1609] ;
  assign n6057 = Ng2525;
  assign n6066 = Ng2527;
  assign n6075 = Ng2529;
  assign n6084 = Ng2355;
  assign n6093 = Ng2357;
  assign n6102 = Ng2359;
  assign n6111 = Ng2361;
  assign n6120 = Ng2363;
  assign n6124 = Ng13455;
  assign n6128 = Ng2365;
  assign n6147 = Ng11578;
  assign n6151 = Ng2417;
  assign n6155 = Ng11579;
  assign n6159 = Ng2425;
  assign n6163 = Ng11580;
  assign n6167 = Ng2427;
  assign n6171 = Ng11581;
  assign n6175 = Ng2432;
  assign n6179 = Ng11582;
  assign n6183 = Ng2440;
  assign n6187 = Ng11583;
  assign n6191 = Ng2442;
  assign n6195 = Ng11584;
  assign n6199 = Ng2447;
  assign n6203 = Ng11585;
  assign n6207 = Ng2455;
  assign n6211 = Ng11586;
  assign n6215 = Ng2457;
  assign n6219 = Ng11587;
  assign n6223 = Ng2462;
  assign n6227 = Ng11588;
  assign n6231 = Ng2470;
  assign n6235 = Ng11589;
  assign n6239 = Ng2472;
  assign n6263 = Ng2587;
  assign n6267 = Ng2597;
  assign n6272 = Ng11593;
  assign n6276 = Ng2638;
  assign n6281 = Ng11596;
  assign n6285 = Ng2644;
  assign n6290 = Ng11597;
  assign n6294 = Ng2646;
  assign n6299 = Ng11598;
  assign n6303 = Ng2648;
  assign n6308 = Ng11594;
  assign n6312 = Ng2640;
  assign n6317 = Ng11595;
  assign n6321 = Ng2642;
  assign n6399 = Ng2602;
  assign n6403 = Ng2609;
  assign n6412 = Ng2617;
  assign n6426 = Ng2623;
  assign n6435 = Ng2632;
  assign n6574 = Ng8311;
  assign n6587 = Pg16437;
  assign n7160 = Pg3234;
  assign n7163 = Pg5388;
  assign n7167 = Pg16496;
  always @ (posedge clock) begin
    Pg8021 <= n270_1;
    Ng2817 <= n274_1;
    Ng2933 <= n279_1;
    Ng13457 <= n284_1;
    Ng2883 <= n289_1;
    Ng2888 <= n294_1;
    Ng2896 <= n299_1;
    Ng2892 <= n304_1;
    Ng2903 <= n309_1;
    Ng2900 <= n314_1;
    Ng2908 <= n319_1;
    Ng2912 <= n324_1;
    Ng2917 <= n329;
    Ng2924 <= n334_1;
    Ng2920 <= n339;
    Ng2984 <= n344;
    Ng2985 <= n349_1;
    Ng2929 <= n353_1;
    Ng2879 <= n358_1;
    Ng2934 <= n362_1;
    Ng2935 <= n366_1;
    Ng2938 <= n370_1;
    Ng2941 <= n374_1;
    Ng2944 <= n378_1;
    Ng2947 <= n382_1;
    Ng2953 <= n386;
    Ng2956 <= n390_1;
    Ng2959 <= n394;
    Ng2962 <= n398_1;
    Ng2963 <= n402_1;
    Ng2966 <= n406;
    Ng2969 <= n410_1;
    Ng2972 <= n414_1;
    Ng2975 <= n418_1;
    Ng2978 <= n422_1;
    Ng2981 <= n426_1;
    Ng2874 <= n430_1;
    Ng1506 <= n435_1;
    Ng1501 <= n440_1;
    Ng1496 <= n445_1;
    Ng1491 <= n450_1;
    Ng1486 <= n455_1;
    Ng1481 <= n460_1;
    Ng1476 <= n465;
    Ng1471 <= n470_1;
    Ng13439 <= n475_1;
    Pg8251 <= n480_1;
    Ng813 <= n483_1;
    Pg4090 <= n488_1;
    Ng809 <= n491_1;
    Pg4323 <= n496_1;
    Ng805 <= n499_1;
    Pg4590 <= n504_1;
    Ng801 <= n507;
    Pg6225 <= n512_1;
    Ng797 <= n515_1;
    Pg6442 <= n520_1;
    Ng793 <= n523_1;
    Pg6895 <= n528_1;
    Ng789 <= n531_1;
    Pg7334 <= n536_1;
    Ng785 <= n539_1;
    Pg7519 <= n544_1;
    Ng13423 <= n547_1;
    Pg8249 <= n552_1;
    Ng125 <= n555_1;
    Pg4088 <= n560_1;
    Ng121 <= n563_1;
    Pg4321 <= n568_1;
    Ng117 <= n571_1;
    Pg8023 <= n576_1;
    Ng113 <= n579;
    Pg8175 <= n584_1;
    Ng109 <= n587_1;
    Pg3993 <= n592_1;
    Ng105 <= n595_1;
    Pg4200 <= n600_1;
    Ng101 <= n603_1;
    Pg4450 <= n608_1;
    Ng97 <= n611_1;
    Pg8096 <= n616;
    Ng13407 <= n619_1;
    Ng2200 <= n624_1;
    Ng2195 <= n629_1;
    Ng2190 <= n634_1;
    Ng2185 <= n639_1;
    Ng2180 <= n644_1;
    Ng2175 <= n649_1;
    Ng2170 <= n654_1;
    Ng2165 <= n659_1;
    Ng13455 <= n664_1;
    Ng3210 <= n669_1;
    Ng3211 <= n674;
    Ng3084 <= n679_1;
    Ng3085 <= n684_1;
    Ng3086 <= n689_1;
    Ng3087 <= n694;
    Ng3091 <= n699_1;
    Ng3092 <= n704_1;
    Ng3093 <= n709_1;
    Ng3094 <= n714_1;
    Ng3095 <= n719_1;
    Ng3096 <= n724_1;
    Ng3097 <= n729;
    Ng3098 <= n734_1;
    Ng3099 <= n739_1;
    Ng3100 <= n744_1;
    Ng3101 <= n749_1;
    Ng3102 <= n754_1;
    Ng3103 <= n759_1;
    Ng3104 <= n764_1;
    Ng3105 <= n769_1;
    Ng3106 <= n774;
    Ng3107 <= n779;
    Ng3108 <= n784_1;
    Ng3155 <= n789_1;
    Ng3158 <= n794_1;
    Ng3161 <= n799_1;
    Ng3164 <= n804_1;
    Ng3167 <= n809_1;
    Ng3170 <= n814_1;
    Ng3173 <= n819_1;
    Ng3176 <= n824_1;
    Ng3179 <= n829_1;
    Ng3182 <= n834_1;
    Ng3185 <= n839_1;
    Ng3088 <= n844_1;
    Ng3191 <= n848_1;
    Ng3128 <= n853_1;
    Ng3126 <= n858_1;
    Ng3125 <= n863_1;
    Ng3123 <= n868_1;
    Ng3120 <= n872_1;
    Ng3110 <= n876_1;
    Ng3139 <= n880_1;
    Ng3135 <= n884_1;
    Ng3147 <= n888_1;
    Ng185 <= n893_1;
    Ng130 <= n898_1;
    Ng131 <= n903_1;
    Ng129 <= n908_1;
    Ng133 <= n913_1;
    Ng134 <= n918_1;
    Ng132 <= n923_1;
    Ng142 <= n928;
    Ng143 <= n933_1;
    Ng141 <= n938_1;
    Ng145 <= n943_1;
    Ng146 <= n948_1;
    Ng144 <= n953_1;
    Ng148 <= n958;
    Ng149 <= n963_1;
    Ng147 <= n968_1;
    Ng151 <= n973_1;
    Ng152 <= n978_1;
    Ng150 <= n983_1;
    Ng154 <= n988_1;
    Ng155 <= n993_1;
    Ng153 <= n998;
    Ng157 <= n1003;
    Ng158 <= n1008_1;
    Ng156 <= n1013_1;
    Ng160 <= n1018;
    Ng161 <= n1023_1;
    Ng159 <= n1028_1;
    Ng163 <= n1033;
    Ng164 <= n1038_1;
    Ng162 <= n1043_1;
    Ng169 <= n1048;
    Ng170 <= n1053;
    Ng168 <= n1058_1;
    Ng172 <= n1063;
    Ng173 <= n1068_1;
    Ng171 <= n1073_1;
    Ng175 <= n1078_1;
    Ng176 <= n1083_1;
    Ng174 <= n1088_1;
    Ng178 <= n1093_1;
    Ng179 <= n1098_1;
    Ng177 <= n1103_1;
    Ng186 <= n1108;
    Ng189 <= n1113_1;
    Ng192 <= n1118_1;
    Ng231 <= n1123_1;
    Ng234 <= n1128_1;
    Ng237 <= n1133_1;
    Ng195 <= n1138_1;
    Ng198 <= n1143_1;
    Ng201 <= n1148_1;
    Ng240 <= n1153_1;
    Ng243 <= n1158_1;
    Ng246 <= n1163_1;
    Ng204 <= n1168_1;
    Ng207 <= n1173_1;
    Ng210 <= n1178;
    Ng249 <= n1183_1;
    Ng252 <= n1188_1;
    Ng255 <= n1193_1;
    Ng213 <= n1198_1;
    Ng216 <= n1203_1;
    Ng219 <= n1208_1;
    Ng258 <= n1213_1;
    Ng261 <= n1218_1;
    Ng264 <= n1223_1;
    Ng222 <= n1228_1;
    Ng225 <= n1233_1;
    Ng228 <= n1238_1;
    Ng267 <= n1243_1;
    Ng270 <= n1248_1;
    Ng273 <= n1253_1;
    Ng92 <= n1258_1;
    Ng88 <= n1263_1;
    Ng83 <= n1268;
    Ng79 <= n1273_1;
    Ng74 <= n1278;
    Ng70 <= n1283_1;
    Ng65 <= n1288;
    Ng61 <= n1293_1;
    Ng56 <= n1298;
    Ng52 <= n1303;
    Ng11497 <= n1308_1;
    Ng11498 <= n1313;
    Ng11499 <= n1318;
    Ng11500 <= n1323_1;
    Ng11501 <= n1328_1;
    Ng11502 <= n1333_1;
    Ng11503 <= n1338_1;
    Ng11504 <= n1343_1;
    Ng11505 <= n1348;
    Ng11506 <= n1353;
    Ng11507 <= n1358_1;
    Ng11508 <= n1363_1;
    Ng408 <= n1368;
    Ng411 <= n1373_1;
    Ng414 <= n1378_1;
    Ng417 <= n1383;
    Ng420 <= n1388;
    Ng423 <= n1393;
    Ng427 <= n1398_1;
    Ng428 <= n1403;
    Ng426 <= n1408_1;
    Ng429 <= n1413;
    Ng432 <= n1418_1;
    Ng435 <= n1423_1;
    Ng438 <= n1428_1;
    Ng441 <= n1433_1;
    Ng444 <= n1438_1;
    Ng448 <= n1443_1;
    Ng449 <= n1448_1;
    Ng447 <= n1453;
    Ng312 <= n1458_1;
    Ng313 <= n1463_1;
    Ng314 <= n1468_1;
    Ng315 <= n1473_1;
    Ng316 <= n1478_1;
    Ng317 <= n1483_1;
    Ng318 <= n1488_1;
    Ng319 <= n1493;
    Ng320 <= n1498;
    Ng322 <= n1503;
    Ng323 <= n1508;
    Ng321 <= n1513_1;
    Ng403 <= n1518_1;
    Ng404 <= n1523_1;
    Ng402 <= n1528;
    Ng450 <= n1533_1;
    Ng451 <= n1537_1;
    Ng452 <= n1542_1;
    Ng453 <= n1546_1;
    Ng454 <= n1551_1;
    Ng279 <= n1555_1;
    Ng280 <= n1560_1;
    Ng281 <= n1564;
    Ng282 <= n1569_1;
    Ng283 <= n1573;
    Ng284 <= n1578;
    Ng285 <= n1582_1;
    Ng286 <= n1587;
    Ng287 <= n1591;
    Ng288 <= n1596;
    Ng289 <= n1600_1;
    Ng290 <= n1604_1;
    Ng291 <= n1608;
    Ng299 <= n1613;
    Ng305 <= n1618_1;
    Ng298 <= n1623_1;
    Ng342 <= n1627_1;
    Ng349 <= n1631;
    Ng350 <= n1635;
    Ng351 <= n1639_1;
    Ng352 <= n1643;
    Ng353 <= n1647_1;
    Ng357 <= n1651;
    Ng364 <= n1655;
    Ng365 <= n1659_1;
    Ng366 <= n1663_1;
    Ng367 <= n1667;
    Ng368 <= n1671_1;
    Ng372 <= n1675_1;
    Ng379 <= n1679_1;
    Ng380 <= n1683_1;
    Ng381 <= n1687_1;
    Ng382 <= n1691_1;
    Ng383 <= n1695;
    Ng387 <= n1699_1;
    Ng394 <= n1703;
    Ng395 <= n1707;
    Ng396 <= n1711_1;
    Ng397 <= n1715;
    Ng324 <= n1719;
    Ng554 <= n1724_1;
    Ng557 <= n1729_1;
    Ng510 <= n1734_1;
    Ng513 <= n1739_1;
    Ng523 <= n1743;
    Ng524 <= n1747;
    Ng564 <= n1752_1;
    Ng569 <= n1756;
    Ng570 <= n1761_1;
    Ng571 <= n1765;
    Ng572 <= n1770_1;
    Ng573 <= n1774_1;
    Ng574 <= n1779_1;
    Ng565 <= n1783_1;
    Ng566 <= n1788;
    Ng567 <= n1792_1;
    Ng568 <= n1797_1;
    Ng489 <= n1801_1;
    Ng486 <= n1806_1;
    Ng487 <= n1811_1;
    Ng488 <= n1816_1;
    Ng11512 <= n1821_1;
    Ng11515 <= n1825_1;
    Ng11516 <= n1829;
    Ng477 <= n1833;
    Ng478 <= n1838;
    Ng479 <= n1843_1;
    Ng480 <= n1848;
    Ng484 <= n1853_1;
    Ng464 <= n1858_1;
    Ng11517 <= n1863;
    Ng11513 <= n1867_1;
    Ng11514 <= n1871_1;
    Ng528 <= n1875_1;
    Ng535 <= n1879_1;
    Ng542 <= n1883_1;
    Ng543 <= n1888;
    Ng544 <= n1892;
    Ng548 <= n1897_1;
    Ng549 <= n1902_1;
    Ng8284 <= n1906_1;
    Ng558 <= n1911_1;
    Ng559 <= n1915_1;
    Ng576 <= n1920_1;
    Ng577 <= n1925;
    Ng575 <= n1930_1;
    Ng579 <= n1935_1;
    Ng580 <= n1940_1;
    Ng578 <= n1945_1;
    Ng582 <= n1950;
    Ng583 <= n1955;
    Ng581 <= n1960_1;
    Ng585 <= n1965;
    Ng586 <= n1970_1;
    Ng584 <= n1975;
    Ng587 <= n1980;
    Ng590 <= n1985;
    Ng593 <= n1990_1;
    Ng596 <= n1995_1;
    Ng599 <= n2000_1;
    Ng602 <= n2005_1;
    Ng614 <= n2010;
    Ng617 <= n2015_1;
    Ng620 <= n2020_1;
    Ng605 <= n2025_1;
    Ng608 <= n2030;
    Ng611 <= n2035_1;
    Ng490 <= n2040;
    Ng493 <= n2045_1;
    Ng496 <= n2050_1;
    Ng506 <= n2054_1;
    Ng507 <= n2059_1;
    Pg16297 <= n2064_1;
    Ng525 <= n2067;
    Ng529 <= n2072_1;
    Ng530 <= n2077_1;
    Ng531 <= n2082;
    Ng532 <= n2087_1;
    Ng533 <= n2092_1;
    Ng534 <= n2097_1;
    Ng536 <= n2102_1;
    Ng537 <= n2107_1;
    Ng538 <= n2112;
    Ng541 <= n2117_1;
    Ng630 <= n2122_1;
    Ng659 <= n2127_1;
    Ng640 <= n2132;
    Ng633 <= n2137;
    Ng653 <= n2142_1;
    Ng646 <= n2147_1;
    Ng660 <= n2152_1;
    Ng672 <= n2157_1;
    Ng666 <= n2162_1;
    Ng679 <= n2167_1;
    Ng686 <= n2172_1;
    Ng692 <= n2177;
    Ng699 <= n2182_1;
    Ng700 <= n2187_1;
    Ng698 <= n2192_1;
    Ng702 <= n2197;
    Ng703 <= n2202;
    Ng701 <= n2207_1;
    Ng705 <= n2212_1;
    Ng706 <= n2217_1;
    Ng704 <= n2222;
    Ng708 <= n2227_1;
    Ng709 <= n2232;
    Ng707 <= n2237_1;
    Ng711 <= n2242;
    Ng712 <= n2247_1;
    Ng710 <= n2252;
    Ng714 <= n2257_1;
    Ng715 <= n2262;
    Ng713 <= n2267;
    Ng717 <= n2272;
    Ng718 <= n2277;
    Ng716 <= n2282;
    Ng720 <= n2287;
    Ng721 <= n2292;
    Ng719 <= n2297_1;
    Ng723 <= n2302;
    Ng724 <= n2307;
    Ng722 <= n2312;
    Ng726 <= n2317;
    Ng727 <= n2322;
    Ng725 <= n2327_1;
    Ng729 <= n2332_1;
    Ng730 <= n2337;
    Ng728 <= n2342;
    Ng732 <= n2347;
    Ng733 <= n2352;
    Ng731 <= n2357;
    Ng735 <= n2362_1;
    Ng736 <= n2367_1;
    Ng734 <= n2372;
    Ng738 <= n2377;
    Ng739 <= n2382;
    Ng737 <= n2387;
    \[1612]  <= n2391;
    \[1594]  <= n2395_1;
    Ng853 <= n2399;
    Ng818 <= n2404;
    Ng819 <= n2409;
    Ng817 <= n2414;
    Ng821 <= n2419;
    Ng822 <= n2424_1;
    Ng820 <= n2429_1;
    Ng830 <= n2434;
    Ng831 <= n2439;
    Ng829 <= n2444_1;
    Ng833 <= n2449;
    Ng834 <= n2454;
    Ng832 <= n2459;
    Ng836 <= n2464;
    Ng837 <= n2469;
    Ng835 <= n2474;
    Ng839 <= n2479;
    Ng840 <= n2484;
    Ng838 <= n2489_1;
    Ng842 <= n2494;
    Ng843 <= n2499_1;
    Ng841 <= n2504_1;
    Ng845 <= n2509;
    Ng846 <= n2514_1;
    Ng844 <= n2519_1;
    Ng848 <= n2524_1;
    Ng849 <= n2529;
    Ng847 <= n2534_1;
    Ng851 <= n2539;
    Ng852 <= n2544;
    Ng850 <= n2549;
    Ng857 <= n2554;
    Ng858 <= n2559;
    Ng856 <= n2564;
    Ng860 <= n2569;
    Ng861 <= n2574;
    Ng859 <= n2579;
    Ng863 <= n2584_1;
    Ng864 <= n2589;
    Ng862 <= n2594;
    Ng866 <= n2599_1;
    Ng867 <= n2604;
    Ng865 <= n2609;
    Ng873 <= n2614;
    Ng876 <= n2619_1;
    Ng879 <= n2624;
    Ng918 <= n2629;
    Ng921 <= n2634;
    Ng924 <= n2639;
    Ng882 <= n2644;
    Ng885 <= n2649;
    Ng888 <= n2654;
    Ng927 <= n2659;
    Ng930 <= n2664;
    Ng933 <= n2669;
    Ng891 <= n2674;
    Ng894 <= n2679;
    Ng897 <= n2684;
    Ng936 <= n2689;
    Ng939 <= n2694_1;
    Ng942 <= n2699_1;
    Ng900 <= n2704_1;
    Ng903 <= n2709;
    Ng906 <= n2714_1;
    Ng945 <= n2719;
    Ng948 <= n2724_1;
    Ng951 <= n2729_1;
    Ng909 <= n2734_1;
    Ng912 <= n2739_1;
    Ng915 <= n2744_1;
    Ng954 <= n2749_1;
    Ng957 <= n2754_1;
    Ng960 <= n2759_1;
    Ng780 <= n2764_1;
    Ng776 <= n2769_1;
    Ng771 <= n2774_1;
    Ng767 <= n2779_1;
    Ng762 <= n2784_1;
    Ng758 <= n2789_1;
    Ng753 <= n2794_1;
    Ng749 <= n2799_1;
    Ng744 <= n2804_1;
    Ng740 <= n2809_1;
    Ng11524 <= n2814_1;
    Ng11525 <= n2819_1;
    Ng11526 <= n2824_1;
    Ng11527 <= n2829_1;
    Ng11528 <= n2834_1;
    Ng11529 <= n2839_1;
    Ng11530 <= n2844_1;
    Ng11531 <= n2849_1;
    Ng11532 <= n2854_1;
    Ng11533 <= n2859_1;
    Ng11534 <= n2864_1;
    Ng11535 <= n2869_1;
    Ng1095 <= n2874_1;
    Ng1098 <= n2879_1;
    Ng1101 <= n2884_1;
    Ng1104 <= n2889;
    Ng1107 <= n2894;
    Ng1110 <= n2899;
    Ng1114 <= n2904;
    Ng1115 <= n2909_1;
    Ng1113 <= n2914_1;
    Ng1116 <= n2919_1;
    Ng1119 <= n2924_1;
    Ng1122 <= n2929_1;
    Ng1125 <= n2934_1;
    Ng1128 <= n2939_1;
    Ng1131 <= n2944_1;
    Ng1135 <= n2949_1;
    Ng1136 <= n2954_1;
    Ng1134 <= n2959_1;
    Ng999 <= n2964_1;
    Ng1000 <= n2969_1;
    Ng1001 <= n2974_1;
    Ng1002 <= n2979_1;
    Ng1003 <= n2984_1;
    Ng1004 <= n2989_1;
    Ng1005 <= n2994_1;
    Ng1006 <= n2999;
    Ng1007 <= n3004_1;
    Ng1009 <= n3009_1;
    Ng1010 <= n3014;
    Ng1008 <= n3019_1;
    Ng1090 <= n3024_1;
    Ng1091 <= n3029_1;
    Ng1089 <= n3034_1;
    Ng1137 <= n3039_1;
    Ng1138 <= n3043_1;
    Ng1139 <= n3048_1;
    Ng1140 <= n3052_1;
    Ng1141 <= n3057_1;
    Ng966 <= n3061_1;
    Ng967 <= n3066_1;
    Ng968 <= n3070;
    Ng969 <= n3075;
    Ng970 <= n3079_1;
    Ng971 <= n3084_1;
    Ng972 <= n3088_1;
    Ng973 <= n3093_1;
    Ng974 <= n3097_1;
    Ng975 <= n3102;
    Ng976 <= n3106_1;
    Ng977 <= n3110_1;
    Ng978 <= n3114_1;
    Ng986 <= n3119_1;
    Ng992 <= n3124_1;
    Ng985 <= n3129_1;
    Ng1029 <= n3133_1;
    Ng1036 <= n3137_1;
    Ng1037 <= n3141_1;
    Ng1038 <= n3145_1;
    Ng1039 <= n3149_1;
    Ng1040 <= n3153_1;
    Ng1044 <= n3157_1;
    Ng1051 <= n3161_1;
    Ng1052 <= n3165_1;
    Ng1053 <= n3169_1;
    Ng1054 <= n3173_1;
    Ng1055 <= n3177_1;
    Ng1059 <= n3181_1;
    Ng1066 <= n3185_1;
    Ng1067 <= n3189_1;
    Ng1068 <= n3193_1;
    Ng1069 <= n3197_1;
    Ng1070 <= n3201_1;
    Ng1074 <= n3205_1;
    Ng1081 <= n3209_1;
    Ng1082 <= n3213_1;
    Ng1083 <= n3217_1;
    Ng1084 <= n3221_1;
    Ng1011 <= n3225_1;
    Ng1240 <= n3230_1;
    Ng1243 <= n3235_1;
    Ng1196 <= n3240_1;
    Ng1199 <= n3245_1;
    Ng1209 <= n3249_1;
    Ng1210 <= n3253_1;
    Ng1250 <= n3258_1;
    Ng1255 <= n3262_1;
    Ng1256 <= n3267_1;
    Ng1257 <= n3271_1;
    Ng1258 <= n3276_1;
    Ng1259 <= n3280_1;
    Ng1260 <= n3285_1;
    Ng1251 <= n3289_1;
    Ng1252 <= n3294_1;
    Ng1253 <= n3298_1;
    Ng1254 <= n3303_1;
    Ng1176 <= n3307_1;
    Ng1173 <= n3312_1;
    Ng1174 <= n3317_1;
    Ng1175 <= n3322_1;
    Ng11539 <= n3327_1;
    Ng11542 <= n3331_1;
    Ng11543 <= n3335_1;
    Ng1164 <= n3339_1;
    Ng1165 <= n3344_1;
    Ng1166 <= n3349_1;
    Ng1167 <= n3354_1;
    Ng1171 <= n3359_1;
    Ng1151 <= n3364_1;
    Ng11544 <= n3369_1;
    Ng11540 <= n3373_1;
    Ng11541 <= n3377_1;
    Ng1214 <= n3381_1;
    Ng1221 <= n3385_1;
    Ng1228 <= n3389_1;
    Ng1229 <= n3394_1;
    Ng1230 <= n3398_1;
    Ng1234 <= n3403_1;
    Ng1235 <= n3408_1;
    Ng8293 <= n3412_1;
    Ng1244 <= n3417_1;
    Ng1245 <= n3421_1;
    Ng1262 <= n3426_1;
    Ng1263 <= n3431_1;
    Ng1261 <= n3436_1;
    Ng1265 <= n3441_1;
    Ng1266 <= n3446_1;
    Ng1264 <= n3451_1;
    Ng1268 <= n3456_1;
    Ng1269 <= n3461_1;
    Ng1267 <= n3466_1;
    Ng1271 <= n3471_1;
    Ng1272 <= n3476_1;
    Ng1270 <= n3481_1;
    Ng1273 <= n3486_1;
    Ng1276 <= n3491_1;
    Ng1279 <= n3496_1;
    Ng1282 <= n3501_1;
    Ng1285 <= n3506_1;
    Ng1288 <= n3511_1;
    Ng1300 <= n3516_1;
    Ng1303 <= n3521_1;
    Ng1306 <= n3526_1;
    Ng1291 <= n3531_1;
    Ng1294 <= n3536_1;
    Ng1297 <= n3541_1;
    Ng1177 <= n3546_1;
    Ng1180 <= n3551_1;
    Ng1183 <= n3556_1;
    Ng1192 <= n3560_1;
    Ng1193 <= n3565_1;
    Pg16355 <= n3570_1;
    Ng1211 <= n3573_1;
    Ng1215 <= n3578_1;
    Ng1216 <= n3583_1;
    Ng1217 <= n3588_1;
    Ng1218 <= n3593_1;
    Ng1219 <= n3598_1;
    Ng1220 <= n3603_1;
    Ng1222 <= n3608_1;
    Ng1223 <= n3613_1;
    Ng1224 <= n3618_1;
    Ng1227 <= n3623_1;
    \[1605]  <= n3628_1;
    \[1603]  <= n3632_1;
    Ng1315 <= n3636_1;
    Ng1316 <= n3641_1;
    Ng1345 <= n3646_1;
    Ng1326 <= n3651_1;
    Ng1319 <= n3656_1;
    Ng1339 <= n3661_1;
    Ng1332 <= n3666_1;
    Ng1346 <= n3671_1;
    Ng1358 <= n3676_1;
    Ng1352 <= n3681_1;
    Ng1365 <= n3686_1;
    Ng1372 <= n3691_1;
    Ng1378 <= n3696_1;
    Ng1385 <= n3701_1;
    Ng1386 <= n3706_1;
    Ng1384 <= n3711_1;
    Ng1388 <= n3716_1;
    Ng1389 <= n3721_1;
    Ng1387 <= n3726_1;
    Ng1391 <= n3731_1;
    Ng1392 <= n3736_1;
    Ng1390 <= n3741_1;
    Ng1394 <= n3746_1;
    Ng1395 <= n3751_1;
    Ng1393 <= n3756_1;
    Ng1397 <= n3761;
    Ng1398 <= n3766_1;
    Ng1396 <= n3771;
    Ng1400 <= n3776_1;
    Ng1401 <= n3781_1;
    Ng1399 <= n3786;
    Ng1403 <= n3791;
    Ng1404 <= n3796_1;
    Ng1402 <= n3801;
    Ng1406 <= n3806;
    Ng1407 <= n3811_1;
    Ng1405 <= n3816;
    Ng1409 <= n3821;
    Ng1410 <= n3826_1;
    Ng1408 <= n3831_1;
    Ng1412 <= n3836_1;
    Ng1413 <= n3841_1;
    Ng1411 <= n3846_1;
    Ng1415 <= n3851_1;
    Ng1416 <= n3856_1;
    Ng1414 <= n3861_1;
    Ng1418 <= n3866;
    Ng1419 <= n3871_1;
    Ng1417 <= n3876_1;
    Ng1421 <= n3881_1;
    Ng1422 <= n3886_1;
    Ng1420 <= n3891;
    Ng1424 <= n3896;
    Ng1425 <= n3901;
    Ng1423 <= n3906;
    Ng1512 <= n3911;
    Ng1513 <= n3916_1;
    Ng1511 <= n3921;
    Ng1515 <= n3926_1;
    Ng1516 <= n3931;
    Ng1514 <= n3936;
    Ng1524 <= n3941_1;
    Ng1525 <= n3946;
    Ng1523 <= n3951;
    Ng1527 <= n3956;
    Ng1528 <= n3961_1;
    Ng1526 <= n3966;
    Ng1530 <= n3971;
    Ng1531 <= n3976;
    Ng1529 <= n3981;
    Ng1533 <= n3986;
    Ng1534 <= n3991;
    Ng1532 <= n3996_1;
    Ng1536 <= n4001_1;
    Ng1537 <= n4006_1;
    Ng1535 <= n4011_1;
    Ng1539 <= n4016_1;
    Ng1540 <= n4021;
    Ng1538 <= n4026;
    Ng1542 <= n4031_1;
    Ng1543 <= n4036;
    Ng1541 <= n4041_1;
    Ng1545 <= n4046;
    Ng1546 <= n4051;
    Ng1544 <= n4056;
    Ng1551 <= n4061;
    Ng1552 <= n4066_1;
    Ng1550 <= n4071_1;
    Ng1554 <= n4076;
    Ng1555 <= n4081_1;
    Ng1553 <= n4086_1;
    Ng1557 <= n4091;
    Ng1558 <= n4096_1;
    Ng1556 <= n4101;
    Ng1560 <= n4106;
    Ng1561 <= n4111_1;
    Ng1559 <= n4116_1;
    Ng1567 <= n4121;
    Ng1570 <= n4126;
    Ng1573 <= n4131;
    Ng1612 <= n4136_1;
    Ng1615 <= n4141;
    Ng1618 <= n4146;
    Ng1576 <= n4151;
    Ng1579 <= n4156;
    Ng1582 <= n4161;
    Ng1621 <= n4166;
    Ng1624 <= n4171;
    Ng1627 <= n4176;
    Ng1585 <= n4181_1;
    Ng1588 <= n4186;
    Ng1591 <= n4191_1;
    Ng1630 <= n4196;
    Ng1633 <= n4201;
    Ng1636 <= n4206;
    Ng1594 <= n4211;
    Ng1597 <= n4216;
    Ng1600 <= n4221;
    Ng1639 <= n4226;
    Ng1642 <= n4231;
    Ng1645 <= n4236_1;
    Ng1603 <= n4241_1;
    Ng1606 <= n4246;
    Ng1609 <= n4251;
    Ng1648 <= n4256;
    Ng1651 <= n4261_1;
    Ng1654 <= n4266;
    Ng1466 <= n4271;
    Ng1462 <= n4276;
    Ng1457 <= n4281_1;
    Ng1453 <= n4286;
    Ng1448 <= n4291_1;
    Ng1444 <= n4296;
    Ng1439 <= n4301;
    Ng1435 <= n4306_1;
    Ng1430 <= n4311_1;
    Ng1426 <= n4316;
    Ng11551 <= n4321;
    Ng11552 <= n4326;
    Ng11553 <= n4331_1;
    Ng11554 <= n4336_1;
    Ng11555 <= n4341_1;
    Ng11556 <= n4346;
    Ng11557 <= n4351;
    Ng11558 <= n4356;
    Ng11559 <= n4361;
    Ng11560 <= n4366;
    Ng11561 <= n4371;
    Ng11562 <= n4376;
    Ng1789 <= n4381;
    Ng1792 <= n4386;
    Ng1795 <= n4391;
    Ng1798 <= n4396;
    Ng1801 <= n4401;
    Ng1804 <= n4406;
    Ng1808 <= n4411;
    Ng1809 <= n4416;
    Ng1807 <= n4421;
    Ng1810 <= n4426;
    Ng1813 <= n4431;
    Ng1816 <= n4436;
    Ng1819 <= n4441;
    Ng1822 <= n4446_1;
    Ng1825 <= n4451_1;
    Ng1829 <= n4456_1;
    Ng1830 <= n4461;
    Ng1828 <= n4466;
    Ng1693 <= n4471;
    Ng1694 <= n4476;
    Ng1695 <= n4481;
    Ng1696 <= n4486;
    Ng1697 <= n4491;
    Ng1698 <= n4496;
    Ng1699 <= n4501;
    Ng1700 <= n4506_1;
    Ng1701 <= n4511;
    Ng1703 <= n4516;
    Ng1704 <= n4521;
    Ng1702 <= n4526;
    Ng1784 <= n4531;
    Ng1785 <= n4536;
    Ng1783 <= n4541;
    Ng1831 <= n4546;
    Ng1832 <= n4550;
    Ng1833 <= n4555;
    Ng1834 <= n4559;
    Ng1835 <= n4564;
    Ng1660 <= n4568;
    Ng1661 <= n4573;
    Ng1662 <= n4577;
    Ng1663 <= n4582;
    Ng1664 <= n4586;
    Ng1665 <= n4591;
    Ng1666 <= n4595;
    Ng1667 <= n4600;
    Ng1668 <= n4604;
    Ng1669 <= n4609;
    Ng1670 <= n4613;
    Ng1671 <= n4617;
    Ng1672 <= n4621;
    Ng1680 <= n4626;
    Ng1686 <= n4631;
    Ng1679 <= n4636;
    Ng1723 <= n4640;
    Ng1730 <= n4644_1;
    Ng1731 <= n4648;
    Ng1732 <= n4652;
    Ng1733 <= n4656;
    Ng1734 <= n4660;
    Ng1738 <= n4664;
    Ng1745 <= n4668;
    Ng1746 <= n4672;
    Ng1747 <= n4676;
    Ng1748 <= n4680;
    Ng1749 <= n4684;
    Ng1753 <= n4688;
    Ng1760 <= n4692;
    Ng1761 <= n4696;
    Ng1762 <= n4700;
    Ng1763 <= n4704;
    Ng1764 <= n4708;
    Ng1768 <= n4712;
    Ng1775 <= n4716;
    Ng1776 <= n4720;
    Ng1777 <= n4724;
    Ng1778 <= n4728;
    Ng1705 <= n4732;
    Ng1934 <= n4737;
    Ng1937 <= n4742;
    Ng1890 <= n4747;
    Ng1893 <= n4752;
    Ng1903 <= n4756;
    Ng1904 <= n4760;
    Ng1944 <= n4765;
    Ng1949 <= n4769;
    Ng1950 <= n4774;
    Ng1951 <= n4778;
    Ng1952 <= n4783;
    Ng1953 <= n4787;
    Ng1954 <= n4792;
    Ng1945 <= n4796;
    Ng1946 <= n4801;
    Ng1947 <= n4805;
    Ng1948 <= n4810;
    Ng1870 <= n4814;
    Ng1867 <= n4819;
    Ng1868 <= n4824;
    Ng1869 <= n4829;
    Ng11566 <= n4834;
    Ng11569 <= n4838;
    Ng11570 <= n4842;
    Ng1858 <= n4846;
    Ng1859 <= n4851;
    Ng1860 <= n4856;
    Ng1861 <= n4861;
    Ng1865 <= n4866;
    Ng1845 <= n4871_1;
    Ng11571 <= n4876;
    Ng11567 <= n4880;
    Ng11568 <= n4884;
    Ng1908 <= n4888;
    Ng1915 <= n4892;
    Ng1922 <= n4896_1;
    Ng1923 <= n4901;
    Ng1924 <= n4905_1;
    Ng1928 <= n4910;
    Ng1929 <= n4915;
    Ng8302 <= n4919;
    Ng1938 <= n4924;
    Ng1939 <= n4928;
    Ng1956 <= n4933;
    Ng1957 <= n4938;
    Ng1955 <= n4943;
    Ng1959 <= n4948;
    Ng1960 <= n4953;
    Ng1958 <= n4958;
    Ng1962 <= n4963;
    Ng1963 <= n4968;
    Ng1961 <= n4973;
    Ng1965 <= n4978;
    Ng1966 <= n4983;
    Ng1964 <= n4988;
    Ng1967 <= n4993;
    Ng1970 <= n4998;
    Ng1973 <= n5003;
    Ng1976 <= n5008;
    Ng1979 <= n5013;
    Ng1982 <= n5018;
    Ng1994 <= n5023;
    Ng1997 <= n5028;
    Ng2000 <= n5033;
    Ng1985 <= n5038;
    Ng1988 <= n5043;
    Ng1991 <= n5048;
    Ng1871 <= n5053;
    Ng1874 <= n5058;
    Ng1877 <= n5063;
    Ng1886 <= n5067;
    Ng1887 <= n5072;
    Pg16399 <= n5077;
    Ng1905 <= n5080;
    Ng1909 <= n5085;
    Ng1910 <= n5090;
    Ng1911 <= n5095;
    Ng1912 <= n5100;
    Ng1913 <= n5105;
    Ng1914 <= n5110;
    Ng1916 <= n5115;
    Ng1917 <= n5120;
    Ng1918 <= n5125;
    Ng1921 <= n5130;
    Ng2010 <= n5135;
    Ng2039 <= n5140;
    Ng2020 <= n5145;
    Ng2013 <= n5150;
    Ng2033 <= n5155;
    Ng2026 <= n5160;
    Ng2040 <= n5165;
    Ng2052 <= n5170;
    Ng2046 <= n5175;
    Ng2059 <= n5180;
    Ng2066 <= n5185;
    Ng2072 <= n5190;
    Ng2079 <= n5195;
    Ng2080 <= n5200;
    Ng2078 <= n5205;
    Ng2082 <= n5210;
    Ng2083 <= n5215;
    Ng2081 <= n5220;
    Ng2085 <= n5225;
    Ng2086 <= n5230;
    Ng2084 <= n5235;
    Ng2088 <= n5240;
    Ng2089 <= n5245;
    Ng2087 <= n5250;
    Ng2091 <= n5255;
    Ng2092 <= n5260;
    Ng2090 <= n5265;
    Ng2094 <= n5270;
    Ng2095 <= n5275;
    Ng2093 <= n5280;
    Ng2097 <= n5285;
    Ng2098 <= n5290;
    Ng2096 <= n5295;
    Ng2100 <= n5300;
    Ng2101 <= n5305;
    Ng2099 <= n5310;
    Ng2103 <= n5315;
    Ng2104 <= n5320;
    Ng2102 <= n5325;
    Ng2106 <= n5330;
    Ng2107 <= n5335;
    Ng2105 <= n5340;
    Ng2109 <= n5345;
    Ng2110 <= n5350;
    Ng2108 <= n5355;
    Ng2112 <= n5360;
    Ng2113 <= n5365;
    Ng2111 <= n5370;
    Ng2115 <= n5375;
    Ng2116 <= n5380;
    Ng2114 <= n5385;
    Ng2118 <= n5390;
    Ng2119 <= n5395;
    Ng2117 <= n5400;
    Ng2206 <= n5405;
    Ng2207 <= n5410;
    Ng2205 <= n5415;
    Ng2209 <= n5420;
    Ng2210 <= n5425;
    Ng2208 <= n5430;
    Ng2218 <= n5435;
    Ng2219 <= n5440;
    Ng2217 <= n5445;
    Ng2221 <= n5450;
    Ng2222 <= n5455;
    Ng2220 <= n5460;
    Ng2224 <= n5465;
    Ng2225 <= n5470;
    Ng2223 <= n5475;
    Ng2227 <= n5480;
    Ng2228 <= n5485;
    Ng2226 <= n5490;
    Ng2230 <= n5495;
    Ng2231 <= n5500;
    Ng2229 <= n5505;
    Ng2233 <= n5510;
    Ng2234 <= n5515;
    Ng2232 <= n5520;
    Ng2236 <= n5525;
    Ng2237 <= n5530;
    Ng2235 <= n5535;
    Ng2239 <= n5540;
    Ng2240 <= n5545;
    Ng2238 <= n5550;
    Ng2245 <= n5555;
    Ng2246 <= n5560;
    Ng2244 <= n5565;
    Ng2248 <= n5570;
    Ng2249 <= n5575;
    Ng2247 <= n5580;
    Ng2251 <= n5585;
    Ng2252 <= n5590;
    Ng2250 <= n5595;
    Ng2254 <= n5600;
    Ng2255 <= n5605;
    Ng2253 <= n5610;
    Ng2261 <= n5615;
    Ng2264 <= n5620;
    Ng2267 <= n5625;
    Ng2306 <= n5630;
    Ng2309 <= n5635;
    Ng2312 <= n5640;
    Ng2270 <= n5645;
    Ng2273 <= n5650;
    Ng2276 <= n5655;
    Ng2315 <= n5660;
    Ng2318 <= n5665;
    Ng2321 <= n5670;
    Ng2279 <= n5675;
    Ng2282 <= n5680;
    Ng2285 <= n5685;
    Ng2324 <= n5690;
    Ng2327 <= n5695;
    Ng2330 <= n5700;
    Ng2288 <= n5705;
    Ng2291 <= n5710;
    Ng2294 <= n5715;
    Ng2333 <= n5720;
    Ng2336 <= n5725;
    Ng2339 <= n5730;
    Ng2297 <= n5735;
    Ng2300 <= n5740;
    Ng2303 <= n5745;
    Ng2342 <= n5750;
    Ng2345 <= n5755;
    Ng2348 <= n5760;
    Ng2160 <= n5765;
    Ng2156 <= n5770;
    Ng2151 <= n5775;
    Ng2147 <= n5780;
    Ng2142 <= n5785;
    Ng2138 <= n5790;
    Ng2133 <= n5795;
    Ng2129 <= n5800;
    Ng2124 <= n5805;
    Ng2120 <= n5810;
    Ng2256 <= n5815;
    \[1609]  <= n5819;
    Ng2257 <= n5823;
    Ng11578 <= n5828;
    Ng11579 <= n5833;
    Ng11580 <= n5838;
    Ng11581 <= n5843;
    Ng11582 <= n5848;
    Ng11583 <= n5853;
    Ng11584 <= n5858;
    Ng11585 <= n5863;
    Ng11586 <= n5868;
    Ng11587 <= n5873;
    Ng11588 <= n5878;
    Ng11589 <= n5883;
    Ng2483 <= n5888;
    Ng2486 <= n5893;
    Ng2489 <= n5898;
    Ng2492 <= n5903;
    Ng2495 <= n5908;
    Ng2498 <= n5913;
    Ng2502 <= n5918;
    Ng2503 <= n5923;
    Ng2501 <= n5928;
    Ng2504 <= n5933;
    Ng2507 <= n5938;
    Ng2510 <= n5943;
    Ng2513 <= n5948;
    Ng2516 <= n5953;
    Ng2519 <= n5958;
    Ng2523 <= n5963;
    Ng2524 <= n5968;
    Ng2522 <= n5973;
    Ng2387 <= n5978;
    Ng2388 <= n5983;
    Ng2389 <= n5988;
    Ng2390 <= n5993;
    Ng2391 <= n5998;
    Ng2392 <= n6003;
    Ng2393 <= n6008;
    Ng2394 <= n6013;
    Ng2395 <= n6018;
    Ng2397 <= n6023;
    Ng2398 <= n6028;
    Ng2396 <= n6033;
    Ng2478 <= n6038;
    Ng2479 <= n6043;
    Ng2477 <= n6048;
    Ng2525 <= n6053;
    Ng2526 <= n6057;
    Ng2527 <= n6062;
    Ng2528 <= n6066;
    Ng2529 <= n6071;
    Ng2354 <= n6075;
    Ng2355 <= n6080;
    Ng2356 <= n6084;
    Ng2357 <= n6089;
    Ng2358 <= n6093;
    Ng2359 <= n6098;
    Ng2360 <= n6102;
    Ng2361 <= n6107;
    Ng2362 <= n6111;
    Ng2363 <= n6116;
    Ng2364 <= n6120;
    Ng2365 <= n6124;
    Ng2366 <= n6128;
    Ng2374 <= n6133;
    Ng2380 <= n6138;
    Ng2373 <= n6143;
    Ng2417 <= n6147;
    Ng2424 <= n6151;
    Ng2425 <= n6155;
    Ng2426 <= n6159;
    Ng2427 <= n6163;
    Ng2428 <= n6167;
    Ng2432 <= n6171;
    Ng2439 <= n6175;
    Ng2440 <= n6179;
    Ng2441 <= n6183;
    Ng2442 <= n6187;
    Ng2443 <= n6191;
    Ng2447 <= n6195;
    Ng2454 <= n6199;
    Ng2455 <= n6203;
    Ng2456 <= n6207;
    Ng2457 <= n6211;
    Ng2458 <= n6215;
    Ng2462 <= n6219;
    Ng2469 <= n6223;
    Ng2470 <= n6227;
    Ng2471 <= n6231;
    Ng2472 <= n6235;
    Ng2399 <= n6239;
    Ng2628 <= n6244;
    Ng2631 <= n6249;
    Ng2584 <= n6254;
    Ng2587 <= n6259;
    Ng2597 <= n6263;
    Ng2598 <= n6267;
    Ng2638 <= n6272;
    Ng2643 <= n6276;
    Ng2644 <= n6281;
    Ng2645 <= n6285;
    Ng2646 <= n6290;
    Ng2647 <= n6294;
    Ng2648 <= n6299;
    Ng2639 <= n6303;
    Ng2640 <= n6308;
    Ng2641 <= n6312;
    Ng2642 <= n6317;
    Ng2564 <= n6321;
    Ng2561 <= n6326;
    Ng2562 <= n6331;
    Ng2563 <= n6336;
    Ng11593 <= n6341;
    Ng11596 <= n6345;
    Ng11597 <= n6349;
    Ng2552 <= n6353;
    Ng2553 <= n6358;
    Ng2554 <= n6363;
    Ng2555 <= n6368;
    Ng2559 <= n6373;
    Ng2539 <= n6378;
    Ng11598 <= n6383;
    Ng11594 <= n6387;
    Ng11595 <= n6391;
    Ng2602 <= n6395;
    Ng2609 <= n6399;
    Ng2616 <= n6403;
    Ng2617 <= n6408;
    Ng2618 <= n6412;
    Ng2622 <= n6417;
    Ng2623 <= n6422;
    Ng8311 <= n6426;
    Ng2632 <= n6431;
    Ng2633 <= n6435;
    Ng2650 <= n6440;
    Ng2651 <= n6445;
    Ng2649 <= n6450;
    Ng2653 <= n6455;
    Ng2654 <= n6460;
    Ng2652 <= n6465;
    Ng2656 <= n6470;
    Ng2657 <= n6475;
    Ng2655 <= n6480;
    Ng2659 <= n6485;
    Ng2660 <= n6490;
    Ng2658 <= n6495;
    Ng2661 <= n6500;
    Ng2664 <= n6505;
    Ng2667 <= n6510;
    Ng2670 <= n6515;
    Ng2673 <= n6520;
    Ng2676 <= n6525;
    Ng2688 <= n6530;
    Ng2691 <= n6535;
    Ng2694 <= n6540;
    Ng2679 <= n6545;
    Ng2682 <= n6550;
    Ng2685 <= n6555;
    Ng2565 <= n6560;
    Ng2568 <= n6565;
    Ng2571 <= n6570;
    Ng2580 <= n6574;
    Ng2581 <= n6579;
    Pg16437 <= n6584;
    Ng2599 <= n6587;
    Ng2603 <= n6592;
    Ng2604 <= n6597;
    Ng2605 <= n6602;
    Ng2606 <= n6607;
    Ng2607 <= n6612;
    Ng2608 <= n6617;
    Ng2610 <= n6622;
    Ng2611 <= n6627;
    Ng2612 <= n6632;
    Ng2615 <= n6637;
    Ng2704 <= n6642;
    Ng2733 <= n6647;
    Ng2714 <= n6652;
    Ng2707 <= n6657;
    Ng2727 <= n6662;
    Ng2720 <= n6667;
    Ng2734 <= n6672;
    Ng2746 <= n6677;
    Ng2740 <= n6682;
    Ng2753 <= n6687;
    Ng2760 <= n6692;
    Ng2766 <= n6697;
    Ng2773 <= n6702;
    Ng2774 <= n6707;
    Ng2772 <= n6712;
    Ng2776 <= n6717;
    Ng2777 <= n6722;
    Ng2775 <= n6727;
    Ng2779 <= n6732;
    Ng2780 <= n6737;
    Ng2778 <= n6742;
    Ng2782 <= n6747;
    Ng2783 <= n6752;
    Ng2781 <= n6757;
    Ng2785 <= n6762;
    Ng2786 <= n6767;
    Ng2784 <= n6772;
    Ng2788 <= n6777;
    Ng2789 <= n6782;
    Ng2787 <= n6787;
    Ng2791 <= n6792;
    Ng2792 <= n6797;
    Ng2790 <= n6802;
    Ng2794 <= n6807;
    Ng2795 <= n6812;
    Ng2793 <= n6817;
    Ng2797 <= n6822;
    Ng2798 <= n6827;
    Ng2796 <= n6832;
    Ng2800 <= n6837;
    Ng2801 <= n6842;
    Ng2799 <= n6847;
    Ng2803 <= n6852;
    Ng2804 <= n6857;
    Ng2802 <= n6862;
    Ng2806 <= n6867;
    Ng2807 <= n6872;
    Ng2805 <= n6877;
    Ng2809 <= n6882;
    Ng2810 <= n6887;
    Ng2808 <= n6892;
    Ng2812 <= n6897;
    Ng2813 <= n6902;
    Ng2811 <= n6907;
    Ng3054 <= n6912;
    Ng3079 <= n6917;
    Ng13475 <= n6922;
    Ng3043 <= n6926;
    Ng3044 <= n6931;
    Ng3045 <= n6936;
    Ng3046 <= n6941;
    Ng3047 <= n6946;
    Ng3048 <= n6951;
    Ng3049 <= n6956;
    Ng3050 <= n6961;
    Ng3051 <= n6966;
    Ng3052 <= n6971;
    Ng3053 <= n6976;
    Ng3055 <= n6981;
    Ng3056 <= n6986;
    Ng3057 <= n6991;
    Ng3058 <= n6996;
    Ng3059 <= n7001;
    Ng3060 <= n7006;
    Ng3061 <= n7011;
    Ng3062 <= n7016;
    Ng3063 <= n7021;
    Ng3064 <= n7026;
    Ng3065 <= n7031;
    Ng3066 <= n7036;
    Ng3067 <= n7041;
    Ng3068 <= n7046;
    Ng3069 <= n7051;
    Ng3070 <= n7056;
    Ng3071 <= n7061;
    Ng3072 <= n7066;
    Ng3073 <= n7071;
    Ng3074 <= n7076;
    Ng3075 <= n7081;
    Ng3076 <= n7086;
    Ng3077 <= n7091;
    Ng3078 <= n7096;
    Ng2997 <= n7101;
    Ng2993 <= n7106;
    Ng2998 <= n7111;
    Ng3006 <= n7116;
    Ng3002 <= n7121;
    Ng3013 <= n7126;
    Ng3010 <= n7131;
    Ng3024 <= n7136;
    Ng3018 <= n7141;
    Ng3028 <= n7146;
    Ng3036 <= n7151;
    Ng3032 <= n7156;
    Pg5388 <= n7160;
    Ng2986 <= n7163;
    Ng2987 <= n7167;
    Pg8275 <= n7172;
    Pg8274 <= n7176;
    Pg8273 <= n7180;
    Pg8272 <= n7184;
    Pg8268 <= n7188;
    Pg8269 <= n7192;
    Pg8270 <= n7196;
    Pg8271 <= n7200;
    Ng3083 <= n7204;
    Pg8267 <= n7209;
    Ng2992 <= n7213;
    Pg8266 <= n7218;
    Pg8265 <= n7222;
    Pg8264 <= n7226;
    Pg8262 <= n7230;
    Pg8263 <= n7234;
    Pg8260 <= n7238;
    Pg8261 <= n7242;
    Pg8259 <= n7246;
    Ng2990 <= n7250;
    Ng2991 <= n7255;
    Pg8258 <= n7260;
  end
endmodule


