// Benchmark "TOP" written by ABC on Tue Mar  5 09:54:52 2019

module apex2 ( 
    i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_,
    i_11_, i_12_, i_13_, i_14_, i_16_, i_17_, i_18_, i_19_, i_20_,
    i_21_, i_22_, i_23_, i_24_, i_25_, i_26_, i_27_, i_28_, i_29_, i_30_,
    i_31_, i_32_, i_33_, i_34_, i_35_, i_36_, i_37_, i_38_,
    o_0_, o_1_, o_2_  );
  input  i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_,
    i_10_, i_11_, i_12_, i_13_, i_14_, i_16_, i_17_, i_18_, i_19_,
    i_20_, i_21_, i_22_, i_23_, i_24_, i_25_, i_26_, i_27_, i_28_, i_29_,
    i_30_, i_31_, i_32_, i_33_, i_34_, i_35_, i_36_, i_37_, i_38_;
  output o_0_, o_1_, o_2_;
  wire n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
    n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
    n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
    n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
    n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
    n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
    n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
    n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
    n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
    n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
    n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
    n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
    n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
    n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
    n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
    n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
    n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
    n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
    n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
    n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
    n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
    n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
    n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
    n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
    n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
    n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
    n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
    n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
    n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
    n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
    n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
    n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
    n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
    n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
    n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
    n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
    n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
    n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
    n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
    n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
    n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
    n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
    n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
    n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
    n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
    n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
    n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
    n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
    n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
    n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
    n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
    n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
    n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
    n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
    n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
    n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
    n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
    n977, n978, n979, n980, n981, n982, n983;
  assign o_0_ = ~n965 | ~n966 | n49 | ~n964 | n47 | n48 | n45 | n46;
  assign o_1_ = ~n603;
  assign o_2_ = ~n350;
  assign n45 = ~n798 & n686 & n229 & ~n379;
  assign n46 = ~n684 & n528 & i_35_ & n526;
  assign n47 = ~n693 & ~n805 & (~i_13_ | ~i_14_);
  assign n48 = ~n524 & (~n939 | (~n205 & ~n473));
  assign n49 = n804 | ~n968 | n734 | n736 | n732 | n733 | ~n208 | n731;
  assign n50 = ~i_27_ & ~n161;
  assign n51 = ~i_30_ & n300;
  assign n52 = i_36_ & (~n938 | (n50 & n51));
  assign n53 = ~i_12_ & ~i_13_;
  assign n54 = ~i_7_ & (n53 | ~n803);
  assign n55 = ~i_11_ & ~i_19_;
  assign n56 = ~i_24_ & (~n80 | (n55 & ~n81));
  assign n57 = i_19_ & ~i_13_ & i_18_;
  assign n58 = ~i_13_ & i_18_;
  assign n59 = ~i_22_ & (n57 | (i_11_ & n58));
  assign n60 = ~i_24_ & (~n86 | (n55 & ~n87));
  assign n61 = i_17_ & i_12_;
  assign n62 = i_14_ & i_13_;
  assign n63 = i_22_ & (n61 | n62);
  assign n64 = ~i_10_ & ~i_24_;
  assign n65 = ~n90 & (n64 | (i_13_ & ~i_24_));
  assign n66 = ~i_24_ & (n61 | n62);
  assign n67 = n610 | i_1_ | n746;
  assign n68 = ~i_18_ | ~n237;
  assign n69 = i_6_ | n113;
  assign n70 = (n68 | n69) & (n67 | ~n237);
  assign n71 = i_11_ & ~i_13_;
  assign n72 = n71 & (~n773 | (i_18_ & ~n149));
  assign n73 = i_9_ & n71;
  assign n74 = n73 & (~n67 | (i_18_ & ~n69));
  assign n75 = ~n635 | ~n280 | ~n324;
  assign n76 = ~n324 | n747;
  assign n77 = n75 & (n76 | ~n128);
  assign n78 = ~n280 | n106 | n140;
  assign n79 = n78 & (~n128 | ~n259 | ~n328);
  assign n80 = n764 | i_9_ | i_18_;
  assign n81 = n313 | n100;
  assign n82 = n80 & (~n55 | n81);
  assign n83 = n113 | i_6_ | n744;
  assign n84 = n316 | n745;
  assign n85 = n83 & (~i_9_ | n84);
  assign n86 = i_18_ | n759;
  assign n87 = n313 | n98;
  assign n88 = n86 & (~n55 | n87);
  assign n89 = i_10_ & ~i_13_;
  assign n90 = i_9_ | n760;
  assign n91 = (i_32_ | n88) & (n89 | n90);
  assign n92 = n754 | ~i_9_ | n745;
  assign n93 = ~i_11_ | i_12_;
  assign n94 = ~i_11_ | n744;
  assign n95 = (n67 | n94) & (n92 | n93);
  assign n96 = (~n73 | n84) & (~n71 | n83);
  assign n97 = (~i_18_ | n96) & (i_13_ | n95);
  assign n98 = i_7_ | n763;
  assign n99 = i_32_ | ~i_38_;
  assign n100 = i_8_ | n763;
  assign n101 = (n98 | n99) & (n100 | ~n262);
  assign n102 = ~n278 | n98 | n107;
  assign n103 = ~n328 | n100 | n116;
  assign n104 = i_25_ | n743;
  assign n105 = n102 & n103 & (n101 | n104);
  assign n106 = i_32_ | ~n324;
  assign n107 = i_32_ | n743;
  assign n108 = (n104 | n106) & (n107 | ~n328);
  assign n109 = n757 | n419;
  assign n110 = n313 | n765;
  assign n111 = (i_19_ | n110) & (i_18_ | n109);
  assign n112 = n316 | n468;
  assign n113 = i_12_ | n313;
  assign n114 = i_6_ | ~n214;
  assign n115 = (n113 | n114) & (i_8_ | n112);
  assign n116 = i_31_ | n743;
  assign n117 = i_35_ | n749;
  assign n118 = n117 | n116 | n111;
  assign n119 = ~n262 | i_32_ | n111;
  assign n120 = n119 & (i_2_ | ~n259 | ~n324);
  assign n121 = ~n104 | ~n971;
  assign n122 = i_38_ & (~n118 | (~n115 & n121));
  assign n123 = n867 & (~n635 | n774);
  assign n124 = (~i_38_ | n91) & (n82 | ~n262);
  assign n125 = n866 & (i_10_ | n85 | ~n324);
  assign n126 = n123 & (i_28_ | (n124 & n125));
  assign n127 = ~i_24_ & (~n869 | ~n871 | ~n873);
  assign n128 = ~i_28_ & ~n161;
  assign n129 = n128 & (~n876 | ~n878 | ~n880);
  assign n130 = ~n271 | i_30_ | n160;
  assign n131 = (n190 | ~n269) & (n104 | n768);
  assign n132 = ~i_38_ | n762;
  assign n133 = n130 & n131 & (~n51 | n132);
  assign n134 = i_28_ | n175;
  assign n135 = i_22_ | ~n257;
  assign n136 = n143 | ~n324;
  assign n137 = (n135 | n136) & (n134 | ~n269);
  assign n138 = n135 | n143;
  assign n139 = n175 | ~n328;
  assign n140 = i_28_ | i_31_ | i_30_;
  assign n141 = (n139 | n140) & (n138 | ~n262);
  assign n142 = n104 | i_30_ | ~i_38_;
  assign n143 = i_30_ | n743;
  assign n144 = n142 & (n143 | ~n278);
  assign n145 = (~n64 | n83) & (n84 | ~n272);
  assign n146 = ~i_18_ | ~n257;
  assign n147 = i_13_ | ~n257;
  assign n148 = (n95 | n147) & (n96 | n146);
  assign n149 = n742 | n316;
  assign n150 = i_10_ | i_6_ | ~i_9_;
  assign n151 = (n113 | n150) & (i_10_ | n149);
  assign n152 = ~n262 | i_8_ | i_30_;
  assign n153 = n119 & (n89 | n101 | n313);
  assign n154 = n152 & n153 & (n151 | n106);
  assign n155 = ~n65 & (i_32_ | ~n60);
  assign n156 = n155 & (i_30_ | ~n336);
  assign n157 = (n156 | ~n278) & (~n56 | n282);
  assign n158 = n865 & (n76 | ~n272);
  assign n159 = n157 & n158 & (n154 | ~n257);
  assign n160 = ~i_34_ | ~n324;
  assign n161 = i_24_ | i_26_;
  assign n162 = (n161 | ~n328) & (n160 | ~n257);
  assign n163 = n98 | n161 | ~n278 | ~n310;
  assign n164 = n162 | n167;
  assign n165 = i_31_ | i_33_ | n160 | ~n267;
  assign n166 = n163 & (n100 | (n164 & n165));
  assign n167 = i_31_ | ~n300;
  assign n168 = (n116 | n135) & (n167 | ~n280);
  assign n169 = (n160 | ~n265) & (~n128 | ~n328);
  assign n170 = n750 | n160 | ~n267;
  assign n171 = (i_31_ | n199) & (n168 | n106);
  assign n172 = i_29_ | n541;
  assign n173 = n170 & n171 & (n169 | n172);
  assign n174 = n135 | n143 | i_32_ | ~i_38_;
  assign n175 = i_22_ | n161;
  assign n176 = n174 & (n175 | ~n278 | ~n635);
  assign n177 = n176 | n761;
  assign n178 = i_3_ | i_8_ | ~i_10_ | n141;
  assign n179 = i_3_ | n744;
  assign n180 = n177 & n178 & (n137 | n179);
  assign n181 = (i_29_ | ~n128) & (i_28_ | n175);
  assign n182 = i_2_ | n744;
  assign n183 = i_24_ | ~i_12_ | i_22_;
  assign n184 = i_10_ | n744;
  assign n185 = (n183 | n184) & (n182 | ~n342);
  assign n186 = i_26_ | ~i_38_ | ~n51 | n117;
  assign n187 = i_29_ | ~n219;
  assign n188 = n186 & (i_28_ | n187 | n132);
  assign n189 = ~n654 | ~i_38_ | ~n51;
  assign n190 = i_26_ | ~n300;
  assign n191 = i_30_ | n106;
  assign n192 = n189 & (n190 | n191);
  assign n193 = ~i_19_ | i_24_;
  assign n194 = ~i_19_ | ~n257;
  assign n195 = (n192 | n194) & (n188 | n193);
  assign n196 = (n107 | n135) & (~n265 | n509);
  assign n197 = (~n128 | n224) & (~n267 | n318);
  assign n198 = n196 & n197 & (~n280 | ~n310);
  assign n199 = n139 | i_32_ | i_28_;
  assign n200 = n199 & (n198 | ~n324);
  assign n201 = ~i_31_ | ~n235;
  assign n202 = n201 & (~n235 | (~i_30_ & ~i_32_));
  assign n203 = i_23_ | ~n739;
  assign n204 = i_27_ | n740;
  assign n205 = ~i_14_ | n580;
  assign n206 = (n204 | n205) & (n203 | ~n307);
  assign n207 = n684 | n738 | ~i_20_ | ~n537;
  assign n208 = n207 & (n206 | ~n235 | ~n531);
  assign n209 = i_22_ | ~n237;
  assign n210 = ~n59 & (i_3_ | n209);
  assign n211 = (i_8_ | n141) & (i_7_ | n176);
  assign n212 = (n79 | n210) & (n211 | n68);
  assign n213 = ~i_22_ & ~n193;
  assign n214 = ~i_7_ & ~i_8_;
  assign n215 = n214 & ~n144 & n213;
  assign n216 = i_12_ & n58;
  assign n217 = n216 & (n215 | (i_11_ & ~n211));
  assign n218 = ~i_34_ | n769;
  assign n219 = ~i_30_ & ~i_32_;
  assign n220 = n218 & (i_28_ | ~i_34_ | n219);
  assign n221 = (~i_22_ | n220) & (n219 | ~n303);
  assign n222 = i_29_ | n572;
  assign n223 = n221 & (i_28_ | n222);
  assign n224 = i_29_ | n749;
  assign n225 = (i_28_ | n224) & (i_25_ | ~n310);
  assign n226 = i_31_ | n752;
  assign n227 = (i_8_ | n226) & (n111 | n172);
  assign n228 = i_33_ & n235;
  assign n229 = i_33_ & i_34_;
  assign n230 = i_14_ & (n228 | (~i_24_ & n229));
  assign n231 = n785 & n112;
  assign n232 = i_2_ | ~n214;
  assign n233 = (i_30_ | n232) & (i_32_ | n231);
  assign n234 = i_22_ & (n230 | (~n202 & n203));
  assign n235 = ~i_34_ & i_35_;
  assign n236 = ~n259 & (~n853 | (n63 & n235));
  assign n237 = ~i_13_ & i_19_;
  assign n238 = ~n179 & (n71 | n237);
  assign n239 = ~i_24_ & (n238 | (n58 & ~n94));
  assign n240 = i_13_ | n744;
  assign n241 = ~n239 & (~i_18_ | n193 | n240);
  assign n242 = n68 & (~i_18_ | ~n71);
  assign n243 = (n94 | ~n216) & (n182 | n242);
  assign n244 = ~i_12_ | n744;
  assign n245 = n243 & (n68 | n244);
  assign n246 = i_12_ & n71;
  assign n247 = n246 & i_18_ & ~i_22_;
  assign n248 = ~n761 & n213 & ~i_13_ & ~i_8_ & i_12_;
  assign n249 = (n106 | n138) & (n139 | ~n635);
  assign n250 = (n77 | n210) & (i_7_ | n176);
  assign n251 = ~i_10_ & ~n249 & (~i_2_ | i_12_);
  assign n252 = ~i_3_ & i_11_;
  assign n253 = ~i_22_ & i_12_ & ~i_13_;
  assign n254 = n252 & (~n847 | (~n77 & n253));
  assign n255 = (~n55 | n90) & (i_8_ | n86);
  assign n256 = ~n225 & ~n89 & ~i_24_ & ~n87;
  assign n257 = ~i_24_ & ~i_25_;
  assign n258 = n257 & n51 & ~i_7_ & ~i_32_;
  assign n259 = ~i_31_ & n219;
  assign n260 = (~i_22_ | ~i_23_) & (~n63 | n259);
  assign n261 = (~i_38_ | n155) & (~n56 | ~n262);
  assign n262 = ~i_31_ & n324;
  assign n263 = ~n823 & ~i_29_ & n262;
  assign n264 = i_8_ | ~n51 | ~n257 | ~n262;
  assign n265 = ~i_28_ & n257;
  assign n266 = n265 & (n263 | (~n184 & ~n768));
  assign n267 = ~i_24_ & n300;
  assign n268 = ~n823 & ~i_31_ & n328;
  assign n269 = ~i_30_ & n328;
  assign n270 = n267 & (n268 | (~n184 & n269));
  assign n271 = ~i_25_ & n300;
  assign n272 = n64 & i_9_;
  assign n273 = n271 & (~n261 | (~n191 & n272));
  assign n274 = i_29_ | n769;
  assign n275 = ~n66 | n274;
  assign n276 = i_38_ & (n256 | n258 | ~n842);
  assign n277 = (n104 | n261) & (n142 | ~n336);
  assign n278 = ~i_33_ & i_38_;
  assign n279 = n278 & ~i_7_ & ~n161;
  assign n280 = ~i_25_ & ~n161;
  assign n281 = ~i_32_ & (n279 | (n262 & n280));
  assign n282 = i_33_ | ~n262;
  assign n283 = ~n281 & (i_8_ | n161 | n282);
  assign n284 = ~i_25_ & (~n770 | (n51 & n214));
  assign n285 = ~n89 & (~n90 | (~i_32_ & ~n87));
  assign n286 = n829 & (~n310 | (~n280 & ~n299));
  assign n287 = n830 & (~n267 | n318);
  assign n288 = i_32_ | ~n235;
  assign n289 = n286 & n287 & (~n271 | n288);
  assign n290 = ~n190 & (~n115 | (~i_7_ & n219));
  assign n291 = n565 | n87 | ~n300;
  assign n292 = i_29_ | i_34_ | i_33_;
  assign n293 = n291 & (i_28_ | n90 | n292);
  assign n294 = (n117 | ~n128) & (~n265 | ~n654);
  assign n295 = i_33_ | n755;
  assign n296 = i_24_ | i_28_;
  assign n297 = i_33_ | ~n300;
  assign n298 = (n161 | n297) & (n295 | n296);
  assign n299 = ~i_33_ & n235;
  assign n300 = ~i_28_ & ~i_29_;
  assign n301 = ~n115 & (~n298 | (n299 & n300));
  assign n302 = ~n255 & (~n827 | (n280 & n300));
  assign n303 = n300 & i_34_;
  assign n304 = n257 & (~n828 | (~n115 & n303));
  assign n305 = n235 & (n284 | ~n832 | ~n834);
  assign n306 = ~i_27_ & n300;
  assign n307 = n53 & i_14_;
  assign n308 = ~i_16_ & n655;
  assign n309 = n308 & n306 & n307;
  assign n310 = ~i_32_ & n300;
  assign n311 = n310 & ~n151 & ~n161;
  assign n312 = (~n56 | n167) & (~n259 | ~n267);
  assign n313 = i_5_ | n741;
  assign n314 = i_12_ | i_6_;
  assign n315 = i_5_ | i_6_;
  assign n316 = i_1_ | n741;
  assign n317 = (n315 | n316) & (n313 | n314);
  assign n318 = ~i_34_ | n749;
  assign n319 = (~n272 | n318) & (n184 | ~n280);
  assign n320 = (i_29_ | n145) & (n187 | ~n272);
  assign n321 = ~i_24_ & ~n317 & (~n814 | ~n815);
  assign n322 = n213 & (~n104 | ~n971);
  assign n323 = (~n816 | ~n817) & (~n819 | ~n820);
  assign n324 = ~i_35_ & i_38_;
  assign n325 = n324 & (~n821 | ~n822 | ~n825);
  assign n326 = ~n181 & (n268 | (~n255 & n278));
  assign n327 = ~n180 & (n246 | (i_12_ & n237));
  assign n328 = ~i_33_ & n324;
  assign n329 = n328 & (n311 | (~n143 & ~n185));
  assign n330 = n306 & ~n473;
  assign n331 = n229 & (n309 | (~n205 & n330));
  assign n332 = n228 & n300 & n259;
  assign n333 = i_14_ & (n332 | (n128 & i_33_));
  assign n334 = i_9_ & (~n848 | ~n850 | ~n852);
  assign n335 = i_10_ & (n247 | (n252 & n253));
  assign n336 = ~i_24_ & n214;
  assign n337 = ~n144 & (n248 | (n335 & n336));
  assign n338 = ~i_28_ & (n234 | n236 | ~n975);
  assign n339 = i_10_ & (~n857 | (i_12_ & ~n212));
  assign n340 = n73 & (~n859 | (~n137 & ~n771));
  assign n341 = n203 & (~n860 | (n128 & ~n219));
  assign n342 = ~i_22_ & n64;
  assign n343 = ~n313 & (~n864 | (~n105 & n342));
  assign n344 = ~n325 & (~i_27_ | n175 | ~n421);
  assign n345 = n887 & (n77 | n209 | n748);
  assign n346 = n886 & (~n66 | n219 | ~n303);
  assign n347 = ~n333 & n890 & (~n51 | n283);
  assign n348 = ~n329 & n888 & (n132 | n312);
  assign n349 = n897 & n896 & n895 & n893 & n892 & n891 & ~n339 & ~n340;
  assign n350 = n349 & n348 & n347 & n346 & n345 & n344 & ~n326 & ~n327;
  assign n351 = ~i_34_ | ~i_37_;
  assign n352 = i_29_ | n510;
  assign n353 = ~i_37_ | ~n235;
  assign n354 = (n351 | n352) & (~n306 | n353);
  assign n355 = n523 | i_29_ | ~n427;
  assign n356 = ~i_34_ | ~n427;
  assign n357 = n355 & (~n306 | n356);
  assign n358 = ~n654 | ~i_37_ | ~n306;
  assign n359 = n358 & (i_32_ | n355);
  assign n360 = n793 | n313 | n361;
  assign n361 = i_17_ | n581;
  assign n362 = i_10_ | n763;
  assign n363 = n360 & (n313 | n361 | n362);
  assign n364 = n413 | n397 | n788 | n362;
  assign n365 = n488 | ~i_37_ | n468;
  assign n366 = n863 | ~n427 | n788;
  assign n367 = n364 & (n361 | (n365 & n366));
  assign n368 = n788 | ~n391 | n766;
  assign n369 = n778 | i_7_ | i_0_;
  assign n370 = n368 & (i_12_ | n369);
  assign n371 = ~i_23_ & ~n161;
  assign n372 = n371 & (~n921 | (~n370 & ~n493));
  assign n373 = n463 | n500 | n782;
  assign n374 = i_11_ | n581;
  assign n375 = n590 | n98 | n788;
  assign n376 = ~n372 & n373 & (n374 | n375);
  assign n377 = i_14_ | ~n427;
  assign n378 = (~i_21_ | ~n546) & (~n51 | n377);
  assign n379 = n737 & n361;
  assign n380 = n379 & (i_33_ | ~n544);
  assign n381 = n87 | n604;
  assign n382 = i_10_ | n581;
  assign n383 = n381 & (n87 | n382);
  assign n384 = n380 | n450 | ~i_31_ | ~n51;
  assign n385 = n384 & (~n330 | n383);
  assign n386 = n523 | n800 | ~i_29_ | n367;
  assign n387 = n796 | i_29_ | n690 | n444;
  assign n388 = (~i_37_ | n376) & (n351 | n385);
  assign n389 = n923 & (i_31_ | n378 | n540);
  assign n390 = n389 & n388 & n386 & n387;
  assign n391 = ~i_27_ & n421;
  assign n392 = n655 & i_22_;
  assign n393 = n391 & n392 & (~n379 | ~n784);
  assign n394 = ~i_33_ | n541;
  assign n395 = ~i_25_ | ~n655;
  assign n396 = ~n393 & (~n51 | n394 | n395);
  assign n397 = i_33_ | ~n427;
  assign n398 = n377 & (i_13_ | n397);
  assign n399 = n382 & n604;
  assign n400 = i_10_ | n580;
  assign n401 = (n397 | n400) & (n399 | ~n427);
  assign n402 = ~n365 & (~n485 | (~i_33_ & ~n474));
  assign n403 = i_20_ | ~n776;
  assign n404 = i_20_ | n740;
  assign n405 = (i_16_ | n404) & (i_12_ | n403);
  assign n406 = n900 & (n764 | n500 | n786);
  assign n407 = i_19_ | n740;
  assign n408 = n406 & (n81 | n407 | n374);
  assign n409 = n786 | n764 | n501;
  assign n410 = i_11_ | n580;
  assign n411 = n409 & (n81 | n407 | n410);
  assign n412 = n399 & (i_33_ | n400);
  assign n413 = i_17_ | n580;
  assign n414 = (n397 | n413) & (n361 | ~n427);
  assign n415 = n918 & (i_19_ | n765 | n417);
  assign n416 = n415 & (n398 | n314 | n403);
  assign n417 = n414 | i_23_ | i_20_;
  assign n418 = ~i_3_ | n780;
  assign n419 = i_9_ | n315;
  assign n420 = n419 | i_18_ | n417 | n418;
  assign n421 = ~i_28_ & i_29_;
  assign n422 = ~n404 & n421 & (n402 | ~n917);
  assign n423 = n438 | i_13_ | n787;
  assign n424 = n423 | ~n310 | n397;
  assign n425 = ~i_32_ & n421;
  assign n426 = n425 & (~n420 | (~n416 & ~n788));
  assign n427 = ~i_35_ & i_37_;
  assign n428 = n427 & (~n919 | (n310 & ~n556));
  assign n429 = n898 & (n758 | n501 | n786);
  assign n430 = n429 & (n87 | n407 | n410);
  assign n431 = i_18_ | ~n655;
  assign n432 = i_19_ | ~n655;
  assign n433 = (n110 | n432) & (n109 | n431);
  assign n434 = ~i_37_ | n749;
  assign n435 = i_30_ | ~i_31_ | n434 | ~n544;
  assign n436 = n362 | n313 | n413;
  assign n437 = n436 | ~i_37_ | n117;
  assign n438 = i_16_ | n740;
  assign n439 = i_13_ | ~n214;
  assign n440 = i_23_ | n580;
  assign n441 = i_12_ | ~n214;
  assign n442 = (n440 | n441) & (n438 | n439);
  assign n443 = n397 | n472 | ~i_34_ | ~n308;
  assign n444 = i_34_ | n566;
  assign n445 = n443 & (i_33_ | n442 | n444);
  assign n446 = n371 & (~n435 | ~n437 | ~n913);
  assign n447 = n915 & (n430 | n565 | n566);
  assign n448 = ~n446 & n447 & (i_30_ | n445);
  assign n449 = ~n659 | n690;
  assign n450 = i_27_ | ~n655;
  assign n451 = n449 & (~n303 | n450);
  assign n452 = n462 | i_8_ | n759;
  assign n453 = i_11_ | n783;
  assign n454 = n452 & (n90 | n453);
  assign n455 = i_7_ | i_28_ | n226 | n288;
  assign n456 = n495 | i_9_ | n89 | ~n537 | n789;
  assign n457 = n455 & n456 & (n451 | n454);
  assign n458 = (i_10_ | n90) & (i_30_ | ~n214);
  assign n459 = n438 | n354 | n458;
  assign n460 = n912 & (~n427 | n751 | n767);
  assign n461 = n459 & n460 & (~i_37_ | n457);
  assign n462 = i_18_ | n779;
  assign n463 = n468 | n418;
  assign n464 = n463 | n462 | i_8_;
  assign n465 = ~i_9_ & (~n464 | (~n453 & ~n789));
  assign n466 = n465 & (~i_14_ | (~i_13_ & ~i_33_));
  assign n467 = ~n789 & (~n737 | (~i_33_ & ~n784));
  assign n468 = i_7_ | n315;
  assign n469 = n434 | n413 | n468;
  assign n470 = ~n488 & (~n469 | (~n414 & ~n745));
  assign n471 = ~n470 & (~i_37_ | (~n466 & ~n467));
  assign n472 = i_8_ | ~n53;
  assign n473 = i_17_ | ~n655;
  assign n474 = i_8_ | n580;
  assign n475 = (n473 | n474) & (~n308 | n472);
  assign n476 = i_33_ | n752;
  assign n477 = n623 & n972;
  assign n478 = (n477 | n224) & (n475 | n476);
  assign n479 = ~n543 | n737;
  assign n480 = n969 & (~i_29_ | n471 | n800);
  assign n481 = n479 & n480 & (~n427 | n478);
  assign n482 = n394 | n799 | ~i_25_ | i_28_;
  assign n483 = n482 & (~n330 | n397 | n474);
  assign n484 = i_8_ | n803;
  assign n485 = i_8_ | n581;
  assign n486 = (~n308 | n484) & (n473 | n485);
  assign n487 = i_33_ | i_9_ | i_10_ | n789;
  assign n488 = i_1_ | n780;
  assign n489 = n487 & (n315 | n117 | n488);
  assign n490 = n434 | n369 | ~n371;
  assign n491 = n490 & (~i_37_ | n489 | ~n537);
  assign n492 = i_20_ | n580;
  assign n493 = i_20_ | n581;
  assign n494 = (~n427 | n493) & (n397 | n492);
  assign n495 = i_20_ | n779;
  assign n496 = (n398 | n495) & (i_12_ | n494);
  assign n497 = n299 & ~i_7_ & i_37_;
  assign n498 = n300 & (n497 | (i_25_ & n228));
  assign n499 = ~n498 & (~n235 | ~n421 | ~n738);
  assign n500 = i_9_ | n581;
  assign n501 = i_9_ | n580;
  assign n502 = (n397 | n501) & (~n427 | n500);
  assign n503 = (n356 | n423) & (n430 | n351);
  assign n504 = n760 | n784;
  assign n505 = n783 | i_11_ | n90;
  assign n506 = n504 & (i_13_ | (n505 & n452));
  assign n507 = n84 | n413;
  assign n508 = (n356 | n507) & (n506 | n351);
  assign n509 = i_32_ | n755;
  assign n510 = i_24_ | n777;
  assign n511 = (n509 | n510) & (n288 | ~n306);
  assign n512 = n907 & (n758 | n500 | n786);
  assign n513 = n512 & (n87 | n407 | n374);
  assign n514 = ~n310 | n450;
  assign n515 = n81 | n400;
  assign n516 = (n436 | n514) & (~n330 | n515);
  assign n517 = n204 | ~n310;
  assign n518 = (n318 | ~n330) & (~n299 | n517);
  assign n519 = (n511 | n513) & (n516 | n762);
  assign n520 = n908 & n909 & (n518 | n802);
  assign n521 = n760 | n737;
  assign n522 = n519 & n520 & (n451 | n521);
  assign n523 = i_26_ | n777;
  assign n524 = (~n229 | ~n306) & (~i_33_ | n523);
  assign n525 = ~n664 & i_25_ & i_20_ & ~i_23_;
  assign n526 = ~i_34_ & n421;
  assign n527 = ~i_27_ & n697;
  assign n528 = i_22_ & n797;
  assign n529 = i_35_ & n526 & (n527 | n528);
  assign n530 = i_25_ & n797;
  assign n531 = n300 & i_33_;
  assign n532 = n235 & (n525 | (n530 & n531));
  assign n533 = n906 & (~i_34_ | ~n391 | ~n686);
  assign n534 = ~n532 & n533 & (n395 | n524);
  assign n535 = ~n413 & i_34_ & n391;
  assign n536 = ~i_20_ & ~i_21_;
  assign n537 = n371 & n391;
  assign n538 = ~n737 | ~n784;
  assign n539 = n538 & n537 & n536 & i_2_;
  assign n540 = i_34_ | n161;
  assign n541 = i_31_ | i_32_;
  assign n542 = ~i_22_ | n540 | n541 | ~n546;
  assign n543 = i_29_ & n392;
  assign n544 = ~n413 | ~n784;
  assign n545 = ~n523 & n543 & (~n361 | n544);
  assign n546 = ~i_30_ & n421;
  assign n547 = n392 & (n535 | (n546 & ~n751));
  assign n548 = n112 | n413;
  assign n549 = n112 | n474;
  assign n550 = (n514 | n548) & (~n330 | n549);
  assign n551 = n905 & (n442 | n476 | n510);
  assign n552 = (~n330 | n794) & (n514 | n796);
  assign n553 = n551 & n552 & (i_33_ | n550);
  assign n554 = ~n655 | i_28_ | n318;
  assign n555 = n973 & n411;
  assign n556 = n438 | i_14_ | n787;
  assign n557 = (n509 | n556) & (n555 | n295);
  assign n558 = ~n226 & (~n554 | (n128 & ~n565));
  assign n559 = n795 | ~n303 | n450;
  assign n560 = ~n558 & n559 & (n510 | n557);
  assign n561 = (n297 | n549) & (~n310 | n383);
  assign n562 = n794 | ~n300 | n444;
  assign n563 = n562 & (n561 | n353);
  assign n564 = n379 | ~i_37_ | n288;
  assign n565 = i_34_ | n749;
  assign n566 = ~i_35_ | ~i_37_;
  assign n567 = n564 & (~n544 | n565 | n566);
  assign n568 = n492 | n370 | ~n371;
  assign n569 = n463 | n501 | n782;
  assign n570 = n568 & n569 & (n410 | n375);
  assign n571 = i_27_ | n769;
  assign n572 = ~i_31_ | ~i_34_;
  assign n573 = (~n235 | n571) & (n510 | n572);
  assign n574 = (~n306 | n572) & (~i_31_ | n523);
  assign n575 = n274 | n204 | ~n235;
  assign n576 = n740 | ~i_20_ | n573;
  assign n577 = n575 & n576 & (n574 | n473);
  assign n578 = n308 & ~n574;
  assign n579 = (n578 | ~n902) & (n53 | ~n803);
  assign n580 = i_16_ | i_13_;
  assign n581 = i_16_ | i_14_;
  assign n582 = ~n579 & (n577 | (n580 & n581));
  assign n583 = i_34_ | i_24_ | n143 | n394;
  assign n584 = n583 & (i_28_ | ~n228 | ~n259);
  assign n585 = ~n51 | n540;
  assign n586 = (~i_20_ | n584) & (n394 | n585);
  assign n587 = (n363 | n514) & (n408 | n352);
  assign n588 = (n397 | n410) & (n374 | ~n427);
  assign n589 = n753 | n494 | ~n537;
  assign n590 = i_19_ | n781;
  assign n591 = n589 & (n588 | n100 | n590);
  assign n592 = ~n308 | i_14_ | n69;
  assign n593 = n592 & (n433 | n361);
  assign n594 = ~i_30_ & (~n911 | (i_34_ & ~n483));
  assign n595 = n502 | n745 | n782 | n418;
  assign n596 = i_0_ | i_8_ | n496 | n709;
  assign n597 = n924 & (n503 | n224 | n510);
  assign n598 = n926 & n927 & (n473 | ~n899);
  assign n599 = (~i_25_ | n586) & (n356 | n587);
  assign n600 = (n591 | n788) & (n359 | n593);
  assign n601 = n928 & (n690 | (n904 & n929));
  assign n602 = n936 & n935 & n933 & n932 & n931 & n930 & ~n594 & ~n804;
  assign n603 = n602 & n601 & n600 & n599 & n598 & n597 & n595 & n596;
  assign n604 = ~i_13_ | n581;
  assign n605 = (i_12_ | n604) & (~i_13_ | n361);
  assign n606 = n413 & n361;
  assign n607 = (i_10_ | n413) & (~i_13_ | n361);
  assign n608 = i_5_ | ~i_3_ | i_4_;
  assign n609 = n608 | n462 | i_6_;
  assign n610 = i_4_ | n315;
  assign n611 = ~i_2_ & (i_8_ | n610 | ~n735);
  assign n612 = ~n610 & i_36_ & ~i_7_ & ~i_32_;
  assign n613 = ~n607 & (~n611 | n612);
  assign n614 = ~i_13_ & (~n609 | (~n453 & ~n610));
  assign n615 = ~i_32_ & n735;
  assign n616 = ~i_9_ & (n613 | (n614 & n615));
  assign n617 = n957 & (~n259 | ~n735 | n958);
  assign n618 = i_31_ | n610 | ~n615 | n958;
  assign n619 = n617 & (~i_29_ | (~n616 & n618));
  assign n620 = n974 & n515;
  assign n621 = n794 & n549;
  assign n622 = (~i_36_ | n621) & (n620 | ~n735);
  assign n623 = n433 | n413;
  assign n624 = (~n615 | n623) & (n473 | n622);
  assign n625 = n485 & n474;
  assign n626 = n472 & n484;
  assign n627 = (n473 | n625) & (~n308 | n626);
  assign n628 = n972 & n592;
  assign n629 = (n627 | n226) & (n628 | n172);
  assign n630 = n425 & ~n610;
  assign n631 = i_9_ | n610;
  assign n632 = n400 & n604;
  assign n633 = n631 | n632 | ~n214 | ~n421;
  assign n634 = ~i_21_ & n776;
  assign n635 = ~i_28_ & n219;
  assign n636 = n54 & n634 & (n630 | n635);
  assign n637 = ~n809 & (~n633 | (~i_28_ & ~n621));
  assign n638 = n310 & (~n898 | ~n907);
  assign n639 = n410 | n631 | i_19_ | ~n214;
  assign n640 = n114 | i_18_ | n608 | n501;
  assign n641 = ~n306 | ~n371;
  assign n642 = i_21_ | ~n655;
  assign n643 = n641 & (n523 | n642);
  assign n644 = ~n648 & (~n449 | ~n643);
  assign n645 = n371 & (~n504 | ~n521);
  assign n646 = n330 & (~n621 | (~i_32_ & ~n978));
  assign n647 = n352 | n651 | n438;
  assign n648 = n796 & n548;
  assign n649 = ~n646 & n647 & (n514 | n648);
  assign n650 = n978 | n204 | ~n310;
  assign n651 = n790 & n801;
  assign n652 = n650 & (~n306 | n438 | n651);
  assign n653 = (i_7_ | ~n259) & (n204 | n621);
  assign n654 = ~i_35_ & ~i_32_ & i_34_;
  assign n655 = ~i_23_ & ~i_24_;
  assign n656 = n655 & ~n226 & n654;
  assign n657 = ~n511 & (~n430 | ~n907);
  assign n658 = ~n451 & (~n506 | ~n521);
  assign n659 = ~i_29_ & n235;
  assign n660 = ~i_28_ & (n656 | (~n653 & n659));
  assign n661 = n306 & (n645 | (~n623 & n654));
  assign n662 = ~i_32_ & (n644 | (~i_7_ & ~n812));
  assign n663 = n50 & (n636 | n637 | n638);
  assign n664 = ~i_33_ | n777;
  assign n665 = (~n235 | n664) & (~n229 | n510);
  assign n666 = n973 & n900;
  assign n667 = n411 & (i_31_ | n666);
  assign n668 = n951 & (n678 | n172 | n510);
  assign n669 = (~n330 | n620) & (n514 | n947);
  assign n670 = n668 & n669 & (n667 | n352);
  assign n671 = n140 & (i_31_ | ~n421 | n610);
  assign n672 = ~i_8_ & ~n812;
  assign n673 = ~n751 & n306 & ~n628;
  assign n674 = ~i_31_ & (n672 | (~n643 & ~n980));
  assign n675 = n50 & (~n950 | (n300 & ~n411));
  assign n676 = ~n371 | i_31_ | n62 | n777 | n787;
  assign n677 = n676 & (~n537 | n631 | ~n813);
  assign n678 = n423 & n556;
  assign n679 = n678 | ~n50 | n167;
  assign n680 = ~n226 & ~i_34_ & n128;
  assign n681 = ~i_14_ & ~i_25_;
  assign n682 = i_28_ | i_30_ | n394 | n681;
  assign n683 = ~n421 | i_24_ | ~n259;
  assign n684 = n379 & ~n544;
  assign n685 = n683 & (~i_29_ | n510 | n684);
  assign n686 = n655 & i_21_;
  assign n687 = n686 & (~n682 | (~n571 & ~n807));
  assign n688 = (n222 | n510) & (~n50 | n769);
  assign n689 = n688 & (n201 | ~n306);
  assign n690 = i_23_ | n777;
  assign n691 = (n450 | n218) & (n690 | n201);
  assign n692 = n779 | ~i_21_ | n691;
  assign n693 = n692 & (n689 | n438);
  assign n694 = i_11_ | n806;
  assign n695 = ~i_3_ | n806;
  assign n696 = (i_18_ | n695) & (i_19_ | n694);
  assign n697 = i_21_ & ~i_23_;
  assign n698 = n697 & i_25_ & ~n664;
  assign n699 = i_22_ & n259 & n421;
  assign n700 = ~n379 & (n698 | (n530 & n531));
  assign n701 = n608 | i_18_ | n98;
  assign n702 = n701 & (i_7_ | ~n55 | n631);
  assign n703 = i_9_ | ~i_2_ | ~i_3_;
  assign n704 = n703 & (n100 | n608 | ~n735);
  assign n705 = ~n611 & ~i_9_ & n55;
  assign n706 = n421 & (n705 | (~i_18_ & ~n704));
  assign n707 = ~n706 & (~i_36_ | ~n425 | n702);
  assign n708 = ~n981 & (i_31_ | n288 | ~n546);
  assign n709 = ~n371 | n778;
  assign n710 = n709 & (~n537 | n610);
  assign n711 = n523 | n187 | n473;
  assign n712 = n711 & (~n51 | n204 | n288);
  assign n713 = ~n219 | ~i_34_ | ~i_36_;
  assign n714 = (~n330 | n713) & (~i_36_ | n712);
  assign n715 = ~n615 | i_2_ | n140;
  assign n716 = ~n983 & (~n52 | ~n214 | n438);
  assign n717 = (i_7_ | n714) & (n809 | ~n940);
  assign n718 = n970 & (~i_21_ | n691 | n729);
  assign n719 = n716 & (i_16_ | (n717 & n718));
  assign n720 = (n431 | n695) & (n432 | n694);
  assign n721 = ~n697 | n573 | n696;
  assign n722 = n721 & (n574 | n720);
  assign n723 = (i_17_ | n205) & (i_16_ | ~n307);
  assign n724 = n394 | n585;
  assign n725 = ~n332 & n724 & (~i_21_ | n584);
  assign n726 = i_31_ | i_30_ | n627 | n808;
  assign n727 = n726 & (~n54 | ~n308 | n713);
  assign n728 = (~n371 | n571) & (~i_31_ | n449);
  assign n729 = i_12_ | n805;
  assign n730 = (n689 | n729) & (~n52 | n441);
  assign n731 = ~i_21_ & (~n982 | (i_20_ & ~n708));
  assign n732 = n235 & (n699 | n700 | ~n943);
  assign n733 = i_34_ & (~n396 | n687 | ~n946);
  assign n734 = n615 & (~n679 | n680 | ~n948);
  assign n735 = ~i_35_ & i_36_;
  assign n736 = n735 & (n673 | n674 | n675);
  assign n737 = i_12_ | n581;
  assign n738 = i_21_ | i_22_;
  assign n739 = ~i_16_ & ~i_27_;
  assign n740 = i_23_ | i_17_;
  assign n741 = i_2_ | i_4_;
  assign n742 = ~i_9_ | n315;
  assign n743 = i_28_ | i_26_;
  assign n744 = i_8_ | ~i_9_;
  assign n745 = i_8_ | n315;
  assign n746 = i_2_ | i_3_;
  assign n747 = i_33_ | ~n219;
  assign n748 = ~i_9_ | n746;
  assign n749 = i_33_ | i_32_;
  assign n750 = i_31_ | n749;
  assign n751 = ~i_34_ | n541;
  assign n752 = i_30_ | i_29_;
  assign n753 = i_8_ | n314;
  assign n754 = i_4_ | n746;
  assign n755 = i_29_ | ~i_34_;
  assign n756 = ~i_9_ | ~n58;
  assign n757 = ~i_3_ | n741;
  assign n758 = n757 | n468;
  assign n759 = i_9_ | n758;
  assign n760 = n313 | n114;
  assign n761 = ~i_10_ | i_3_ | i_7_;
  assign n762 = i_35_ | i_33_ | ~i_34_;
  assign n763 = i_9_ | i_6_;
  assign n764 = n745 | n757;
  assign n765 = i_11_ | n763;
  assign n766 = i_7_ | n314;
  assign n767 = ~n51 | ~n655;
  assign n768 = ~n324 | n752;
  assign n769 = i_28_ | ~i_31_;
  assign n770 = n187 | i_7_ | i_28_;
  assign n771 = i_8_ | n746;
  assign n772 = i_22_ | ~n421 | n684 | ~n697;
  assign n773 = n754 | i_12_ | n742;
  assign n774 = ~i_38_ | i_2_ | i_7_;
  assign n775 = n61 | n62;
  assign n776 = ~i_16_ & ~i_23_;
  assign n777 = i_27_ | i_28_;
  assign n778 = i_30_ | n777;
  assign n779 = i_16_ | i_17_;
  assign n780 = i_0_ | i_4_;
  assign n781 = ~n537 | i_17_ | i_20_;
  assign n782 = i_18_ | n781;
  assign n783 = i_19_ | n779;
  assign n784 = i_12_ | n580;
  assign n785 = n313 | n766;
  assign n786 = i_18_ | n740;
  assign n787 = n315 | n316;
  assign n788 = i_5_ | n780;
  assign n789 = n114 | n788;
  assign n790 = n90 | ~i_13_ | i_14_;
  assign n791 = n313 | n753;
  assign n792 = i_23_ | n581;
  assign n793 = ~i_13_ | n763;
  assign n794 = n112 | n485;
  assign n795 = n84 | n361;
  assign n796 = n112 | n361;
  assign n797 = ~i_23_ & ~i_27_;
  assign n798 = ~i_25_ | n777;
  assign n799 = ~i_20_ | ~n655;
  assign n800 = i_20_ | ~n655;
  assign n801 = n90 | i_13_ | i_10_;
  assign n802 = n87 | n400;
  assign n803 = i_14_ | i_12_;
  assign n804 = n545 | n547 | n539 | ~n542;
  assign n805 = ~i_7_ | i_9_;
  assign n806 = ~i_7_ | ~i_10_;
  assign n807 = n605 | n806;
  assign n808 = ~i_34_ | ~n735;
  assign n809 = i_21_ | n740;
  assign n810 = i_23_ | ~i_20_ | i_21_;
  assign n811 = i_21_ | n779;
  assign n812 = i_2_ | n62 | n709 | n811;
  assign n813 = (i_13_ & ~i_14_) | (~i_10_ & (~i_13_ | ~i_14_));
  assign n814 = (n104 | n172) & (n167 | n318);
  assign n815 = (~n271 | n751) & (n190 | n750);
  assign n816 = (~n53 | n92) & (n67 | n240);
  assign n817 = (n84 | n756) & (~n58 | n83);
  assign n818 = n297 | ~i_19_ | n161;
  assign n819 = n818 & (i_28_ | n295 | n193);
  assign n820 = ~n322 & (n194 | (n190 & ~n303));
  assign n821 = ~n321 & (~n128 | n184 | n476);
  assign n822 = (~n51 | n319) & (n104 | n320);
  assign n823 = n791 & n84;
  assign n824 = (n148 | ~n303) & (n168 | n823);
  assign n825 = ~n323 & n824 & (n97 | n298);
  assign n826 = n659 & (~n115 | n285);
  assign n827 = (~n265 | n755) & (n135 | n743);
  assign n828 = ~n290 & (n111 | n167 | ~n654);
  assign n829 = n107 | n135;
  assign n830 = (~n128 | n224) & (~n265 | n509);
  assign n831 = n476 | i_28_ | ~n214;
  assign n832 = n831 & (i_7_ | ~n300 | n747);
  assign n833 = ~n271 & n297;
  assign n834 = (n88 | n225) & (n833 | n255);
  assign n835 = n111 | n161 | n167 | n117;
  assign n836 = n835 & (i_25_ | i_28_ | ~n826);
  assign n837 = n836 & (~i_35_ | n89 | n293);
  assign n838 = ~n301 & n837 & (n226 | n294);
  assign n839 = ~n302 & ~n304 & (n138 | n232);
  assign n840 = ~n305 & n839 & (n231 | n289);
  assign n841 = ~n336 | i_30_ | ~n271;
  assign n842 = n841 & (~n65 | n297);
  assign n843 = (~n60 | ~n310) & (i_24_ | n770);
  assign n844 = (n255 | ~n267) & (~n51 | ~n336);
  assign n845 = ~n276 & (~n278 | (n843 & n844));
  assign n846 = i_13_ | i_24_;
  assign n847 = (n192 | n147) & (n188 | n846);
  assign n848 = ~n251 & (n137 | ~n237 | n771);
  assign n849 = n77 | i_2_ | ~n59;
  assign n850 = n849 & (i_13_ | i_3_ | n195);
  assign n851 = ~n214 | n144 | n183;
  assign n852 = ~n254 & n851 & (~i_12_ | n250);
  assign n853 = (i_26_ | ~n66) & (~n659 | ~n775);
  assign n854 = n160 | n151 | n225;
  assign n855 = n854 & (i_28_ | n227 | n132);
  assign n856 = (n223 | n739) & (~i_23_ | ~n303);
  assign n857 = ~n217 & (n79 | ~n252 | ~n253);
  assign n858 = n188 | ~i_18_ | i_24_;
  assign n859 = n858 & (n192 | n146);
  assign n860 = (n202 | ~n300) & (n161 | n769);
  assign n861 = ~n72 & ~n74 & (~i_9_ | n70);
  assign n862 = (n68 | n149) & (~n237 | n773);
  assign n863 = n793 & n362;
  assign n864 = (n89 | n166) & (n863 | n173);
  assign n865 = (n148 | ~n324) & (n145 | ~n328);
  assign n866 = n106 | i_31_ | n875;
  assign n867 = i_2_ | i_8_ | n140 | ~n324;
  assign n868 = n536 | ~i_34_ | ~n421;
  assign n869 = n868 & (n97 | ~n121 | ~n324);
  assign n870 = n150 | n108 | n113;
  assign n871 = n870 & (~i_13_ | n105 | n313);
  assign n872 = n136 | i_2_ | n750;
  assign n873 = ~n122 & n872 & (n104 | n120);
  assign n874 = i_2_ | i_8_ | i_31_ | ~n269;
  assign n875 = n787 & n69;
  assign n876 = n874 & (~n324 | n750 | n875);
  assign n877 = ~n328 | i_10_ | n85;
  assign n878 = n877 & (~i_29_ | (~n775 & n776));
  assign n879 = (n82 | n282) & (n747 | n774);
  assign n880 = n879 & (n91 | ~n278);
  assign n881 = n536 | ~n235 | ~n421;
  assign n882 = n881 & (~n71 | n77 | n748);
  assign n883 = n882 & (~i_9_ | ~i_12_ | n79);
  assign n884 = ~n127 & ~n129 & (n126 | ~n280);
  assign n885 = ~n342 | n108 | n149;
  assign n886 = n885 & (n145 | n833 | n160);
  assign n887 = n142 | i_35_ | n185;
  assign n888 = ~n331 & (~i_38_ | (n838 & n840));
  assign n889 = n976 & n945 & n845 & n275 & ~n273 & ~n270 & n264 & ~n266;
  assign n890 = (~i_34_ | n889) & (i_29_ | n277);
  assign n891 = ~n334 & ~n337 & (~n50 | n772);
  assign n892 = (n133 | n241) & (n137 | n245);
  assign n893 = ~n338 & (i_24_ | (n855 & n856));
  assign n894 = ~n341 & (n200 | (n861 & n862));
  assign n895 = ~n343 & n894 & (n195 | n756);
  assign n896 = (n141 | n244) & (n159 | n190);
  assign n897 = n208 & (i_22_ | (n884 & n883));
  assign n898 = n785 | n440;
  assign n899 = ~n357 & (~n974 | (~n81 & ~n382));
  assign n900 = n791 | n792;
  assign n901 = n274 | n203 | ~n235;
  assign n902 = n901 & (~i_20_ | n573 | ~n776);
  assign n903 = n752 | ~i_31_ | n567;
  assign n904 = n903 & (n506 | n292 | n566);
  assign n905 = n767 | i_7_ | n750;
  assign n906 = ~n529 & (~n229 | n798 | n799);
  assign n907 = n785 | n792;
  assign n908 = n295 | n438 | n510 | n801;
  assign n909 = ~n214 | i_0_ | i_30_ | n800 | n380 | n523;
  assign n910 = n441 | n354 | n792;
  assign n911 = n910 & (n357 | n486);
  assign n912 = ~n259 | i_7_ | i_23_ | ~n267 | n351;
  assign n913 = (~n427 | n795) & (n397 | n507);
  assign n914 = n438 | n801 | ~i_37_ | ~n299;
  assign n915 = n914 & (n318 | ~n427 | n477);
  assign n916 = n62 | ~i_2_ | i_16_;
  assign n917 = n916 & (n401 | n100 | n788);
  assign n918 = n404 | n412 | ~i_37_ | n98;
  assign n919 = (n297 | n555) & (~n300 | n408);
  assign n920 = i_30_ | ~i_31_ | ~n306 | n379;
  assign n921 = n920 & (i_14_ | n495 | n369);
  assign n922 = n488 | n315 | n377 | n495 | ~n537;
  assign n923 = n922 & (n363 | ~n427 | n641);
  assign n924 = n450 | n508 | n297;
  assign n925 = n751 | ~n546 | ~n686;
  assign n926 = n925 & (n354 | n438 | n790);
  assign n927 = n495 | i_13_ | n491;
  assign n928 = (n434 | n570) & (~i_7_ | n582);
  assign n929 = n548 | n224 | n353;
  assign n930 = (n204 | n563) & (~n427 | n560);
  assign n931 = (n684 | n534) & (n553 | n351);
  assign n932 = (~i_37_ | n522) & (~n259 | n499);
  assign n933 = (i_14_ | n461) & (n481 | n523);
  assign n934 = n977 & n772 & ~n428 & ~n426 & ~n422 & n424;
  assign n935 = (~n50 | n934) & (~n306 | n448);
  assign n936 = (~i_34_ | n396) & (i_32_ | n390);
  assign n937 = n752 | ~i_34_ | n510;
  assign n938 = n937 & (i_30_ | ~n235 | ~n306);
  assign n939 = (n379 | n395) & (~n307 | ~n308);
  assign n940 = n50 & (~n715 | (i_0_ & n421));
  assign n941 = n274 | ~n544 | n696 | ~n797;
  assign n942 = n941 & (~n527 | n769 | n807);
  assign n943 = n942 & (~n391 | n684 | n810);
  assign n944 = n807 | n274 | n450;
  assign n945 = n767 | ~i_14_ | n394;
  assign n946 = n944 & n945 & (n685 | n810);
  assign n947 = n360 & n436;
  assign n948 = (n947 | n641) & (n677 | n811);
  assign n949 = n671 | n626 | ~n634;
  assign n950 = n949 & (n666 | n167);
  assign n951 = n450 | n980 | n167;
  assign n952 = n537 & (~n639 | ~n640);
  assign n953 = n203 | n288 | ~n51 | ~n54;
  assign n954 = n953 & (i_17_ | i_21_ | ~n952);
  assign n955 = n954 & (i_7_ | n751 | n767);
  assign n956 = (~n235 | n652) & (~i_34_ | n649);
  assign n957 = n232 | n606 | i_30_ | ~i_36_;
  assign n958 = n737 & n784;
  assign n959 = ~i_36_ | ~n54 | n187 | ~n308;
  assign n960 = n479 & n959 & (n629 | ~n735);
  assign n961 = (n619 | n642) & (i_29_ | n624);
  assign n962 = n723 | n665 | ~n697;
  assign n963 = n962 & (n730 | (n440 & n792));
  assign n964 = n963 & (n728 | n807);
  assign n965 = (n681 | n725) & (~n306 | n727);
  assign n966 = (~n544 | n722) & (n62 | n719);
  assign n967 = (~i_36_ | ~n979) & (n670 | n808);
  assign n968 = n967 & (n523 | (n961 & n960));
  assign n969 = n515 | i_29_ | n473 | n397;
  assign n970 = n441 | n710 | i_21_ | ~i_36_;
  assign n971 = i_33_ | n743;
  assign n972 = ~n308 | i_13_ | n69;
  assign n973 = n440 | n791;
  assign n974 = n81 | n604;
  assign n975 = ~n278 | n175 | n233;
  assign n976 = n260 | i_24_ | i_28_;
  assign n977 = i_0_ | n398 | n405 | ~n635;
  assign n978 = n381 & n802;
  assign n979 = n660 | n661 | n657 | n658 | ~n955 | ~n956 | n662 | n663;
  assign n980 = n507 & n795;
  assign n981 = n526 & ~n161 & n259;
  assign n982 = n413 | n707 | i_23_ | ~n50;
  assign n983 = n634 & n421 & n50 & i_0_ & ~i_12_;
endmodule


