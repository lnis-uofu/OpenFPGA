// Benchmark "TOP" written by ABC on Mon Feb  4 17:34:12 2019

module spla ( 
    i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_,
    i_11_, i_12_, i_13_, i_14_, i_15_,
    o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_,
    o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_,
    o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_,
    o_31_, o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_, o_40_,
    o_41_, o_42_, o_43_, o_44_, o_45_  );
  input  i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_,
    i_10_, i_11_, i_12_, i_13_, i_14_, i_15_;
  output o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_,
    o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_,
    o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_,
    o_31_, o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_, o_40_,
    o_41_, o_42_, o_43_, o_44_, o_45_;
  wire n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
    n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
    n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
    n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
    n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
    n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
    n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
    n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
    n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
    n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
    n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
    n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
    n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
    n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
    n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
    n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
    n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
    n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
    n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
    n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
    n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
    n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
    n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
    n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
    n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
    n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
    n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
    n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
    n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
    n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
    n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
    n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
    n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
    n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
    n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
    n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
    n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
    n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
    n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
    n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
    n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
    n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
    n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
    n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
    n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
    n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
    n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
    n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
    n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
    n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
    n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
    n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
    n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
    n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
    n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
    n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
    n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
    n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
    n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
    n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
    n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
    n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
    n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
    n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
    n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
    n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
    n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
    n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
    n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
    n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
    n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
    n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
    n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
    n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
    n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
    n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
    n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
    n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
    n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
    n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
    n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
    n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
    n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
    n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
    n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
    n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
    n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
    n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
    n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
    n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
    n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
    n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
    n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
    n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
    n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
    n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
    n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
    n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
    n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
    n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
    n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
    n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
    n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
    n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
    n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
    n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
    n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
    n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
    n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
    n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
    n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
    n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
    n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
    n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
    n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
    n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
    n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
    n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
    n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
    n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
    n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
    n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
    n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
    n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
    n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
    n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
    n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
    n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
    n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
    n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
    n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
    n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
    n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
    n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
    n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
    n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
    n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
    n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
    n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
    n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
    n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
    n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
    n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
    n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
    n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
    n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
    n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
    n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
    n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
    n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
    n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
    n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
    n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
    n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
    n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
    n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
    n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
    n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
    n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
    n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
    n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
    n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
    n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
    n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
    n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
    n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
    n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
    n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
    n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
    n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
    n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
    n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
    n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
    n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
    n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
    n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
    n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
    n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
    n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
    n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
    n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
    n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
    n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
    n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
    n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
    n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
    n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
    n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
    n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
    n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
    n2296, n2297, n2298;
  assign o_0_ = ~n211;
  assign o_1_ = ~n125;
  assign o_2_ = n184 & ~n1084 & (~n984 | ~n1074);
  assign o_3_ = ~n210;
  assign o_4_ = ~n206;
  assign o_5_ = ~n566;
  assign o_6_ = ~n205;
  assign o_7_ = ~n514;
  assign o_8_ = i_3_ & ~i_0_ & ~i_1_;
  assign o_9_ = ~n203;
  assign o_10_ = ~n202;
  assign o_11_ = ~n201;
  assign o_12_ = ~n1064;
  assign o_13_ = ~n200;
  assign o_14_ = ~n1032;
  assign o_15_ = ~n1024;
  assign o_16_ = ~n195;
  assign o_17_ = ~n1017;
  assign o_18_ = ~n186;
  assign o_19_ = n184 & i_5_ & i_3_ & ~i_4_ & ~n1074;
  assign o_20_ = ~n1074 & n184 & n185;
  assign o_21_ = n183 | n181 | n182;
  assign o_22_ = ~n180;
  assign o_23_ = ~n179;
  assign o_24_ = n172 & ~n1083;
  assign o_25_ = n172 & n173;
  assign o_26_ = n163 | n167 | n171 | n158;
  assign o_27_ = n162 | n168 | ~n174 | ~n2250;
  assign o_28_ = n167 | n168 | n169 | n170;
  assign o_29_ = n164 | n162 | n163 | ~n174 | n165 | n166;
  assign o_30_ = n161 | n159 | n160 | n158 | ~n156 | n157;
  assign o_31_ = n955 | n956 | ~n1605 | ~n2244;
  assign o_32_ = ~n954;
  assign o_33_ = ~n952;
  assign o_34_ = ~n156;
  assign o_35_ = ~n153;
  assign o_36_ = ~n937;
  assign o_37_ = ~n146;
  assign o_38_ = ~n873;
  assign o_39_ = ~n788;
  assign o_40_ = ~n145;
  assign o_41_ = n144 & n142 & n143;
  assign o_42_ = ~n141;
  assign o_43_ = ~n138;
  assign o_44_ = ~n134;
  assign o_45_ = ~n126;
  assign n108 = ~n469 & (~n497 | ~n1574);
  assign n109 = ~n349 & (~n484 | ~n1105);
  assign n110 = n555 & n1101;
  assign n111 = ~n781 | ~n1224;
  assign n112 = n110 & (n111 | ~n463);
  assign n113 = ~n796 & (~n845 | ~n849);
  assign n114 = n218 | ~n268;
  assign n115 = ~n405 & (n114 | ~n779);
  assign n116 = ~n225 & (~n377 | ~n636);
  assign n117 = n110 & (~n1105 | ~n1202);
  assign n118 = ~n1458 | ~n1468;
  assign n119 = ~n405 & (n118 | ~n1151 | ~n1231);
  assign n120 = n385 | ~n945;
  assign n121 = ~n796 & (n120 | ~n1005);
  assign n122 = n1084 | ~n1515;
  assign n123 = i_7_ | i_6_;
  assign n124 = n122 | n123;
  assign n125 = n983 & (~n144 | n984 | n985);
  assign n126 = n517 & n669 & (n667 | n670);
  assign n127 = n743 & n708 & n704 & n742 & n721 & n735 & n744 & n745;
  assign n128 = n1649 & n1648 & n1647 & n1645 & n1644 & n409 & ~n701 & n1646;
  assign n129 = n1655 & n1654 & n1653 & n1652 & n1650 & n1651 & n700;
  assign n130 = n1643 & n749 & n1642 & n1641 & n336 & n1640;
  assign n131 = n2160 & (n405 | (n1006 & n1547));
  assign n132 = n675 & n1677 & n698 & n1662 & n1669 & n1674 & n1684;
  assign n133 = n2159 & n2158 & n2157 & n2156 & n2155 & n195 & ~n115 & ~n119;
  assign n134 = n132 & n131 & n130 & n129 & n127 & n128 & n133 & ~n752;
  assign n135 = n1699 & n1698 & n1697 & n1696 & ~n767 & ~n765 & ~n217 & n757;
  assign n136 = ~n430 | n1115;
  assign n137 = ~n430 | n1200;
  assign n138 = n137 & n136 & n127 & n135;
  assign n139 = n196 & n240 & (n241 | n242);
  assign n140 = n197 & n480 & (n481 | n242);
  assign n141 = n139 & n140;
  assign n142 = ~i_11_ & ~i_9_ & ~i_10_;
  assign n143 = ~i_8_ & n1119;
  assign n144 = ~n1084 & n1700;
  assign n145 = n768 & n519 & (n769 | n568);
  assign n146 = n912 & n911 & n910 & n909 & n708 & n908 & n913 & n914;
  assign n147 = ~n948 & (n456 | (n747 & n944));
  assign n148 = n2239 & (n943 | n755);
  assign n149 = n2241 & n2242 & (n746 | n405);
  assign n150 = n1359 & n1322 & n307 & n1488 & n367 & n420;
  assign n151 = n1611 & n585 & n649 & n1779 & n807 & n1761;
  assign n152 = n2238 & n2237 & n1909 & n1896 & n1857 & n1258 & ~n121 & ~n947;
  assign n153 = ~n950 & n152 & n151 & n150 & n149 & n147 & n148 & ~n949;
  assign n154 = n1080 & n1079 & n1078 & n1077 & n1075 & n1076 & n1081 & n1082;
  assign n155 = n663 & n661;
  assign n156 = n154 & n155;
  assign n157 = ~n525 & ~n1787;
  assign n158 = n963 | n964 | n965 | n966 | ~n2246 | n967 | n968;
  assign n159 = n957 | n958 | n959 | n960 | ~n2247 | n961 | n962;
  assign n160 = ~n516 & ~n525;
  assign n161 = ~n525 & n1529;
  assign n162 = n1521 | n1785 | n1786;
  assign n163 = n1522 | n971 | n1783 | n1531;
  assign n164 = ~n516 & ~n1214;
  assign n165 = ~n1214 & n1529;
  assign n166 = ~n1214 & ~n1787;
  assign n167 = n1703 | n1784 | n1788 | n1789 | ~n124 | n978 | n1523 | n1532;
  assign n168 = n972 | n973 | n974 | n975 | ~n2248 | n976 | n977;
  assign n169 = ~n515 & n1529;
  assign n170 = ~n515 & (~n516 | ~n1787);
  assign n171 = ~n2249 & n185 & ~n1512;
  assign n172 = ~n1512 & (n185 | n222);
  assign n173 = ~i_6_ & i_7_;
  assign n174 = n518 & (n969 | n970);
  assign n175 = n774 & (n304 | n516);
  assign n176 = n522 & (n516 | (n523 & n524));
  assign n177 = ~n1525 & ~n1534;
  assign n178 = n122 & ~n958;
  assign n179 = ~n1704 & ~n980 & ~n183 & n178 & n177 & n176 & n174 & n175;
  assign n180 = n520 & n981 & (~n979 | n982);
  assign n181 = ~n665 & n555 & n556;
  assign n182 = ~n1117 & n556 & ~n665;
  assign n183 = n1784 | n1783 | n966 | n974 | n1785 | n959;
  assign n184 = ~n985 & n1700;
  assign n185 = ~i_5_ & i_3_ & i_4_;
  assign n186 = n1001 & n1000 & n999 & n998 & n875 & n997 & n1002 & n1003;
  assign n187 = n684 | n1354;
  assign n188 = n543 | n684;
  assign n189 = ~n120 | n684;
  assign n190 = n1262 | n684;
  assign n191 = n684 | n1309;
  assign n192 = n684 | n535;
  assign n193 = n684 | n1340;
  assign n194 = n686 & n1842 & n1305 & n1633 & n1621 & n908;
  assign n195 = n192 & n191 & n190 & n189 & n187 & n188 & n193 & n194;
  assign n196 = n1142 & n1140 & n1141;
  assign n197 = n1476 & n1475 & n1474 & n479;
  assign n198 = n603 & n602 & n600 & n601;
  assign n199 = n590 & n1747 & n604;
  assign n200 = n155 & n199 & n198 & n196 & n197;
  assign n201 = n209 & ~n1704 & (n770 | n771);
  assign n202 = n1071 & n1070 & n1069 & n1068 & n440 & n291 & n1072 & n1073;
  assign n203 = n392 & n391 & n390 & n389 & n387 & n388 & n393 & n394;
  assign n204 = n517 & n521 & n520 & n518 & n519;
  assign n205 = n204 & n122 & n176;
  assign n206 = ~n1536 & n177 & ~n1520;
  assign n207 = n176 & (n770 | n771);
  assign n208 = n122 & ~n1704;
  assign n209 = n981 & n768 & n777 & n774;
  assign n210 = n209 & n204 & n207 & n208;
  assign n211 = ~n1515 & (~n144 | n985 | n1074);
  assign n212 = n1099 & n1101;
  assign n213 = n212 & (~n1118 | ~n1136);
  assign n214 = ~n349 & (~n725 | ~n1634);
  assign n215 = ~n469 & (~n1208 | ~n1224);
  assign n216 = n1086 & n143;
  assign n217 = ~n1261 & (n216 | ~n755);
  assign n218 = ~n781 | ~n987;
  assign n219 = ~n225 & (n218 | ~n570);
  assign n220 = n1101 & n143;
  assign n221 = n220 & (~n781 | ~n1127);
  assign n222 = i_3_ & i_5_ & i_4_;
  assign n223 = n225 | n1111;
  assign n224 = n225 | n1110;
  assign n225 = ~n555 | ~n1093;
  assign n226 = n1090 | n1091;
  assign n227 = n223 & n224 & (n225 | n226);
  assign n228 = n1198 & n1204;
  assign n229 = n1118 & n237;
  assign n230 = n352 & n374;
  assign n231 = n1088 | n1095;
  assign n232 = n1095 | n1109;
  assign n233 = n824 & n235;
  assign n234 = n233 & n232 & n231 & n230 & n228 & n229;
  assign n235 = n1109 | n1167;
  assign n236 = n1109 | n1163;
  assign n237 = n1090 | n1109;
  assign n238 = n1103 | n1122;
  assign n239 = n238 & n237 & n236 & n235 & n232;
  assign n240 = n1747 & n2027 & (n2028 | n265);
  assign n241 = i_11_ | ~i_9_ | ~i_10_;
  assign n242 = n984 | ~n1138;
  assign n243 = n1074 | ~n1086;
  assign n244 = n1088 | n1104;
  assign n245 = n1104 | n1109;
  assign n246 = (n243 | n244) & (~n212 | n245);
  assign n247 = n419 & n456;
  assign n248 = ~n815 & ~n379 & n247 & ~n250;
  assign n249 = ~n1154 & (~n728 | ~n987);
  assign n250 = ~n349 | ~n796;
  assign n251 = ~n988 & (n250 | ~n488 | ~n1166);
  assign n252 = ~n249 & (n1164 | (n780 & n1129));
  assign n253 = ~n219 & (~n277 | (n1111 & n1151));
  assign n254 = ~n251 & n2040 & (n236 | n2012);
  assign n255 = n1538 & n588 & n471 & n890 & n1771 & n921 & n639 & n635;
  assign n256 = n2043 & n2044 & n2046 & n2045 & n658 & n246 & n2042 & n2041;
  assign n257 = n1721 & n848 & n837 & n790 & n455 & n410 & n467 & n631;
  assign n258 = n395 & n399 & n2039 & n627 & n641 & n462 & n1691 & n1690;
  assign n259 = n719 & n1625 & n404 & n408 & n1641 & n415 & n2035 & n2038;
  assign n260 = n257 & n256 & n255 & n254 & n252 & n253 & n258 & n259;
  assign n261 = n1120 | ~n1138;
  assign n262 = ~n142 | n261;
  assign n263 = n478 | n261;
  assign n264 = n1131 | n261;
  assign n265 = i_11_ | i_9_ | ~i_10_;
  assign n266 = n263 & n264 & (n265 | n261);
  assign n267 = n225 | n1217;
  assign n268 = n1226 & n1224 & n1225;
  assign n269 = n1126 | n1196;
  assign n270 = n267 & (n225 | (n268 & n269));
  assign n271 = n539 | ~n796;
  assign n272 = ~n1210 & (n271 | ~n488);
  assign n273 = n220 | ~n456;
  assign n274 = n273 & (~n824 | ~n1204 | ~n1232);
  assign n275 = ~n377 | ~n1307;
  assign n276 = ~n1154 & (~n268 | n275 | ~n1213);
  assign n277 = ~n243 | ~n405;
  assign n278 = ~n226 | ~n1353;
  assign n279 = n277 & (n278 | ~n1203 | ~n1231);
  assign n280 = ~n243 | n818;
  assign n281 = ~n488 | ~n349 | ~n456;
  assign n282 = ~n1200 & (n271 | n280 | n281);
  assign n283 = ~n274 & (n1197 | (n469 & n1157));
  assign n284 = ~n272 & (n2010 | (n643 & n1207));
  assign n285 = ~n276 & n2013 & (n1218 | n2014);
  assign n286 = n889 & n1078 & n920 & n915 & n1768 & n2009 & n587 & n638;
  assign n287 = n2020 & n2018 & n2017 & n2016 & ~n279 & ~n282;
  assign n288 = n789 & n411 & n451 & n454 & n458 & n634 & n836 & n847;
  assign n289 = n396 & n400 & n626 & n461 & n1722 & n630 & n1688 & n2008;
  assign n290 = n2007 & n1591 & n1586 & n1626 & n407 & n403 & n2003 & n2006;
  assign n291 = n288 & n287 & n286 & n285 & n283 & n284 & n289 & n290;
  assign n292 = n236 | ~n421;
  assign n293 = n456 | n1153;
  assign n294 = n232 | ~n818;
  assign n295 = n456 | n530;
  assign n296 = n456 | n1149;
  assign n297 = n236 | ~n925;
  assign n298 = n1579 & n1566 & n577 & n1726 & n1618 & n591;
  assign n299 = n1996 & n1995 & n1689 & n1630 & n1279 & n1267 & ~n217 & n655;
  assign n300 = n1989 & n1705 & n1716 & n1694 & n718 & n1990 & n1986 & n1982;
  assign n301 = n298 & n297 & n296 & n295 & n293 & n294 & n299 & n300;
  assign n302 = n405 & n419;
  assign n303 = n238 | n302;
  assign n304 = n1089 | n1113;
  assign n305 = n1089 | n1128;
  assign n306 = n304 & n305;
  assign n307 = n1306 & n303 & n1305 & n188 & n1303 & n1304;
  assign n308 = n1302 & n1301 & n1300 & n1299 & n1297 & n1298;
  assign n309 = n1294 & n1293 & n1292 & n1291 & n1289 & n1290 & n1295 & n1296;
  assign n310 = n1287 & n1286 & n1285 & n1284 & n1282 & n1283 & n1288;
  assign n311 = n1973 & n1974 & (~n216 | n238);
  assign n312 = n1751 & n1686 & n1631 & n1559 & n1772 & n1749 & n1710 & n1972;
  assign n313 = n1971 & n812 & n1752 & n1619 & n595 & n1583;
  assign n314 = n1968 & n1657 & n1970 & n1969 & n1678 & n1596;
  assign n315 = n312 & n311 & n310 & n309 & n307 & n308 & n313 & n314;
  assign n316 = n1091 | n1167;
  assign n317 = ~n220 | n316;
  assign n318 = n456 | n316;
  assign n319 = ~n818 | n824;
  assign n320 = n456 | n484;
  assign n321 = n456 | n1228;
  assign n322 = ~n925 | n1227;
  assign n323 = n1584 & n594 & n580 & n1565 & n1715;
  assign n324 = n1330 & n1337 & n1953 & n1713 & n1767 & n1955 & n1954 & n1322;
  assign n325 = n1950 & n786 & n785 & n1706 & n1951 & n1952 & n1949;
  assign n326 = n323 & n322 & n321 & n320 & n318 & n319 & n324 & n325;
  assign n327 = n1352 & n1351 & n1350 & n1349 & n1347 & n1348;
  assign n328 = n1346 & n1345 & n1344 & n1343 & n1341 & n1342;
  assign n329 = n1934 & (~n818 | n970);
  assign n330 = (n419 | n726) & (~n216 | n1232);
  assign n331 = n1933 & (n243 | n1045);
  assign n332 = n1931 & n1632 & n1711 & n1628 & n1687 & n1932;
  assign n333 = n596 & n1753 & n1545 & n811 & n1620 & n1616 & n582 & n1930;
  assign n334 = n1928 & n1654 & n1672 & n1663 & n693 & n1656;
  assign n335 = n332 & n331 & n330 & n329 & n327 & n328 & n333 & n334;
  assign n336 = n243 | n1212;
  assign n337 = n243 | n1097;
  assign n338 = n1110 | n405;
  assign n339 = n243 | n1225;
  assign n340 = n243 | n1135;
  assign n341 = n717 & n1595 & n1594 & n1610 & n1682 & n1681;
  assign n342 = n1915 & n1575 & n579 & n1568 & n1567 & n1671 & n1651 & n1914;
  assign n343 = n1359 & n1368 & n1919 & n1627 & n1922 & n1561 & n1921 & n1918;
  assign n344 = n341 & n340 & n339 & n338 & n336 & n337 & n342 & n343;
  assign n345 = n1088 | n1102;
  assign n346 = n1102 | n1109;
  assign n347 = ~n892 & n345 & n346;
  assign n348 = n1214 & n780;
  assign n349 = ~n555 | ~n1086;
  assign n350 = (n348 | n349) & (n347 | ~n430);
  assign n351 = n349 | n1127;
  assign n352 = n1208 & n1127;
  assign n353 = n643 & n1129;
  assign n354 = n351 & (~n430 | (n352 & n353));
  assign n355 = ~n879 & n1136;
  assign n356 = n355 | ~n421;
  assign n357 = n225 | n1339;
  assign n358 = n405 | n1340;
  assign n359 = n349 | n1339;
  assign n360 = n349 | n726;
  assign n361 = n225 | n1232;
  assign n362 = n469 | n1339;
  assign n363 = n1161 | n1340;
  assign n364 = n1846 & n1843 & n1845 & n1844 & n193 & n1697;
  assign n365 = n362 & n361 & n360 & n359 & n357 & n358 & n363 & n364;
  assign n366 = (~n385 | n419) & (n225 | n995);
  assign n367 = n366 & n365;
  assign n368 = ~n984 & n1101;
  assign n369 = n368 & (~n1232 | ~n1340);
  assign n370 = ~n110 | n780;
  assign n371 = n2298 | n225;
  assign n372 = ~n879 & n1215;
  assign n373 = n370 & n371 & (~n110 | n372);
  assign n374 = n345 & n346;
  assign n375 = n1394 & ~n385 & n1280;
  assign n376 = n375 & n374 & n231;
  assign n377 = n515 & n1215;
  assign n378 = n377 & ~n892;
  assign n379 = ~n243 | n368;
  assign n380 = n379 & (~n233 | ~n374);
  assign n381 = n212 | n110;
  assign n382 = ~n346 | ~n1281;
  assign n383 = n381 & (n382 | n111);
  assign n384 = n277 & (~n990 | ~n1133);
  assign n385 = ~n1261 | ~n1308;
  assign n386 = n368 & (n385 | ~n648);
  assign n387 = (~n250 | ~n275) & (n243 | n1606);
  assign n388 = (~n385 | n684) & (n302 | n652);
  assign n389 = (n352 | n405) & (n355 | n796);
  assign n390 = (n1152 | n738) & (n1781 | n1161);
  assign n391 = n2069 & n2070 & n373 & n1076 & n418 & n367;
  assign n392 = n291 & n260 & n335 & n326 & n301 & n315 & n227 & n2071;
  assign n393 = n2058 & n2060 & n2062 & n2065 & n2067 & n2068 & n2056 & n2055;
  assign n394 = n2054 & n2053 & n2051 & n2050 & n2049 & n2048 & ~n213 & n2047;
  assign n395 = n225 | n1123;
  assign n396 = n225 | n231;
  assign n397 = n1089 | n1095;
  assign n398 = n395 & n396 & (n225 | n397);
  assign n399 = n225 | n1124;
  assign n400 = n225 | n1204;
  assign n401 = n1089 | n1090;
  assign n402 = n399 & n400 & (n225 | n401);
  assign n403 = n405 | n231;
  assign n404 = n405 | n232;
  assign n405 = ~n1086 | n1117;
  assign n406 = n403 & n404 & (n405 | n397);
  assign n407 = n405 | n1204;
  assign n408 = n405 | n237;
  assign n409 = n407 & n408 & (n405 | n401);
  assign n410 = n225 | n1136;
  assign n411 = n225 | n1198;
  assign n412 = n1089 | n1106;
  assign n413 = n410 & n411 & (n225 | n412);
  assign n414 = n405 | n1198;
  assign n415 = n405 | n1118;
  assign n416 = n414 & n415 & (n405 | n412);
  assign n417 = n349 | n1261;
  assign n418 = n1406 & n190 & n1405 & n1019 & n1403 & n1404;
  assign n419 = ~n1093 | n1117;
  assign n420 = n417 & n418 & (n419 | n235);
  assign n421 = ~n349 | n430;
  assign n422 = ~n1136 & (n421 | ~n796);
  assign n423 = n1431 & n1430 & n1429 & n1428 & n1426 & n1427 & n1432 & n1433;
  assign n424 = n1377 & n2090 & (~n539 | n1124);
  assign n425 = (~n815 | n1149) & (n243 | n1153);
  assign n426 = (n2088 | n1261) & (n1461 | n346);
  assign n427 = n2089 & (n235 | (~n539 & n1461));
  assign n428 = ~n422 & (n1127 | (~n421 & n1459));
  assign n429 = n426 & n425 & n424 & n420 & n301 & n423 & n427 & n428;
  assign n430 = n1086 & n1099;
  assign n431 = ~n1208 & (n430 | ~n1459);
  assign n432 = n469 | n1307;
  assign n433 = n469 | n1219;
  assign n434 = ~n431 & (n824 | (n1461 & n1462));
  assign n435 = (~n546 | n1309) & (n231 | n2087);
  assign n436 = n1517 | n1307;
  assign n437 = (n1461 | n345) & (n1463 | n1219);
  assign n438 = (n2088 | n1308) & (n2066 | n1228);
  assign n439 = n326 & n1075 & (~n212 | n1224);
  assign n440 = n437 & n436 & n435 & n434 & n432 & n433 & n438 & n439;
  assign n441 = n368 & (~n636 | ~n1467);
  assign n442 = n469 | n632;
  assign n443 = n469 | n1465;
  assign n444 = n469 | n628;
  assign n445 = ~n110 | n632;
  assign n446 = n2085 & (~n212 | (n463 & n632));
  assign n447 = (~n381 | n642) & (n684 | n1467);
  assign n448 = n1473 & n1472 & n1471 & n1470 & ~n441 & n1469;
  assign n449 = n2086 & (~n679 | n1481);
  assign n450 = n447 & n446 & n445 & n444 & n442 & n443 & n448 & n449;
  assign n451 = ~n220 | n231;
  assign n452 = n397 & n232;
  assign n453 = n451 & (~n220 | n452);
  assign n454 = n456 | n1198;
  assign n455 = n1118 | n456;
  assign n456 = ~n1101 | n1120;
  assign n457 = n454 & n455 & (n456 | n412);
  assign n458 = ~n220 | n1198;
  assign n459 = n412 & n1118;
  assign n460 = n458 & (~n220 | n459);
  assign n461 = n456 | n1208;
  assign n462 = n456 | n1127;
  assign n463 = n1089 | n1126;
  assign n464 = n461 & n462 & (n456 | n463);
  assign n465 = ~n233 | ~n482;
  assign n466 = n220 & (n465 | ~n486);
  assign n467 = n469 | n1123;
  assign n468 = n469 | n231;
  assign n469 = ~n1101 | n1114;
  assign n470 = n467 & n468 & (n469 | n397);
  assign n471 = n469 | n1136;
  assign n472 = n469 | n1198;
  assign n473 = n471 & n472 & (n469 | n412);
  assign n474 = n2076 & (~n1053 | (n945 & n1048));
  assign n475 = ~n368 | n725;
  assign n476 = n475 & n474 & n470 & n473;
  assign n477 = ~n1099 | ~n1138;
  assign n478 = ~i_11_ | i_9_ | i_10_;
  assign n479 = n477 | n478;
  assign n480 = n2075 & (n2028 | n478);
  assign n481 = ~i_11_ | ~i_9_ | i_10_;
  assign n482 = n1089 | n1167;
  assign n483 = n482 | n349;
  assign n484 = n1091 | n1102;
  assign n485 = n1481 & n1480 & n589 & n1465 & n1467;
  assign n486 = n1108 | n1167;
  assign n487 = n486 & n485 & n484 & n226 & n316;
  assign n488 = n225 & n302;
  assign n489 = ~n421 & ~n818;
  assign n490 = ~n1051 & n488 & n489;
  assign n491 = n1090 | n1108;
  assign n492 = n482 & n401 & n491 & n486;
  assign n493 = ~n212 | n2293;
  assign n494 = n493 & (~n212 | n491);
  assign n495 = n1108 | n1126;
  assign n496 = n1108 | n1163;
  assign n497 = n1102 | n1108;
  assign n498 = n497 & n495 & n496;
  assign n499 = n381 & (~n346 | ~n495);
  assign n500 = ~n796 & (~n397 | ~n530);
  assign n501 = ~n419 | ~n850;
  assign n502 = n501 & (~n1123 | ~n1136 | ~n1458);
  assign n503 = n501 | ~n1154;
  assign n504 = n503 & (~n530 | ~n1219 | ~n1307);
  assign n505 = ~n488 & (~n463 | ~n482 | ~n781);
  assign n506 = (n397 | n1460) & (~n277 | n1458);
  assign n507 = (n1157 | n487) & (n1155 | n482);
  assign n508 = (n1483 | n496) & (n1807 | n530);
  assign n509 = (n2099 | n1479) & (n2011 | n725);
  assign n510 = n2098 & n2097 & n2095 & ~n505 & ~n502 & ~n504;
  assign n511 = n2093 & n2094 & n1708 & n896 & n1560 & n1540;
  assign n512 = n1617 & n1624 & n1629 & n1647 & n844 & n1707 & n2091 & n1587;
  assign n513 = n2104 & n2106 & n2108 & n2112 & n2110 & n2109 & n2114 & n2113;
  assign n514 = n511 & n510 & n509 & n508 & n506 & n507 & n512 & n513;
  assign n515 = n1106 | n1201;
  assign n516 = ~n1099 | n1513;
  assign n517 = ~n160 & ~n164 & (n515 | n516);
  assign n518 = n970 | n516;
  assign n519 = n1514 | n985;
  assign n520 = n1514 | n665;
  assign n521 = (n1514 | n776) & (n304 | n516);
  assign n522 = ~n1119 | n1513;
  assign n523 = n652 & n1230;
  assign n524 = n1045 & n990;
  assign n525 = n1089 | n1107;
  assign n526 = n370 & (~n110 | n525);
  assign n527 = ~n110 | n1215;
  assign n528 = ~n382 & n1392;
  assign n529 = n526 & n527 & (~n212 | n528);
  assign n530 = n1104 | n1108;
  assign n531 = ~n117 & (~n110 | (~n382 & n530));
  assign n532 = n1088 | n1107;
  assign n533 = ~n213 & n531 & (~n212 | n532);
  assign n534 = n1448 & n1447 & n1446 & n1445 & n1443 & n1444 & n1449 & n1450;
  assign n535 = n1103 | n1206;
  assign n536 = n534 & (~n368 | n535);
  assign n537 = ~n1202 & (~n225 | n430);
  assign n538 = ~n532 & (n110 | ~n1517);
  assign n539 = ~n984 & n1093;
  assign n540 = ~n1110 & (n421 | n539);
  assign n541 = ~n1354 & (~n225 | ~n1161);
  assign n542 = n1455 & n1454 & n800 & n1453 & n1451 & n1452 & n1456 & n1457;
  assign n543 = n1089 | n1122;
  assign n544 = n542 & (~n368 | n543);
  assign n545 = ~n220 & n302;
  assign n546 = ~n225 | n273;
  assign n547 = ~n543 & (n546 | ~n1161);
  assign n548 = (~n430 | n1129) & (n349 | n780);
  assign n549 = (n405 | n990) & (~n220 | n1121);
  assign n550 = (n304 | ~n815) & (~n421 | n1111);
  assign n551 = (n545 | n1133) & (n1463 | n1046);
  assign n552 = ~n547 & (n525 | (~n212 & n1517));
  assign n553 = n2115 & n1388 & n223;
  assign n554 = n551 & n550 & n549 & n548 & n544 & n315 & n552 & n553;
  assign n555 = i_8_ & ~n1083;
  assign n556 = n1092 & ~n1512;
  assign n557 = ~n776 & n555 & n556;
  assign n558 = n1099 & n556;
  assign n559 = n558 & ~n667;
  assign n560 = n260 & n429 & (n796 | n235);
  assign n561 = n554 & n1528 & n529 & n533;
  assign n562 = (~n430 | n530) & (~n539 | n1111);
  assign n563 = (~n110 | n781) & (n1225 | n2107);
  assign n564 = n2133 & n2134 & (n2010 | n1121);
  assign n565 = n2130 & n2120 & n2121 & n2124 & n2123 & n2131 & n2129 & n2128;
  assign n566 = ~n1525 & n565 & n564 & n563 & n562 & n560 & n561 & ~n1520;
  assign n567 = ~n1117 & n556 & ~n776;
  assign n568 = n1074 | ~n1602;
  assign n569 = n568 & (~n1099 | ~n1602);
  assign n570 = n1109 | n1128;
  assign n571 = n495 & n570;
  assign n572 = n1087 | n1201;
  assign n573 = (n469 | n572) & (~n368 | n571);
  assign n574 = ~n368 | n1153;
  assign n575 = n1578 & n1577 & n444 & n1575 & n1576;
  assign n576 = n574 & n575 & (~n368 | ~n465);
  assign n577 = n469 | n1153;
  assign n578 = n469 | n824;
  assign n579 = n469 | n1134;
  assign n580 = n469 | n316;
  assign n581 = n469 | n1133;
  assign n582 = n469 | n726;
  assign n583 = n469 | n727;
  assign n584 = n443 & (n469 | n482);
  assign n585 = n582 & n581 & n580 & n579 & n577 & n578 & n583 & n584;
  assign n586 = ~n368 | n397;
  assign n587 = ~n220 | n1200;
  assign n588 = ~n220 | n1115;
  assign n589 = n1106 | n1108;
  assign n590 = n587 & n588 & (~n220 | n589);
  assign n591 = n469 | n1124;
  assign n592 = n469 | n1204;
  assign n593 = n1110 | n469;
  assign n594 = n226 | n469;
  assign n595 = n1111 | n469;
  assign n596 = n469 | n1338;
  assign n597 = n469 | n1353;
  assign n598 = n442 & (n469 | n401);
  assign n599 = n596 & n595 & n594 & n593 & n591 & n592 & n597 & n598;
  assign n600 = n456 | n245;
  assign n601 = n456 | n613;
  assign n602 = n456 | n1216;
  assign n603 = (~n220 | n1574) & (~n273 | n747);
  assign n604 = ~n220 | n613;
  assign n605 = n1132 | n1201;
  assign n606 = n604 & (n605 | ~n1053);
  assign n607 = n615 & n412 & ~n385 & n401;
  assign n608 = n486 & n1573;
  assign n609 = n608 & n607 & n374;
  assign n610 = n1128 | n1201;
  assign n611 = n269 & n610;
  assign n612 = (n469 | n495) & (~n368 | n611);
  assign n613 = n1107 | n1201;
  assign n614 = n613 | n469;
  assign n615 = n1096 | n1201;
  assign n616 = ~n220 | n615;
  assign n617 = ~n220 | n605;
  assign n618 = n2291 | n456;
  assign n619 = n1932 & n1922 & n1955;
  assign n620 = n756 & n1391;
  assign n621 = n618 & n619 & (~n220 | n620);
  assign n622 = n1209 & n632 & n1130;
  assign n623 = n456 | n622;
  assign n624 = n1466 & n737;
  assign n625 = n456 | n624;
  assign n626 = ~n220 | n1207;
  assign n627 = ~n220 | n1125;
  assign n628 = n1091 | n1096;
  assign n629 = n626 & n627 & (~n220 | n628);
  assign n630 = ~n220 | n1209;
  assign n631 = ~n220 | n1130;
  assign n632 = n1087 | n1091;
  assign n633 = n630 & n631 & (~n220 | n632);
  assign n634 = n456 | n1214;
  assign n635 = n456 | n780;
  assign n636 = n1091 | n1107;
  assign n637 = n634 & n635 & (n456 | n636);
  assign n638 = ~n220 | n1214;
  assign n639 = ~n220 | n780;
  assign n640 = n638 & n639 & (~n220 | n636);
  assign n641 = n456 | n1129;
  assign n642 = n1091 | n1128;
  assign n643 = n1128 | n1196;
  assign n644 = n641 & (n456 | (n642 & n643));
  assign n645 = n1339 & n1465 & n1280;
  assign n646 = n456 | n645;
  assign n647 = n1545 & n1544 & n1543 & n293 & n1542 & n318 & n646;
  assign n648 = n535 & n543 & n1309;
  assign n649 = n647 & (n648 | n456);
  assign n650 = n1005 & n992 & n1006 & n1548 & n792;
  assign n651 = n491 & n1546;
  assign n652 = n1104 | n1196;
  assign n653 = n1133 & n1134;
  assign n654 = n653 & n652 & n651 & n650 & ~n385 & n610;
  assign n655 = n1273 & n1272 & n1271 & n1270 & n1269 & n1268 & ~n221 & n828;
  assign n656 = n1223 & n1241 & n1240 & n1238 & n1239;
  assign n657 = (n456 | n1547) & (~n220 | n654);
  assign n658 = n1148 & n1175 & n827 & n1173 & n1174;
  assign n659 = n2146 & n1764 & n2145 & n1844 & n1405 & n2144;
  assign n660 = n2147 & n621 & n1572 & n1570 & n1563 & n1557;
  assign n661 = n659 & n658 & n657 & n309 & n655 & n656 & n660;
  assign n662 = n993 | n456;
  assign n663 = n662 & (~n220 | n572);
  assign n664 = n1115 & n589;
  assign n665 = n1104 | n1201;
  assign n666 = (n469 | n665) & (~n368 | n664);
  assign n667 = n1214 & n525 & n515;
  assign n668 = ~n558 | n667;
  assign n669 = n1605 & ~n1535 & n668 & n663 & n154 & n661;
  assign n670 = n771 & n1604;
  assign n671 = n405 | n1143;
  assign n672 = n405 | n615;
  assign n673 = n405 | n1217;
  assign n674 = (~n277 | n939) & (n243 | n1573);
  assign n675 = n674 & n673 & n671 & n672;
  assign n676 = ~n405 & (~n645 | ~n1133 | ~n1210);
  assign n677 = ~n243 & (~n233 | ~n1607);
  assign n678 = ~n277 | n482;
  assign n679 = ~n984 & n1086;
  assign n680 = n679 & (~n1228 | ~n1613 | ~n2148);
  assign n681 = n679 & (~n874 | ~n1466);
  assign n682 = ~n1224 | ~n610 | ~n987;
  assign n683 = n679 & (n682 | ~n1537 | ~n1614);
  assign n684 = ~n1086 | n1114;
  assign n685 = n1467 & n944;
  assign n686 = n684 | n685;
  assign n687 = ~n243 & (~n688 | ~n1115);
  assign n688 = n613 & n1200;
  assign n689 = n405 | n688;
  assign n690 = n243 | n1204;
  assign n691 = n237 | n243;
  assign n692 = n243 | n1124;
  assign n693 = n243 | n1338;
  assign n694 = n1110 | n243;
  assign n695 = n243 | n1205;
  assign n696 = n1116 | n243;
  assign n697 = n2154 & (n1111 | n243);
  assign n698 = n695 & n694 & n693 & n692 & n690 & n691 & n696 & n697;
  assign n699 = n1089 | n1102;
  assign n700 = n699 | n405;
  assign n701 = ~n405 & (n278 | ~n1111);
  assign n702 = n231 | ~n430;
  assign n703 = n845 & n397 & n628;
  assign n704 = n702 & (~n430 | n703);
  assign n705 = n349 | n1216;
  assign n706 = n349 | n245;
  assign n707 = (~n430 | n1007) & (~n421 | n747);
  assign n708 = n707 & n705 & n706;
  assign n709 = n143 & n1138;
  assign n710 = n709 & (~n241 | ~n481 | ~n1112);
  assign n711 = n636 & n632;
  assign n712 = ~n421 | n711;
  assign n713 = n349 | n1124;
  assign n714 = n349 | n1204;
  assign n715 = n2290 | n349;
  assign n716 = n349 | n1338;
  assign n717 = n349 | n1353;
  assign n718 = n349 | n237;
  assign n719 = n349 | n1116;
  assign n720 = n2005 & (n349 | (n401 & n491));
  assign n721 = n718 & n717 & n716 & n715 & n713 & n714 & n719 & n720;
  assign n722 = n653 & n316 & n1465;
  assign n723 = n1207 & n1125;
  assign n724 = n482 & n723 & n703 & n722;
  assign n725 = n1095 | n1108;
  assign n726 = n1167 | n1201;
  assign n727 = n1103 | n1167;
  assign n728 = n1153 & n653;
  assign n729 = n728 & n727 & n725 & n645 & n316 & ~n465 & n726;
  assign n730 = n349 | n1280;
  assign n731 = n232 | ~n430;
  assign n732 = (~n430 | n729) & (n349 | n724);
  assign n733 = ~n421 | n809;
  assign n734 = n1316 & n1948 & n1849 & n360 & n1357 & n1850;
  assign n735 = n734 & n733 & n732 & n731 & n359 & n730;
  assign n736 = n572 & n491;
  assign n737 = n652 & n1281;
  assign n738 = n530 & n1105;
  assign n739 = n738 & n737 & n736 & n613 & n610 & n401 & ~n114 & ~n385;
  assign n740 = n1199 & n994;
  assign n741 = ~n918 & n740 & n650 & ~n275 & n412;
  assign n742 = n1637 & n1636 & ~n710 & n712;
  assign n743 = n1337 & n1279 & n308 & n1416 & n1035 & n1368;
  assign n744 = n2152 & n2153 & (n349 | n610);
  assign n745 = n2151 & n2150 & n2149 & n2037 & ~n214 & n2004;
  assign n746 = n1574 & n990 & n1203;
  assign n747 = n665 & n497;
  assign n748 = n610 & n589 & n746 & n747;
  assign n749 = n397 | n243;
  assign n750 = ~n650 | ~n353 | ~n374;
  assign n751 = ~n1458 | ~n1045 | ~n1231;
  assign n752 = ~n243 & (n750 | n751 | ~n986);
  assign n753 = n755 | n970;
  assign n754 = n755 | n1121;
  assign n755 = ~n1086 | n1120;
  assign n756 = n1091 | n1113;
  assign n757 = n753 & n754 & (n755 | n756);
  assign n758 = n1468 & n1227;
  assign n759 = n755 | n758;
  assign n760 = n216 & (~n756 | ~n1231 | ~n1685);
  assign n761 = n496 & n740;
  assign n762 = n755 | n761;
  assign n763 = n216 | ~n755;
  assign n764 = ~n945 | ~n1467;
  assign n765 = n763 & (n764 | ~n1308);
  assign n766 = ~n238 | ~n1232;
  assign n767 = n216 & (n766 | ~n944);
  assign n768 = n985 | n775;
  assign n769 = n770 & n1701;
  assign n770 = n970 & n667;
  assign n771 = n1074 | n1513;
  assign n772 = ~n173 | n1513;
  assign n773 = n304 & n523;
  assign n774 = n772 & (n771 | (n773 & n524));
  assign n775 = n1117 | n1513;
  assign n776 = n1113 | n1201;
  assign n777 = n775 | n776;
  assign n778 = n1215 & n1224;
  assign n779 = n463 & n352;
  assign n780 = n1103 | n1107;
  assign n781 = n1108 | n1128;
  assign n782 = n525 & n780 & n491 & n245 & n778 & n779 & n781 & n632;
  assign n783 = n1708 & n1707 & n445 & n1705 & n1706;
  assign n784 = n1172 & n1267 & (~n110 | n532);
  assign n785 = ~n212 | n1204;
  assign n786 = ~n110 | n1208;
  assign n787 = n493 & n2161 & (~n212 | n782);
  assign n788 = n787 & n786 & n785 & n784 & n783 & n533 & ~n112 & n529;
  assign n789 = n268 | n419;
  assign n790 = ~n218 | n419;
  assign n791 = n789 & n790 & (n779 | n419);
  assign n792 = n642 & n463;
  assign n793 = n225 | n792;
  assign n794 = n645 | n796;
  assign n795 = n1133 & n1606;
  assign n796 = ~n1093 | n1114;
  assign n797 = n794 & (n795 | n796);
  assign n798 = n605 | n469;
  assign n799 = n469 | n643;
  assign n800 = n469 | n1129;
  assign n801 = ~n215 & (~n110 | n1614);
  assign n802 = n2183 & (n456 | n495);
  assign n803 = n2184 & n1485 & n644 & n791 & n1714 & n909;
  assign n804 = n2182 & n2158 & n2000 & n1875 & n1471 & n1325 & ~n115 & n1292;
  assign n805 = n877 & n2021 & n2074 & n2025 & n1792 & n1247 & n1249 & n2181;
  assign n806 = n1963 & n1943 & n2136 & n1942 & n1366 & n1980 & n1367 & n2180;
  assign n807 = n804 & n803 & n802 & n801 & n799 & n800 & n805 & n806;
  assign n808 = n539 & (n465 | ~n1607);
  assign n809 = n605 & n608;
  assign n810 = (n615 | n796) & (~n271 | n809);
  assign n811 = n225 | n1207;
  assign n812 = n225 | n1125;
  assign n813 = n628 & n1213;
  assign n814 = n811 & n812 & (n813 | n225);
  assign n815 = ~n225 | n818;
  assign n816 = n815 & (~n482 | ~n486);
  assign n817 = ~n225 & (~n1401 | ~n1465);
  assign n818 = n1093 & n1099;
  assign n819 = ~n645 | ~n1573;
  assign n820 = n818 & (~n605 | ~n728 | n819);
  assign n821 = ~n850 & (n465 | ~n645);
  assign n822 = ~n419 & (n465 | ~n615);
  assign n823 = ~n501 | n809;
  assign n824 = n1088 | n1167;
  assign n825 = n482 & n235 & n824 & n653 & n486 & n316;
  assign n826 = ~n605 & (~n225 | n368);
  assign n827 = ~n220 | n1143;
  assign n828 = ~n220 | n1123;
  assign n829 = n1634 | n469;
  assign n830 = n456 | ~n465;
  assign n831 = ~n826 & (n1217 | (~n368 & n469));
  assign n832 = n1240 & (~n1053 | (n486 & n1143));
  assign n833 = n1147 & n1764 & n1975 & n1872 & n2142 & n1347 & n1146 & n1145;
  assign n834 = n1736 & n810 & n1677 & n675 & n1000 & n1723 & n1738 & n2179;
  assign n835 = n832 & n831 & n830 & n829 & n827 & n828 & n833 & n834;
  assign n836 = n1395 | n419;
  assign n837 = n1396 | n419;
  assign n838 = n836 & n837 & (n622 | n419);
  assign n839 = ~n1338 | ~n1353;
  assign n840 = ~n225 & (~n632 | ~n651 | n839);
  assign n841 = ~n539 | n622;
  assign n842 = n1395 & n1396;
  assign n843 = n841 & (~n539 | n842);
  assign n844 = ~n539 | n849;
  assign n845 = n1635 & n1123 & n1213;
  assign n846 = n844 & (~n539 | n845);
  assign n847 = n2295 | n850;
  assign n848 = n2294 | n850;
  assign n849 = n231 & n452;
  assign n850 = n1074 | ~n1093;
  assign n851 = n847 & n848 & (n849 | n850);
  assign n852 = n629 & n2167 & (n243 | n1197);
  assign n853 = n1881 & n1803 & n2165 & n1835 & n1900 & n2081 & n1802 & n2164;
  assign n854 = n1795 & n2163 & n1284 & n1344 & n1834 & n1891 & n1010 & n1793;
  assign n855 = n2034 & n2007 & n1961 & n1409 & n1636 & n2151 & n2162 & n1873;
  assign n856 = n853 & n852 & n704 & n130 & n846 & n851 & n854 & n855;
  assign n857 = (n736 | n1398) & (n243 | ~n278);
  assign n858 = (n2171 | n401) & (n2172 | n481);
  assign n859 = (~n539 | n1025) & (n1168 | n1546);
  assign n860 = n2080 & (n632 | (~n212 & n1152));
  assign n861 = n2173 & n494 & n633 & n843 & n856 & n698;
  assign n862 = n1860 & n1446 & n1508 & n1820 & n1452 & n1445 & n1837 & n2170;
  assign n863 = n1906 & n1839 & n1289 & n1323 & n1351 & n1435 & n1493 & n2169;
  assign n864 = n2004 & n1474 & n1411 & n1301 & n2037 & n1853 & n1266 & n2168;
  assign n865 = n862 & n861 & n860 & n859 & n857 & n858 & n863 & n864;
  assign n866 = ~n1154 & (~n268 | ~n987);
  assign n867 = n212 & (n111 | ~n779 | ~n1614);
  assign n868 = n2191 & (~n368 | n463);
  assign n869 = n865 & n1621 & n1662 & n807 & n835 & n1746;
  assign n870 = n2188 & n2190 & (n1769 | n938);
  assign n871 = n2001 & n1911 & n1897 & n1858 & ~n221 & ~n866;
  assign n872 = n1310 & n1791 & n1863 & n1346 & n1282 & n1430 & n2185 & n2187;
  assign n873 = n870 & n869 & n868 & n573 & n612 & n354 & n871 & n872;
  assign n874 = n1574 & n747;
  assign n875 = (n225 | n613) & (~n815 | n874);
  assign n876 = ~n539 | n2297;
  assign n877 = n2166 | n796;
  assign n878 = n876 & n877 & (~n275 | ~n539);
  assign n879 = ~n525 | ~n532;
  assign n880 = n818 & (n275 | ~n636 | n879);
  assign n881 = (~n212 | n780) & (~n368 | n636);
  assign n882 = (n589 | ~n1051) & (~n430 | n2211);
  assign n883 = (n2171 | n412) & (n2172 | n241);
  assign n884 = n1674 & n398 & n640 & n878 & n1001 & n199;
  assign n885 = n1799 & n1188 & n2210 & n1078 & n1869 & n1314 & n1257 & n2208;
  assign n886 = n1181 & n1183 & n1171 & n1862 & n1498 & n1712 & n1426 & n2207;
  assign n887 = n1941 & n1960 & n1825 & n1899 & n1274 & n1833 & n1854 & n2205;
  assign n888 = n885 & n884 & n883 & n882 & n881 & n460 & n886 & n887;
  assign n889 = n419 | ~n892;
  assign n890 = n738 | n419;
  assign n891 = n889 & n890 & (n624 | n419);
  assign n892 = ~n1045 | ~n1203;
  assign n893 = ~n225 & (n892 | ~n1548);
  assign n894 = n1114 | ~n1138;
  assign n895 = n261 & n894;
  assign n896 = n2296 | n796;
  assign n897 = ~n275 & n355;
  assign n898 = n896 & (n897 | n796);
  assign n899 = n2297 | n419;
  assign n900 = ~n275 | n419;
  assign n901 = n419 | n613;
  assign n902 = n2196 & n1011 & (n993 | n225);
  assign n903 = n1263 & n1907 & n1841 & n2031 & n1489 & n1264;
  assign n904 = n898 & n1386 & n2197 & n473 & n457 & n373 & n1669 & n2198;
  assign n905 = n662 & n1882 & n1926 & n2083 & n1840 & n1444 & n2195 & n2194;
  assign n906 = n904 & n903 & n902 & n901 & n899 & n900 & n905;
  assign n907 = ~n243 & (~n530 | ~n1045);
  assign n908 = n1626 & n1625 & n1624 & n1623 & ~n681 & n1622;
  assign n909 = n1709 & n264 & n798 & n797;
  assign n910 = n246 & n350 & n198 & n666;
  assign n911 = n906 & n856 & n835 & n875 & n888 & n1761;
  assign n912 = n2222 & n2217 & n2218 & n2219 & n2220 & n2221 & n2216 & n2215;
  assign n913 = n1326 & n1912 & n1191 & n1254 & n1293 & n1876 & n1379 & n2214;
  assign n914 = n1429 & n1311 & n1496 & n2022 & n2213 & n1250 & n267 & n2212;
  assign n915 = n1231 | n850;
  assign n916 = n2291 | n419;
  assign n917 = n915 & n916 & (n620 | n850);
  assign n918 = ~n756 | ~n1468;
  assign n919 = ~n225 & (n918 | ~n1151);
  assign n920 = n1231 | n419;
  assign n921 = n1151 | n419;
  assign n922 = n920 & n921 & (~n118 | n419);
  assign n923 = ~n225 & (~n776 | ~n994);
  assign n924 = ~n349 & (~n2223 | ~n2224);
  assign n925 = n1093 & n143;
  assign n926 = n925 & (~n1231 | ~n1468 | ~n1613);
  assign n927 = n236 & n756 & n589 & n725;
  assign n928 = ~n496 & (n368 | ~n1769);
  assign n929 = (n1156 | n1612) & (n1152 | n1468);
  assign n930 = n1231 | n243;
  assign n931 = (~n118 | n1460) & (~n368 | n664);
  assign n932 = (~n280 | n1638) & (~n430 | n927);
  assign n933 = n2079 & n1910 & n1378 & n1241 & n1233 & ~n928 & n1189;
  assign n934 = n1022 & n1779 & n1692 & n1719 & n888 & n865 & n917 & n2234;
  assign n935 = n1877 & n1291 & n1870 & n1312 & n1271 & n1507 & n1175 & n2232;
  assign n936 = n1335 & n1361 & n1334 & n1276 & n1299 & n1360 & n1851 & n2230;
  assign n937 = n934 & n933 & n932 & n931 & n929 & n930 & n935 & n936;
  assign n938 = n610 & n495;
  assign n939 = n605 & n486;
  assign n940 = n496 & n944;
  assign n941 = n940 & n939 & n938 & ~n764 & n482 & n747;
  assign n942 = n985 & n1479;
  assign n943 = n942 & ~n764 & ~n385 & n761;
  assign n944 = n942 & n1144 & n1218;
  assign n945 = n1089 | n1206;
  assign n946 = n945 & n495 & n944 & n665;
  assign n947 = n250 & (~n809 | ~n1780);
  assign n948 = ~n419 & (~n824 | ~n1573);
  assign n949 = ~n349 & (~n650 | ~n722 | ~n1127);
  assign n950 = ~n225 & (~n1210 | ~n1465 | ~n1574);
  assign n951 = n518 & (n769 | n1603);
  assign n952 = n951 & n208 & n207 & n175 & ~n183 & n517;
  assign n953 = ~n958 & n2243 & (n569 | n769);
  assign n954 = n953 & n669 & n177;
  assign n955 = n1119 & n556;
  assign n956 = n173 & n556;
  assign n957 = n1119 & n1530;
  assign n958 = n1119 & n1518;
  assign n959 = ~n304 & n1782;
  assign n960 = n1119 & n1702;
  assign n961 = ~n304 & n558;
  assign n962 = ~n304 & n1529;
  assign n963 = ~n990 & n1529;
  assign n964 = ~n1083 & n1530;
  assign n965 = ~n1083 & n1518;
  assign n966 = ~n990 & n1782;
  assign n967 = n558 & ~n990;
  assign n968 = ~n1083 & n1702;
  assign n969 = n670 & ~n979;
  assign n970 = n1113 | n1196;
  assign n971 = ~n652 & ~n2245;
  assign n972 = n173 & n1530;
  assign n973 = n173 & n1518;
  assign n974 = ~n1230 & n1782;
  assign n975 = n173 & n1702;
  assign n976 = n558 & ~n1230;
  assign n977 = ~n1230 & n1529;
  assign n978 = ~n1045 & ~n2245;
  assign n979 = n143 & n1602;
  assign n980 = ~n1701 & (n979 | ~n1604);
  assign n981 = n665 | n775;
  assign n982 = n970 & n1701;
  assign n983 = n2288 & (i_0_ | ~i_2_);
  assign n984 = i_8_ | ~n173;
  assign n985 = n1122 | n1201;
  assign n986 = n1639 & n1638 & n736 & n607 & n740 & n737;
  assign n987 = n305 & n1135;
  assign n988 = n1096 | n1109;
  assign n989 = n632 & n1338;
  assign n990 = n1089 | n1104;
  assign n991 = n988 & n613 & n987 & n268 & n986 & n650 & n989 & n990;
  assign n992 = n776 & n1547;
  assign n993 = n1200 & n664;
  assign n994 = n1109 | n1113;
  assign n995 = n648 & n1354 & n1340;
  assign n996 = n995 & n993 & n992 & n605 & ~n764 & n994;
  assign n997 = n1754 & n1753 & n1752 & n1751 & ~n893 & n1750;
  assign n998 = n1768 & ~n919 & n1767;
  assign n999 = n1739 & ~n840 & n227 & n402;
  assign n1000 = n1727 & n1356 & n1726 & n1725 & n319 & n1724 & n1728 & n1729;
  assign n1001 = n1749 & n1748 & ~n880 & n1484;
  assign n1002 = n328 & n310 & n1315 & n1714 & n413 & n423;
  assign n1003 = n2253 & n2252 & n2251 & n2163 & n2039 & n1237 & ~n116 & n371;
  assign n1004 = ~n539 | n572;
  assign n1005 = n1262 & n995;
  assign n1006 = n1537 & n945 & ~n1027;
  assign n1007 = n589 & n1574;
  assign n1008 = n1007 & n1006 & n1005 & n688 & n651 & ~n114 & ~n385;
  assign n1009 = n620 | n796;
  assign n1010 = ~n539 | n2166;
  assign n1011 = n993 | n796;
  assign n1012 = ~n121 & (~n271 | (n992 & n1780));
  assign n1013 = n1501 & n1500 & n1499 & n1498 & n1496 & n1497 & n1502 & n1503;
  assign n1014 = n1251 & n1250 & n1249 & n1248 & n1246 & n1247 & n1252 & n1253;
  assign n1015 = n1187 & (~n539 | n1008);
  assign n1016 = n1738 & n846 & n843 & n878 & n1798 & n898 & n810 & n797;
  assign n1017 = n1014 & n1013 & n1012 & n1011 & n1009 & n1010 & n1015 & n1016;
  assign n1018 = n1161 | n1308;
  assign n1019 = n1261 | n1161;
  assign n1020 = n1161 | n1309;
  assign n1021 = n1161 | n535;
  assign n1022 = n1772 & n1771 & n1770 & ~n926 & n297 & n322;
  assign n1023 = n1845 & n1303 & (n2240 | n1161);
  assign n1024 = n1022 & n1021 & n363 & n1020 & n1018 & n1019 & n135 & n1023;
  assign n1025 = n572 & n651;
  assign n1026 = n1025 & n1007 & ~n750 & n737 & n613 & ~n118 & n352;
  assign n1027 = n766 | ~n1467;
  assign n1028 = ~n419 & (~n945 | ~n992 | n1027);
  assign n1029 = n1802 & n1801 & n899 & n1800 & n1799 & n901 & n1803 & n1804;
  assign n1030 = n1723 & n791 & n1495;
  assign n1031 = n1260 & n2226 & n2196 & n1709 & n2165 & n1731 & n1195 & n2255;
  assign n1032 = n838 & n851 & n891 & n922 & n1029 & n917 & n1030 & n1031;
  assign n1033 = n796 & n243;
  assign n1034 = ~n456 & (~n1209 | ~n1339);
  assign n1035 = n1412 & n1411 & n1410 & n1409 & n1407 & n1408 & n1413 & n1414;
  assign n1036 = n1383 & n1382 & n1381 & n1380 & n1379 & n1378 & ~n369 & n799;
  assign n1037 = n365 & (~n539 | n1338);
  assign n1038 = (~n430 | n643) & (n349 | n1214);
  assign n1039 = (n1033 | n726) & (n1463 | n1044);
  assign n1040 = ~n1034 & (n225 | (n1045 & n1340));
  assign n1041 = n2256 & (~n220 | n970);
  assign n1042 = n1039 & n1038 & n1037 & n335 & n1035 & n1036 & n1040 & n1041;
  assign n1043 = ~n1053 & ~n815 & ~n421 & ~n220 & n243;
  assign n1044 = n515 & n1211;
  assign n1045 = n1102 | n1201;
  assign n1046 = n1089 | n1096;
  assign n1047 = n1046 & n525 & n1044 & n1045;
  assign n1048 = n699 & n1468 & n463;
  assign n1049 = n776 & n610 & n1048 & n665;
  assign n1050 = ~n2107 & (~n305 | ~n1226);
  assign n1051 = ~n243 | ~n850;
  assign n1052 = n1051 & (~n353 | ~n1391);
  assign n1053 = n368 | ~n469;
  assign n1054 = ~n572 & (n1053 | ~n1398);
  assign n1055 = ~n1281 & (~n243 | n381 | n501);
  assign n1056 = ~n1054 & (n613 | (~n277 & n1166));
  assign n1057 = ~n1052 & (n1159 | (n482 & n1805));
  assign n1058 = n1670 & n2257 & (n2096 | n1049);
  assign n1059 = n2258 & n2259 & n2261 & n2260;
  assign n1060 = n2154 & n876 & n1571 & n1079 & n1655 & n1665 & n2158 & n1646;
  assign n1061 = n1645 & n2150 & n794 & n841 & n1642 & n1739 & n1222 & n1147;
  assign n1062 = n1798 & n1029 & n1552 & n606 & n1766 & n742 & n1042 & n2273;
  assign n1063 = n2264 & n2265 & n2266 & n2267 & n2269 & n2268 & n2263 & n2262;
  assign n1064 = n1061 & n1060 & n1059 & n1058 & n1056 & n1057 & n1062 & n1063;
  assign n1065 = ~n532 & (n212 | n503);
  assign n1066 = ~n226 & (~n225 | ~n349 | ~n1154);
  assign n1067 = n539 & (~n231 | ~n726 | ~n1353);
  assign n1068 = n2287 & (n796 | n824);
  assign n1069 = ~n1536 & ~n1534 & n1042 & n1528;
  assign n1070 = (n1154 | n1219) & (n1164 | n1209);
  assign n1071 = n2286 & (~n273 | n1227);
  assign n1072 = n2284 & n2285 & (n2010 | n970);
  assign n1073 = n2278 & n2279 & n2280 & n2281 & n2283 & n2282 & n2276 & n2275;
  assign n1074 = i_8_ | n123;
  assign n1075 = n1425 & n1464;
  assign n1076 = n1389 & n1386 & n1036 & n1402 & n1377;
  assign n1077 = n2140 & (~n368 | (n572 & n874));
  assign n1078 = ~n368 | n1200;
  assign n1079 = ~n368 | n613;
  assign n1080 = (~n368 | n609) & (n940 | ~n1053);
  assign n1081 = n2139 & n2138 & n2137 & n2136 & n2135 & n2034 & ~n108 & n2007;
  assign n1082 = n1601 & n576 & n1592 & n198 & n590 & n599 & n573 & n2141;
  assign n1083 = ~i_6_ | i_7_;
  assign n1084 = ~i_5_ | i_3_ | i_4_;
  assign n1085 = ~i_2_ & ~i_0_ & ~i_1_;
  assign n1086 = ~n1084 & n1085;
  assign n1087 = i_15_ | n481;
  assign n1088 = ~i_14_ | i_12_ | ~i_13_;
  assign n1089 = ~i_14_ | i_12_ | i_13_;
  assign n1090 = ~i_15_ | n481;
  assign n1091 = i_14_ | ~i_12_ | ~i_13_;
  assign n1092 = ~i_5_ & ~i_3_ & i_4_;
  assign n1093 = n1085 & n1092;
  assign n1094 = ~i_11_ | ~i_9_ | ~i_10_;
  assign n1095 = ~i_15_ | n1094;
  assign n1096 = i_15_ | n1094;
  assign n1097 = n1088 | n1096;
  assign n1098 = n1046 & n1097;
  assign n1099 = ~i_8_ & ~n1083;
  assign n1100 = i_5_ & ~i_3_ & i_4_;
  assign n1101 = n1085 & n1100;
  assign n1102 = ~i_15_ | n265;
  assign n1103 = i_14_ | ~i_12_ | i_13_;
  assign n1104 = i_15_ | n265;
  assign n1105 = n990 & n244;
  assign n1106 = ~i_15_ | n241;
  assign n1107 = i_15_ | n241;
  assign n1108 = ~i_14_ | ~i_12_ | ~i_13_;
  assign n1109 = ~i_14_ | ~i_12_ | i_13_;
  assign n1110 = n1087 | n1088;
  assign n1111 = n1087 | n1089;
  assign n1112 = i_11_ | ~i_9_ | i_10_;
  assign n1113 = i_15_ | n1112;
  assign n1114 = ~i_8_ | ~n173;
  assign n1115 = n1107 | n1109;
  assign n1116 = n1087 | n1109;
  assign n1117 = ~i_8_ | n123;
  assign n1118 = n1106 | n1109;
  assign n1119 = i_6_ & i_7_;
  assign n1120 = ~i_8_ | ~n1119;
  assign n1121 = n1103 | n1113;
  assign n1122 = i_15_ | ~n142;
  assign n1123 = n1096 | n1108;
  assign n1124 = n1087 | n1108;
  assign n1125 = n1096 | n1103;
  assign n1126 = ~i_15_ | n478;
  assign n1127 = n1109 | n1126;
  assign n1128 = i_15_ | n478;
  assign n1129 = n1103 | n1128;
  assign n1130 = n1087 | n1103;
  assign n1131 = ~i_11_ | i_9_ | ~i_10_;
  assign n1132 = i_15_ | n1131;
  assign n1133 = n1089 | n1132;
  assign n1134 = n1088 | n1132;
  assign n1135 = n1088 | n1128;
  assign n1136 = n1107 | n1108;
  assign n1137 = ~i_5_ & ~i_3_ & ~i_4_;
  assign n1138 = n1085 & n1137;
  assign n1139 = ~n555 | ~n1138;
  assign n1140 = n241 | n1139;
  assign n1141 = n265 | n477;
  assign n1142 = n265 | n1139;
  assign n1143 = n1109 | n1132;
  assign n1144 = n1109 | n1122;
  assign n1145 = n1123 | n456;
  assign n1146 = n456 | n1097;
  assign n1147 = n456 | n1046;
  assign n1148 = n1147 & n1145 & n1146;
  assign n1149 = n1108 | n1113;
  assign n1150 = n1088 | n1113;
  assign n1151 = n304 & n1149 & n1150;
  assign n1152 = ~n430 & ~n818;
  assign n1153 = n1108 | n1132;
  assign n1154 = ~n539 & n1152;
  assign n1155 = ~n1051 & n1154;
  assign n1156 = ~n250 & n1155;
  assign n1157 = n488 & n1156;
  assign n1158 = ~n273 & ~n1053;
  assign n1159 = n1157 & n1158;
  assign n1160 = n684 & n1159;
  assign n1161 = ~n1093 | n1120;
  assign n1162 = n1161 & n1160;
  assign n1163 = ~i_15_ | n1112;
  assign n1164 = ~n1051 & ~n271 & n302;
  assign n1165 = n850 & n1154;
  assign n1166 = n469 & n1165;
  assign n1167 = ~i_15_ | n1131;
  assign n1168 = ~n220 & n850;
  assign n1169 = ~n110 | n1115;
  assign n1170 = ~n110 | n245;
  assign n1171 = ~n212 | n1115;
  assign n1172 = n1171 & n1169 & n1170;
  assign n1173 = n1116 | n456;
  assign n1174 = n988 | n456;
  assign n1175 = ~n220 | n994;
  assign n1176 = n1781 | n755;
  assign n1177 = n755 | n1144;
  assign n1178 = n225 | n1143;
  assign n1179 = n456 | n1143;
  assign n1180 = n1179 & n1178 & n706 & n671 & n1176 & n1177 & n600;
  assign n1181 = n355 | ~n539;
  assign n1182 = n245 | n796;
  assign n1183 = ~n539 | n1115;
  assign n1184 = n1151 | n796;
  assign n1185 = ~n539 | n1151;
  assign n1186 = n2026 & n2025 & n2024 & n2023 & n2021 & n2022;
  assign n1187 = n1186 & n1185 & n1184 & n1183 & n1181 & n1182;
  assign n1188 = n1115 | n850;
  assign n1189 = n1151 | n850;
  assign n1190 = n1781 | n419;
  assign n1191 = n738 | n850;
  assign n1192 = n355 | n850;
  assign n1193 = n419 | n245;
  assign n1194 = n2033 & n2032 & n1732 & n2031 & n2029 & n2030;
  assign n1195 = n1193 & n1192 & n1191 & n1190 & n1188 & n1189 & n1194;
  assign n1196 = i_14_ | i_12_ | ~i_13_;
  assign n1197 = n1095 | n1196;
  assign n1198 = n1088 | n1106;
  assign n1199 = n1163 | n1196;
  assign n1200 = n1106 | n1196;
  assign n1201 = i_13_ | i_12_ | i_14_;
  assign n1202 = n1102 | n1103;
  assign n1203 = n1202 & n484;
  assign n1204 = n1088 | n1090;
  assign n1205 = n1090 | n1196;
  assign n1206 = ~i_15_ | ~n142;
  assign n1207 = n1096 | n1196;
  assign n1208 = n1088 | n1126;
  assign n1209 = n1087 | n1196;
  assign n1210 = n727 & n316;
  assign n1211 = n1095 | n1201;
  assign n1212 = n1095 | n1103;
  assign n1213 = n1211 & n1212;
  assign n1214 = n1107 | n1196;
  assign n1215 = n1103 | n1106;
  assign n1216 = n1102 | n1196;
  assign n1217 = n1167 | n1196;
  assign n1218 = n1196 | n1206;
  assign n1219 = n1091 | n1095;
  assign n1220 = n456 | n1219;
  assign n1221 = n456 | n1212;
  assign n1222 = n456 | n1211;
  assign n1223 = n1222 & n1220 & n1221;
  assign n1224 = n1091 | n1126;
  assign n1225 = n1103 | n1126;
  assign n1226 = n1126 | n1201;
  assign n1227 = n1088 | n1163;
  assign n1228 = n1091 | n1163;
  assign n1229 = n1103 | n1163;
  assign n1230 = n1163 | n1201;
  assign n1231 = n1230 & n1228 & n1229;
  assign n1232 = n1122 | n1196;
  assign n1233 = ~n818 | n1231;
  assign n1234 = ~n818 | ~n892;
  assign n1235 = ~n818 | n1205;
  assign n1236 = n225 | n1199;
  assign n1237 = n1236 & n1235 & n1233 & n1234;
  assign n1238 = n456 | n1205;
  assign n1239 = n456 | n1197;
  assign n1240 = ~n220 | n1217;
  assign n1241 = ~n220 | n1199;
  assign n1242 = n1806 | n755;
  assign n1243 = n755 | n1218;
  assign n1244 = n456 | n1217;
  assign n1245 = n602 & n1244 & n705 & n673 & n1242 & n1243 & n262;
  assign n1246 = n1395 | n796;
  assign n1247 = n268 | n796;
  assign n1248 = n796 | n1205;
  assign n1249 = n796 | n269;
  assign n1250 = ~n539 | ~n892;
  assign n1251 = n796 | ~n892;
  assign n1252 = n796 | n1216;
  assign n1253 = n1997 & n1998;
  assign n1254 = n850 | ~n892;
  assign n1255 = ~n275 | n850;
  assign n1256 = n419 | n1216;
  assign n1257 = n850 | n1200;
  assign n1258 = n1806 | n419;
  assign n1259 = n2002 & n2001 & n1730 & n900 & n1999 & n2000;
  assign n1260 = n1259 & n1258 & n1257 & n1256 & n1254 & n1255;
  assign n1261 = n1109 | n1206;
  assign n1262 = n1108 | n1122;
  assign n1263 = ~n110 | n1118;
  assign n1264 = ~n110 | n1136;
  assign n1265 = ~n110 | n1127;
  assign n1266 = ~n212 | n237;
  assign n1267 = n1266 & n1265 & n1263 & n1264;
  assign n1268 = ~n220 | n346;
  assign n1269 = ~n220 | n530;
  assign n1270 = ~n220 | n1136;
  assign n1271 = ~n220 | n1149;
  assign n1272 = n456 | n1136;
  assign n1273 = n1977 & n1975 & n1976;
  assign n1274 = ~n430 | n1118;
  assign n1275 = n349 | n1149;
  assign n1276 = ~n430 | n1149;
  assign n1277 = n349 | n1118;
  assign n1278 = n1981 & n1980 & n1733 & n1756 & n1978 & n1979;
  assign n1279 = n1278 & n292 & n1277 & n1276 & n1274 & n1275;
  assign n1280 = n1103 | n1132;
  assign n1281 = n1103 | n1104;
  assign n1282 = ~n818 | n1129;
  assign n1283 = ~n818 | n1130;
  assign n1284 = ~n818 | n1125;
  assign n1285 = n225 | n1130;
  assign n1286 = n225 | n780;
  assign n1287 = n225 | n1121;
  assign n1288 = ~n818 | n1111;
  assign n1289 = ~n220 | n1111;
  assign n1290 = ~n220 | n1281;
  assign n1291 = ~n220 | n304;
  assign n1292 = n456 | n305;
  assign n1293 = ~n220 | n990;
  assign n1294 = ~n220 | n525;
  assign n1295 = ~n220 | n1129;
  assign n1296 = n1958 & n1956 & n1957;
  assign n1297 = n349 | n304;
  assign n1298 = n349 | n1121;
  assign n1299 = n304 | ~n430;
  assign n1300 = ~n430 | n1121;
  assign n1301 = ~n430 | n1130;
  assign n1302 = n1963 & n1962 & n1961 & n1960 & n1959 & n1757;
  assign n1303 = n238 | n1161;
  assign n1304 = n755 | n238;
  assign n1305 = n238 | n684;
  assign n1306 = n1727 & n1966 & n730 & n1965 & n1724 & n1964;
  assign n1307 = n1091 | n1106;
  assign n1308 = n1088 | n1206;
  assign n1309 = n1091 | n1206;
  assign n1310 = ~n818 | n1208;
  assign n1311 = n345 | ~n818;
  assign n1312 = ~n818 | n1227;
  assign n1313 = ~n818 | n1204;
  assign n1314 = ~n818 | n1198;
  assign n1315 = n1314 & n1313 & n1312 & n1310 & n1311;
  assign n1316 = n349 | n824;
  assign n1317 = n405 | n824;
  assign n1318 = n405 | n1308;
  assign n1319 = n405 | n1309;
  assign n1320 = n225 | n824;
  assign n1321 = n1018 & n1935 & n1020 & n191;
  assign n1322 = n1321 & n1320 & n1319 & n1318 & n1316 & n1317;
  assign n1323 = ~n220 | n226;
  assign n1324 = ~n220 | n345;
  assign n1325 = n456 | n1224;
  assign n1326 = ~n220 | n484;
  assign n1327 = ~n220 | n1307;
  assign n1328 = ~n220 | n1208;
  assign n1329 = n1938 & n1936 & n1937;
  assign n1330 = n1327 & n317 & n1326 & n1325 & n1323 & n1324 & n1328 & n1329;
  assign n1331 = n349 | n1227;
  assign n1332 = n349 | n1228;
  assign n1333 = n349 | n1308;
  assign n1334 = ~n430 | n1227;
  assign n1335 = ~n430 | n1228;
  assign n1336 = n1944 & n1943 & n1942 & n1941 & n1939 & n1940;
  assign n1337 = n1336 & n1335 & n1334 & n1333 & n1331 & n1332;
  assign n1338 = n1090 | n1201;
  assign n1339 = n1132 | n1196;
  assign n1340 = n1201 | n1206;
  assign n1341 = ~n818 | n1209;
  assign n1342 = n225 | n1214;
  assign n1343 = n225 | n970;
  assign n1344 = ~n818 | n1207;
  assign n1345 = n225 | n1209;
  assign n1346 = n643 | ~n818;
  assign n1347 = ~n220 | n726;
  assign n1348 = ~n220 | n1226;
  assign n1349 = ~n220 | n643;
  assign n1350 = n456 | n1226;
  assign n1351 = ~n220 | n1338;
  assign n1352 = n1926 & n1925 & n1923 & n1924;
  assign n1353 = n1090 | n1103;
  assign n1354 = n1088 | n1122;
  assign n1355 = n405 | n535;
  assign n1356 = n225 | n1134;
  assign n1357 = n349 | n727;
  assign n1358 = n405 | n1354;
  assign n1359 = n187 & n1021 & n1358 & n1357 & n1355 & n1356 & n192;
  assign n1360 = ~n430 | n1150;
  assign n1361 = ~n430 | n1229;
  assign n1362 = n349 | n1150;
  assign n1363 = n349 | n1229;
  assign n1364 = ~n430 | n1353;
  assign n1365 = n349 | n1202;
  assign n1366 = n349 | n1135;
  assign n1367 = n349 | n1225;
  assign n1368 = n1365 & n1364 & n1363 & n1362 & n1360 & n1361 & n1366 & n1367;
  assign n1369 = n469 | n1118;
  assign n1370 = ~n368 | n530;
  assign n1371 = n469 | n346;
  assign n1372 = ~n368 | n1118;
  assign n1373 = ~n368 | n1136;
  assign n1374 = n1821 & n1819 & n1820;
  assign n1375 = n1822 & (~n368 | (n236 & n1262));
  assign n1376 = n1817 & n1816 & n1815 & n1814 & n1812 & n1813 & n1818 & n1811;
  assign n1377 = n1374 & n1373 & n1372 & n1371 & n1369 & n1370 & n1375 & n1376;
  assign n1378 = ~n368 | n970;
  assign n1379 = ~n368 | n652;
  assign n1380 = n469 | n1232;
  assign n1381 = n469 | n1045;
  assign n1382 = n1841 & n1840 & n1839 & n1838 & n1836 & n1837;
  assign n1383 = n1835 & n1834 & n1833 & n1832 & n1830 & n1831 & n1829;
  assign n1384 = n469 | n532;
  assign n1385 = n469 | n525;
  assign n1386 = n432 & n1384 & n1385;
  assign n1387 = n469 | n1097;
  assign n1388 = n469 | n1046;
  assign n1389 = n433 & n1387 & n1388;
  assign n1390 = n1281 & n1130;
  assign n1391 = n970 & n1121;
  assign n1392 = n1202 & n738;
  assign n1393 = n419 & n1156;
  assign n1394 = n652 & n1339;
  assign n1395 = ~n278 & n1338;
  assign n1396 = n1111 & n1124 & n1110;
  assign n1397 = ~n1051 & n1152;
  assign n1398 = ~n220 & n1397;
  assign n1399 = ~n1053 & ~n679 & n405 & ~n539;
  assign n1400 = n349 & n1398;
  assign n1401 = n726 & n1210;
  assign n1402 = ~n368 | n2298;
  assign n1403 = n225 | n235;
  assign n1404 = n225 | n1153;
  assign n1405 = n456 | n1262;
  assign n1406 = n1850 & n1849 & n1598 & n1848 & n1675 & n1847;
  assign n1407 = n349 | n1226;
  assign n1408 = n349 | n643;
  assign n1409 = ~n430 | n1207;
  assign n1410 = n349 | n1209;
  assign n1411 = ~n430 | n1338;
  assign n1412 = n349 | n1045;
  assign n1413 = n349 | n652;
  assign n1414 = n1856 & n1855 & n1854 & n1853 & n1851 & n1852;
  assign n1415 = ~n430 | n2290;
  assign n1416 = n1415 & n417 & n356 & n354 & ~n109 & n350;
  assign n1417 = ~n368 | n1228;
  assign n1418 = ~n368 | n1208;
  assign n1419 = n469 | n1228;
  assign n1420 = n469 | n1308;
  assign n1421 = ~n368 | n1204;
  assign n1422 = ~n368 | n484;
  assign n1423 = n469 | n345;
  assign n1424 = n1861 & n1860 & n1859 & n1858 & ~n215 & n1857;
  assign n1425 = n1422 & n1421 & n1420 & n1419 & n1417 & n1418 & n1423 & n1424;
  assign n1426 = ~n818 | n1118;
  assign n1427 = n225 | n236;
  assign n1428 = n225 | n1118;
  assign n1429 = n346 | ~n818;
  assign n1430 = n781 | ~n818;
  assign n1431 = n225 | n1127;
  assign n1432 = n1863 & n1862 & n1741;
  assign n1433 = n1869 & n1868 & n1867 & n1866 & n1864 & n1865 & n1870 & n1871;
  assign n1434 = ~n220 | n1110;
  assign n1435 = ~n220 | n1353;
  assign n1436 = ~n220 | n1135;
  assign n1437 = n456 | n1225;
  assign n1438 = n456 | n1215;
  assign n1439 = ~n220 | n1215;
  assign n1440 = n1874 & n1872 & n1873;
  assign n1441 = n1880 & n1879 & n1878 & n1877 & n1875 & n1876 & n1881 & n1882;
  assign n1442 = n1439 & n1438 & n1437 & n1436 & n1434 & n1435 & n1440 & n1441;
  assign n1443 = ~n368 | n1225;
  assign n1444 = n469 | n1215;
  assign n1445 = ~n368 | n1110;
  assign n1446 = ~n368 | n1353;
  assign n1447 = n469 | n535;
  assign n1448 = n1896 & n1894 & n1895;
  assign n1449 = n1897 & (~n368 | n1354);
  assign n1450 = n1892 & n1891 & n1890 & n1889 & n1887 & n1888 & n1893 & n1886;
  assign n1451 = n469 | n1121;
  assign n1452 = ~n368 | n1111;
  assign n1453 = n469 | n238;
  assign n1454 = n469 | n990;
  assign n1455 = n1911 & n1909 & n1910;
  assign n1456 = n1912 & (n238 | ~n368);
  assign n1457 = n1904 & n1908 & n1907 & n1906 & n1742 & n1905;
  assign n1458 = n1227 & n236;
  assign n1459 = n850 & ~n212 & n302;
  assign n1460 = ~n368 & ~n1051;
  assign n1461 = ~n430 & n1460;
  assign n1462 = n419 & ~n539;
  assign n1463 = n225 & ~n250;
  assign n1464 = (~n368 | n1309) & (~n1053 | n1227);
  assign n1465 = n1091 | n1132;
  assign n1466 = n1091 | n1104;
  assign n1467 = n1091 | n1122;
  assign n1468 = n1089 | n1163;
  assign n1469 = n469 | n756;
  assign n1470 = n469 | n1467;
  assign n1471 = n469 | n642;
  assign n1472 = n469 | n1466;
  assign n1473 = n2083 & n2082 & n2081 & n2080 & n2078 & n2079;
  assign n1474 = n481 | n477;
  assign n1475 = n481 | n1139;
  assign n1476 = n478 | n1139;
  assign n1477 = ~n539 & n1400;
  assign n1478 = n225 & n1400;
  assign n1479 = n1108 | n1206;
  assign n1480 = n628 & n711;
  assign n1481 = n1466 & n756 & n642;
  assign n1482 = ~n815 & n1164;
  assign n1483 = ~n763 & ~n925;
  assign n1484 = n225 | n725;
  assign n1485 = n1484 & n916 & ~n112 & n618;
  assign n1486 = n456 | n486;
  assign n1487 = ~n465 | n796;
  assign n1488 = n1487 & n189 & n1486 & n483;
  assign n1489 = n2296 | n419;
  assign n1490 = n1755 | n419;
  assign n1491 = n2296 | n850;
  assign n1492 = n849 | n419;
  assign n1493 = n2291 | n850;
  assign n1494 = n419 | n491;
  assign n1495 = n1494 & n1493 & n1492 & n1491 & n1489 & n1490;
  assign n1496 = ~n539 | n1755;
  assign n1497 = n1755 | n796;
  assign n1498 = ~n539 | n2296;
  assign n1499 = ~n118 | n796;
  assign n1500 = ~n118 | ~n539;
  assign n1501 = ~n539 | n2291;
  assign n1502 = n796 | n491;
  assign n1503 = n2074 & n2072 & n2073;
  assign n1504 = n456 | n491;
  assign n1505 = n456 | n725;
  assign n1506 = n849 | n456;
  assign n1507 = ~n118 | ~n220;
  assign n1508 = ~n220 | n2291;
  assign n1509 = ~n120 | n456;
  assign n1510 = n2077 & ~n466 & n464 & n460 & n453 & n457;
  assign n1511 = n1508 & n1507 & n830 & n1506 & n1504 & n1505 & n1509 & n1510;
  assign n1512 = i_2_ | i_0_ | ~i_1_;
  assign n1513 = ~n1137 | n1512;
  assign n1514 = ~n555 | n1513;
  assign n1515 = i_0_ & ~i_1_;
  assign n1516 = n1215 & n1212;
  assign n1517 = ~n368 & n1463;
  assign n1518 = n1100 & n1515;
  assign n1519 = ~n271 & ~n679;
  assign n1520 = n557 | n559 | n958 | n181;
  assign n1521 = n558 & ~n970;
  assign n1522 = n558 & ~n652;
  assign n1523 = n558 & ~n1045;
  assign n1524 = n1788 | n973 | n965;
  assign n1525 = n967 | n1521 | n1522 | n976 | n1523 | n955 | n961 | n1524;
  assign n1526 = n1384 & (n1463 | (n1516 & n1097));
  assign n1527 = n2116 & n2117 & n2118 & n1442 & n536 & n344;
  assign n1528 = n1527 & n1526 & n1387 & ~n541 & ~n540 & ~n538 & n224 & ~n537;
  assign n1529 = n556 & ~n1074;
  assign n1530 = n1092 & n1515;
  assign n1531 = ~n652 & n1529;
  assign n1532 = ~n1045 & n1529;
  assign n1533 = n962 | n1789 | n1786 | n964 | n957 | n972;
  assign n1534 = n963 | n977 | n1531 | n1533 | n1532 | n956;
  assign n1535 = n169 | n165 | n161;
  assign n1536 = n1535 | n182 | n567;
  assign n1537 = n269 & n570;
  assign n1538 = ~n220 | n988;
  assign n1539 = ~n220 | n1197;
  assign n1540 = ~n220 | n725;
  assign n1541 = n1540 & n1539 & n1538 & n616;
  assign n1542 = n456 | n1133;
  assign n1543 = n456 | n1134;
  assign n1544 = n456 | n727;
  assign n1545 = n456 | n726;
  assign n1546 = n1205 & n1116;
  assign n1547 = n495 & n940;
  assign n1548 = n1466 & n699;
  assign n1549 = n456 | ~n1027;
  assign n1550 = n456 | n615;
  assign n1551 = n2142 & n2143;
  assign n1552 = n644 & n1549 & n637 & n640 & n633 & n629 & n1550 & n1551;
  assign n1553 = n456 | n990;
  assign n1554 = n456 | n244;
  assign n1555 = n456 | n1202;
  assign n1556 = n456 | n1045;
  assign n1557 = n1556 & n1555 & n1554 & n295 & n1553 & n320 & n625;
  assign n1558 = n456 | n1150;
  assign n1559 = n456 | n304;
  assign n1560 = ~n118 | n456;
  assign n1561 = n456 | n1229;
  assign n1562 = n456 | n1230;
  assign n1563 = n1561 & n321 & n296 & n1560 & n1558 & n1559 & n1562;
  assign n1564 = n1111 | n456;
  assign n1565 = n226 | n456;
  assign n1566 = n1124 | n456;
  assign n1567 = n1110 | n456;
  assign n1568 = n456 | n1353;
  assign n1569 = n456 | n1338;
  assign n1570 = n1569 & n1568 & n1567 & n1566 & n1564 & n1565 & n623;
  assign n1571 = n456 | n605;
  assign n1572 = n1244 & n1179 & n1486 & n1541 & n1571 & n617;
  assign n1573 = n1217 & n1143;
  assign n1574 = n1216 & n245;
  assign n1575 = n469 | n1212;
  assign n1576 = n469 | n1211;
  assign n1577 = n469 | n1125;
  assign n1578 = n469 | n1207;
  assign n1579 = ~n368 | n1123;
  assign n1580 = ~n368 | n1097;
  assign n1581 = n232 | ~n368;
  assign n1582 = n231 | ~n368;
  assign n1583 = ~n368 | n1046;
  assign n1584 = ~n368 | n1219;
  assign n1585 = n1584 & n1583 & n1582 & n1581 & n1579 & n1580 & n586;
  assign n1586 = n469 | n1200;
  assign n1587 = n469 | n589;
  assign n1588 = n469 | n1115;
  assign n1589 = n1588 & n1587 & n1586 & n614;
  assign n1590 = n469 | n994;
  assign n1591 = n469 | n1199;
  assign n1592 = n829 & n1590 & n1591;
  assign n1593 = n316 | ~n368;
  assign n1594 = ~n368 | n727;
  assign n1595 = ~n368 | n1134;
  assign n1596 = ~n368 | n1133;
  assign n1597 = ~n368 | n726;
  assign n1598 = n469 | n235;
  assign n1599 = ~n368 | n1280;
  assign n1600 = n1964 & n2084 & n1929 & n585 & n362 & n1585;
  assign n1601 = n1598 & n1597 & n1596 & n1595 & n1593 & n1594 & n1599 & n1600;
  assign n1602 = n1100 & ~n1512;
  assign n1603 = n1512 | n1084 | ~n1099;
  assign n1604 = n1603 & n569;
  assign n1605 = n1512 | n123 | ~n222;
  assign n1606 = n1401 & n1153 & n1134;
  assign n1607 = n645 & n795;
  assign n1608 = n405 | n726;
  assign n1609 = n405 | n1153;
  assign n1610 = n405 | n1134;
  assign n1611 = n1610 & n1609 & ~n676 & n1608;
  assign n1612 = n776 & n740;
  assign n1613 = n1612 & n756 & n496;
  assign n1614 = n495 & n642;
  assign n1615 = ~n679 | n1225;
  assign n1616 = ~n679 | n1226;
  assign n1617 = ~n679 | n779;
  assign n1618 = ~n679 | n781;
  assign n1619 = ~n679 | n1129;
  assign n1620 = n643 | ~n679;
  assign n1621 = n1620 & n1619 & n1618 & n1617 & n1616 & ~n683 & n1615;
  assign n1622 = ~n679 | n1281;
  assign n1623 = n652 | ~n679;
  assign n1624 = ~n679 | n1755;
  assign n1625 = ~n679 | n738;
  assign n1626 = ~n679 | ~n892;
  assign n1627 = ~n679 | n1229;
  assign n1628 = ~n679 | n1230;
  assign n1629 = ~n118 | ~n679;
  assign n1630 = ~n679 | n1149;
  assign n1631 = ~n679 | n1121;
  assign n1632 = ~n679 | n970;
  assign n1633 = n1632 & n1631 & n1630 & n1629 & n1628 & ~n680 & n1627;
  assign n1634 = n615 & n988 & n1197;
  assign n1635 = n1219 & n1098;
  assign n1636 = ~n709 | n1094;
  assign n1637 = n349 | n572;
  assign n1638 = n1151 & n620;
  assign n1639 = n1468 & n725 & n530 & n244 & ~n278 & n1197;
  assign n1640 = n243 | n1211;
  assign n1641 = n988 | n243;
  assign n1642 = n1762 | n243;
  assign n1643 = n1983 & n1947 & n1984 & n1946 & n337 & n1969;
  assign n1644 = n405 | n1205;
  assign n1645 = n405 | n572;
  assign n1646 = n622 | n405;
  assign n1647 = n405 | n491;
  assign n1648 = n1116 | n405;
  assign n1649 = n1927 & n1985 & n338;
  assign n1650 = n405 | n530;
  assign n1651 = n405 | n244;
  assign n1652 = n405 | n346;
  assign n1653 = n405 | n345;
  assign n1654 = n405 | n1045;
  assign n1655 = n624 | n405;
  assign n1656 = n243 | n1226;
  assign n1657 = n243 | n305;
  assign n1658 = n243 | n1224;
  assign n1659 = n243 | n781;
  assign n1660 = n243 | n1127;
  assign n1661 = n243 | n1208;
  assign n1662 = n340 & n1659 & n1658 & n1657 & n339 & n1656 & n1660 & n1661;
  assign n1663 = n405 | n515;
  assign n1664 = n1115 | n405;
  assign n1665 = n2297 | n405;
  assign n1666 = n405 | n1307;
  assign n1667 = n405 | n1215;
  assign n1668 = n1970 & n1988 & n1913;
  assign n1669 = n1666 & n416 & n689 & n1665 & n1663 & n1664 & n1667 & n1668;
  assign n1670 = n2297 | n243;
  assign n1671 = n243 | n1215;
  assign n1672 = n243 | n515;
  assign n1673 = n1990 & n1952 & n1987 & n1951 & n1915 & n1967;
  assign n1674 = n1673 & n1672 & n1671 & n1670 & ~n687 & n136 & n137;
  assign n1675 = n405 | n235;
  assign n1676 = n1762 | n405;
  assign n1677 = n1676 & n1675 & n1611 & n1317 & ~n677 & n678;
  assign n1678 = n405 | n1046;
  assign n1679 = n405 | n1219;
  assign n1680 = n405 | n1123;
  assign n1681 = n405 | n1097;
  assign n1682 = n405 | n1212;
  assign n1683 = n405 | n1211;
  assign n1684 = n1683 & n1682 & n1681 & n1680 & n1678 & n1679 & n406;
  assign n1685 = n758 & n496 & n776;
  assign n1686 = ~n216 | n1121;
  assign n1687 = ~n216 | n970;
  assign n1688 = ~n216 | n1199;
  assign n1689 = ~n216 | n236;
  assign n1690 = ~n216 | n1151;
  assign n1691 = ~n216 | n994;
  assign n1692 = n1691 & n1690 & n1689 & n1688 & n1687 & n1686 & ~n760 & n762;
  assign n1693 = n1231 | n755;
  assign n1694 = n755 | n236;
  assign n1695 = n1151 | n755;
  assign n1696 = n1695 & n1694 & n1693 & n759;
  assign n1697 = n755 | n1232;
  assign n1698 = n1692 & (n942 | n755);
  assign n1699 = n1242 & n1176 & n1177 & n1763 & n1243 & n1304 & n2036 & n2008;
  assign n1700 = ~i_2_ & i_0_ & i_1_;
  assign n1701 = n524 & n773;
  assign n1702 = n1137 & n1515;
  assign n1703 = ~n123 & n1702;
  assign n1704 = n968 | n1703 | n960 | n975;
  assign n1705 = ~n110 | n237;
  assign n1706 = ~n110 | n1204;
  assign n1707 = ~n110 | n491;
  assign n1708 = ~n110 | n2293;
  assign n1709 = n1607 | n419;
  assign n1710 = n225 | n1129;
  assign n1711 = n225 | n643;
  assign n1712 = n1635 | n225;
  assign n1713 = n225 | n1208;
  assign n1714 = n1713 & n1712 & n1711 & n1710 & n793 & n398 & ~n219 & n270;
  assign n1715 = n231 | ~n818;
  assign n1716 = ~n818 | n1123;
  assign n1717 = ~n818 | n1635;
  assign n1718 = n294 & (n397 | ~n818);
  assign n1719 = n1718 & n1717 & n1715 & n1716;
  assign n1720 = n1762 | n419;
  assign n1721 = n728 | n850;
  assign n1722 = n1401 | n850;
  assign n1723 = n1722 & n1721 & n1720 & n823 & ~n821 & ~n822;
  assign n1724 = n225 | n1280;
  assign n1725 = n1634 | n225;
  assign n1726 = n235 | ~n818;
  assign n1727 = n225 | n1133;
  assign n1728 = n1404 & n1403 & n1320;
  assign n1729 = n2009 & n1719 & n1178 & ~n820 & ~n817 & ~n816 & n357 & n814;
  assign n1730 = n2295 | n419;
  assign n1731 = n2166 | n419;
  assign n1732 = n2294 | n419;
  assign n1733 = n349 | n232;
  assign n1734 = n2076 & n1506 & n1808;
  assign n1735 = n2156 & n1684 & n1550 & n1389 & n1239 & n1174 & ~n214 & n470;
  assign n1736 = n1505 & n1733 & n1732 & n1492 & n1730 & n1731 & n1734 & n1735;
  assign n1737 = n1762 | n796;
  assign n1738 = n1737 & n1487 & ~n113 & ~n808;
  assign n1739 = n225 | n572;
  assign n1740 = n796 | n572;
  assign n1741 = n225 | n237;
  assign n1742 = n469 | n1130;
  assign n1743 = n1494 & n1830 & n2029 & n1999;
  assign n1744 = n721 & n599 & n783 & n128 & n999 & n838 & n1570 & n2177;
  assign n1745 = n1246 & n2024 & n1502 & n1794 & n2026 & n1248 & n2176 & n2175;
  assign n1746 = n1743 & n1742 & n1345 & n1285 & n1740 & n1741 & n1744 & n1745;
  assign n1747 = n241 | n477;
  assign n1748 = ~n818 | n1214;
  assign n1749 = n780 | ~n818;
  assign n1750 = n225 | n244;
  assign n1751 = n225 | n990;
  assign n1752 = n225 | n1281;
  assign n1753 = n225 | n652;
  assign n1754 = n225 | n345;
  assign n1755 = n699 & n374;
  assign n1756 = n349 | n530;
  assign n1757 = n349 | n1281;
  assign n1758 = n1979 & n1940 & n1824 & n1423 & ~n108 & n1371;
  assign n1759 = n1497 & n1908 & n1252 & n1182 & n1251 & n2200 & n2023 & n2199;
  assign n1760 = n2203 & n891 & n997 & n129 & n531 & n1557 & n2204 & n2202;
  assign n1761 = n1760 & n1759 & n1758 & n1757 & n1756 & n1412 & ~n109 & n1365;
  assign n1762 = n628 & n723;
  assign n1763 = n755 | n776;
  assign n1764 = n1762 | n456;
  assign n1765 = n2225 & n757 & n2144 & n1009 & n2226 & n2159;
  assign n1766 = n1676 & n1720 & n672 & n1764 & n1763 & n1737 & n601 & n1765;
  assign n1767 = n225 | n1227;
  assign n1768 = n1231 | n225;
  assign n1769 = ~n220 & n1157;
  assign n1770 = ~n925 | n970;
  assign n1771 = ~n925 | n1151;
  assign n1772 = ~n925 | n1121;
  assign n1773 = (n1612 | n419) & (n456 | n496);
  assign n1774 = ~n923 & (n469 | (n572 & n1685));
  assign n1775 = n1836 & n1469 & n1451 & n1343 & n1287 & ~n119 & n1236;
  assign n1776 = n575 & n1563 & n1223 & n814 & n1592 & n1696;
  assign n1777 = n906 & n1746 & n1736 & n998 & n1766 & n922;
  assign n1778 = n2229 & n2228 & n1997 & n1725 & n1499 & n1427 & ~n113 & n1184;
  assign n1779 = n1778 & n1777 & n1776 & n1775 & n1774 & n1773 & ~n924 & n1148;
  assign n1780 = n747 & n610 & n740;
  assign n1781 = n543 & n1262 & n1354;
  assign n1782 = ~n1512 & n143 & ~n1084;
  assign n1783 = ~n652 & n1782;
  assign n1784 = ~n1045 & n1782;
  assign n1785 = ~n970 & n1782;
  assign n1786 = ~n970 & n1529;
  assign n1787 = ~n558 & n670;
  assign n1788 = ~n123 & n1518;
  assign n1789 = ~n123 & n1530;
  assign n1790 = ~n173 & ~n1119;
  assign n1791 = ~n539 | n2292;
  assign n1792 = n2292 | n796;
  assign n1793 = ~n539 | n1762;
  assign n1794 = n622 | n796;
  assign n1795 = ~n539 | n615;
  assign n1796 = n2297 | n796;
  assign n1797 = n2193 & n2200 & n2213 & n1004 & n2231 & n2236;
  assign n1798 = n1740 & n1795 & n1794 & n1793 & n1791 & n1792 & n1796 & n1797;
  assign n1799 = n2297 | n850;
  assign n1800 = n419 | n572;
  assign n1801 = n622 | n850;
  assign n1802 = n850 | n615;
  assign n1803 = n1762 | n850;
  assign n1804 = n2292 | n419;
  assign n1805 = n412 & n397 & n401;
  assign n1806 = n1340 & n1309 & n535;
  assign n1807 = ~n381 & ~n679;
  assign n1808 = n469 | n232;
  assign n1809 = n469 | n236;
  assign n1810 = n469 | n1149;
  assign n1811 = n1810 & n1808 & n1809;
  assign n1812 = n469 | n237;
  assign n1813 = ~n368 | n1127;
  assign n1814 = n469 | n1127;
  assign n1815 = n469 | n781;
  assign n1816 = n237 | ~n368;
  assign n1817 = n469 | n1261;
  assign n1818 = ~n368 | n1149;
  assign n1819 = ~n368 | n781;
  assign n1820 = ~n368 | n1124;
  assign n1821 = n469 | n1262;
  assign n1822 = n469 | n530;
  assign n1823 = ~n368 | n1045;
  assign n1824 = n469 | n652;
  assign n1825 = ~n368 | n515;
  assign n1826 = n469 | n1230;
  assign n1827 = ~n368 | n1230;
  assign n1828 = n469 | n1226;
  assign n1829 = n1828 & n1827 & n1826 & n1825 & n1823 & n1824;
  assign n1830 = n469 | n1209;
  assign n1831 = ~n368 | n1226;
  assign n1832 = ~n368 | n643;
  assign n1833 = ~n368 | n1214;
  assign n1834 = ~n368 | n1211;
  assign n1835 = ~n368 | n1207;
  assign n1836 = n469 | n970;
  assign n1837 = ~n368 | n1338;
  assign n1838 = n469 | n1340;
  assign n1839 = ~n368 | n1209;
  assign n1840 = n469 | n515;
  assign n1841 = n469 | n1214;
  assign n1842 = n1232 | n684;
  assign n1843 = n1842 & (n302 | n1232);
  assign n1844 = n456 | n1340;
  assign n1845 = n1232 | n1161;
  assign n1846 = n225 | n726;
  assign n1847 = n405 | n1261;
  assign n1848 = n405 | n1262;
  assign n1849 = n349 | n235;
  assign n1850 = n349 | n1153;
  assign n1851 = ~n430 | n1230;
  assign n1852 = ~n430 | n970;
  assign n1853 = ~n430 | n1209;
  assign n1854 = ~n430 | n1214;
  assign n1855 = n349 | n1230;
  assign n1856 = n349 | n970;
  assign n1857 = n469 | n1309;
  assign n1858 = ~n368 | n1224;
  assign n1859 = ~n368 | n1198;
  assign n1860 = n226 | ~n368;
  assign n1861 = n469 | n484;
  assign n1862 = n225 | n232;
  assign n1863 = ~n818 | n1127;
  assign n1864 = n225 | n346;
  assign n1865 = n225 | n530;
  assign n1866 = n225 | n1261;
  assign n1867 = n225 | n1262;
  assign n1868 = ~n818 | n1124;
  assign n1869 = ~n818 | n1136;
  assign n1870 = n236 | ~n818;
  assign n1871 = n237 | ~n818;
  assign n1872 = ~n220 | n727;
  assign n1873 = ~n220 | n1212;
  assign n1874 = ~n220 | n1225;
  assign n1875 = n456 | n1135;
  assign n1876 = ~n220 | n244;
  assign n1877 = ~n220 | n1150;
  assign n1878 = n456 | n1354;
  assign n1879 = ~n220 | n1202;
  assign n1880 = ~n220 | n532;
  assign n1881 = ~n220 | n1097;
  assign n1882 = n456 | n532;
  assign n1883 = n469 | n1150;
  assign n1884 = n469 | n1229;
  assign n1885 = ~n368 | n1150;
  assign n1886 = n1885 & n1883 & n1884;
  assign n1887 = n469 | n1225;
  assign n1888 = n244 | ~n368;
  assign n1889 = ~n368 | n1202;
  assign n1890 = ~n368 | n1215;
  assign n1891 = ~n368 | n1212;
  assign n1892 = ~n368 | n1229;
  assign n1893 = n469 | n1135;
  assign n1894 = n469 | n244;
  assign n1895 = n469 | n1202;
  assign n1896 = n469 | n1354;
  assign n1897 = ~n368 | n1135;
  assign n1898 = ~n368 | n990;
  assign n1899 = ~n368 | n780;
  assign n1900 = ~n368 | n1125;
  assign n1901 = n469 | n304;
  assign n1902 = n304 | ~n368;
  assign n1903 = n469 | n305;
  assign n1904 = n1903 & n1902 & n1901 & n1900 & n1898 & n1899;
  assign n1905 = ~n368 | n1129;
  assign n1906 = ~n368 | n1130;
  assign n1907 = n469 | n780;
  assign n1908 = n469 | n1281;
  assign n1909 = n469 | n543;
  assign n1910 = ~n368 | n1121;
  assign n1911 = n305 | ~n368;
  assign n1912 = ~n368 | n1281;
  assign n1913 = n405 | n532;
  assign n1914 = n1667 & n1913 & n694;
  assign n1915 = n243 | n532;
  assign n1916 = n593 & n583 & n1580 & n1543 & n1615 & n597;
  assign n1917 = ~n818 | n1110;
  assign n1918 = n1916 & n1917 & n1558 & n1555 & n1554 & n1544;
  assign n1919 = n1750 & (~n679 | (n1135 & n1150));
  assign n1920 = (~n220 | n1354) & (~n815 | n1353);
  assign n1921 = n1920 & (~n430 | n727);
  assign n1922 = ~n220 | n1229;
  assign n1923 = ~n220 | n1045;
  assign n1924 = ~n220 | n515;
  assign n1925 = ~n220 | n1211;
  assign n1926 = n456 | n515;
  assign n1927 = n405 | n1338;
  assign n1928 = n1683 & n1597 & n716 & n1927 & n1640 & n1608;
  assign n1929 = ~n368 | n1339;
  assign n1930 = n1929 & n1576 & n1569;
  assign n1931 = n1623 & n1556 & n1578 & n1562 & n1770 & n1748;
  assign n1932 = ~n220 | n1230;
  assign n1933 = (~n815 | n1338) & (n302 | n1339);
  assign n1934 = (n349 | n1207) & (~n220 | n1340);
  assign n1935 = n225 | n1308;
  assign n1936 = ~n220 | n1219;
  assign n1937 = ~n220 | n1224;
  assign n1938 = n456 | n1307;
  assign n1939 = n349 | n1198;
  assign n1940 = n349 | n345;
  assign n1941 = ~n430 | n1198;
  assign n1942 = n349 | n1208;
  assign n1943 = n349 | n1224;
  assign n1944 = ~n430 | n1204;
  assign n1945 = n1582 & n578 & n1593;
  assign n1946 = n243 | n1219;
  assign n1947 = n243 | n231;
  assign n1948 = n349 | n231;
  assign n1949 = n1948 & n1947 & n1946 & n1679 & n714 & n702 & n592 & n1945;
  assign n1950 = n1666 & n1653 & n690 & n1658 & n1661;
  assign n1951 = n243 | n1307;
  assign n1952 = n243 | n1198;
  assign n1953 = n1754 & (~n763 | (n1227 & n1308));
  assign n1954 = n1315 & (~n679 | (n1224 & n1228));
  assign n1955 = ~n220 | n1228;
  assign n1956 = ~n220 | n1046;
  assign n1957 = ~n220 | n305;
  assign n1958 = n456 | n525;
  assign n1959 = n349 | n1129;
  assign n1960 = ~n430 | n780;
  assign n1961 = ~n430 | n1125;
  assign n1962 = n349 | n1130;
  assign n1963 = n349 | n305;
  assign n1964 = n469 | n1280;
  assign n1965 = n225 | n238;
  assign n1966 = n405 | n543;
  assign n1967 = n243 | n525;
  assign n1968 = n1967 & n1564 & n581 & n1599;
  assign n1969 = n243 | n1046;
  assign n1970 = n405 | n525;
  assign n1971 = n1542 & n1553 & n1622 & n1577;
  assign n1972 = (n1152 | n1281) & (n306 | ~n679);
  assign n1973 = (n302 | n1280) & (~n212 | n780);
  assign n1974 = (~n818 | n1121) & (n349 | n1125);
  assign n1975 = ~n220 | n1153;
  assign n1976 = n456 | n781;
  assign n1977 = ~n220 | n1124;
  assign n1978 = ~n430 | n1124;
  assign n1979 = n349 | n346;
  assign n1980 = n349 | n781;
  assign n1981 = n237 | ~n430;
  assign n1982 = n731 & n574 & n1581 & n1609 & n1680 & n713;
  assign n1983 = n243 | n1123;
  assign n1984 = n232 | n243;
  assign n1985 = n405 | n1124;
  assign n1986 = n1660 & n1659 & n1985 & n1983 & n1984;
  assign n1987 = n1118 | n243;
  assign n1988 = n405 | n1136;
  assign n1989 = n1988 & n691 & n692 & n1987 & n1650 & n1652;
  assign n1990 = n243 | n1136;
  assign n1991 = ~n271 & ~n421;
  assign n1992 = n419 & n796;
  assign n1993 = (n1991 | n1123) & (n1992 | n1153);
  assign n1994 = ~n430 & ~n539;
  assign n1995 = n1993 & (n1994 | n781);
  assign n1996 = (n243 | n530) & (~n220 | n1262);
  assign n1997 = n1231 | n796;
  assign n1998 = ~n539 | n1231;
  assign n1999 = n419 | n1205;
  assign n2000 = n419 | n269;
  assign n2001 = n268 | n850;
  assign n2002 = n1395 | n850;
  assign n2003 = n472 & n468 & n1539;
  assign n2004 = ~n430 | n1205;
  assign n2005 = n349 | n1205;
  assign n2006 = n695 & n2005 & n2004 & n137 & n753 & n1693 & n1644 & n414;
  assign n2007 = ~n368 | n1197;
  assign n2008 = ~n216 | n1806;
  assign n2009 = ~n818 | n1401;
  assign n2010 = n456 & n1164;
  assign n2011 = n302 & n1156;
  assign n2012 = ~n679 & n1164;
  assign n2013 = (n2011 | n1199) & (n2012 | n1227);
  assign n2014 = ~n216 & n1162;
  assign n2015 = n1168 & ~n1053 & n225 & ~n539;
  assign n2016 = (n1205 | n2015) & (n226 | ~n381);
  assign n2017 = (n268 | n405) & (n316 | ~n421);
  assign n2018 = (n1164 | n1214) & (n1156 | n1232);
  assign n2019 = ~n430 | n726;
  assign n2020 = n1237 & n266 & n656 & n1245 & n1260 & n1014 & n270 & n2019;
  assign n2021 = n570 | n796;
  assign n2022 = ~n539 | n738;
  assign n2023 = n738 | n796;
  assign n2024 = n1396 | n796;
  assign n2025 = ~n218 | n796;
  assign n2026 = n1116 | n796;
  assign n2027 = n241 | n894;
  assign n2028 = n242 & n894;
  assign n2029 = n1116 | n419;
  assign n2030 = n419 | n570;
  assign n2031 = n355 | n419;
  assign n2032 = ~n218 | n850;
  assign n2033 = n1396 | n850;
  assign n2034 = ~n368 | n988;
  assign n2035 = n1588 & n1590 & n2034;
  assign n2036 = ~n216 | n1781;
  assign n2037 = ~n430 | n1116;
  assign n2038 = n1664 & n2037 & n136 & n1695 & n2036 & n754 & n696 & n1648;
  assign n2039 = ~n818 | n1116;
  assign n2040 = (n248 | n1115) & (n2014 | n1144);
  assign n2041 = (n1125 | n2010) & (n239 | ~n273);
  assign n2042 = (~n250 | n653) & (n1116 | n2015);
  assign n2043 = (n994 | n1157) & (~n381 | n1124);
  assign n2044 = (n238 | n1156) & (~n218 | n405);
  assign n2045 = n1172 & (~n220 | n1118);
  assign n2046 = n1180 & n1187 & n1195 & n139;
  assign n2047 = n1717 & n1712 & ~n117 & n715;
  assign n2048 = ~n380 & (n2010 | (n1209 & n1390));
  assign n2049 = ~n383 & (~n273 | (n648 & n1391));
  assign n2050 = ~n384 & (~n212 | (n352 & n1392));
  assign n2051 = ~n386 & (~n818 | (n226 & ~n879));
  assign n2052 = ~n1053 & n1393;
  assign n2053 = (n378 | n225) & (n1573 | n2052);
  assign n2054 = ~n212 | n372;
  assign n2055 = (n376 | n456) & (n230 | ~n679);
  assign n2056 = (~n539 | n842) & (n1635 | n1991);
  assign n2057 = ~n220 & n419;
  assign n2058 = (n653 | n2057) & (n1156 | n1005);
  assign n2059 = ~n271 & n1398;
  assign n2060 = (n1164 | n1391) & (n375 | n2059);
  assign n2061 = ~n271 & ~n501;
  assign n2062 = (n233 | ~n430) & (n234 | n2061);
  assign n2063 = n1399 & n225 & n1398;
  assign n2064 = n1400 & n456 & n1399;
  assign n2065 = (n1574 | n2063) & (n1537 | n2064);
  assign n2066 = ~n216 & ~n925;
  assign n2067 = (n1231 | n2066) & (n1463 | n1213);
  assign n2068 = n740 | n2132;
  assign n2069 = (~n271 | n726) & (~n815 | n1151);
  assign n2070 = (~n110 | n530) & (n1158 | n1227);
  assign n2071 = n1425 & n423 & n1442 & n534 & n344 & n542 & n1416 & n1035;
  assign n2072 = n2291 | n796;
  assign n2073 = ~n539 | n779;
  assign n2074 = n779 | n796;
  assign n2075 = n481 | n894;
  assign n2076 = n469 | n725;
  assign n2077 = n1755 | n456;
  assign n2078 = ~n368 | n1466;
  assign n2079 = ~n368 | n756;
  assign n2080 = ~n368 | n632;
  assign n2081 = ~n368 | n628;
  assign n2082 = ~n368 | n642;
  assign n2083 = n469 | n636;
  assign n2084 = ~n368 | n1465;
  assign n2085 = n2084 & (~n764 | (~n763 & n1161));
  assign n2086 = (n1483 | n1468) & (n2066 | n756);
  assign n2087 = n850 & n796;
  assign n2088 = n419 & ~n271 & ~n368;
  assign n2089 = n2087 | n232;
  assign n2090 = (~n212 | n781) & (n1161 | n1262);
  assign n2091 = n1220 & n1145;
  assign n2092 = ~n763 & n1393;
  assign n2093 = ~n213 & (n2092 | (n1262 & n1309));
  assign n2094 = ~n499 & (n491 | (n225 & n1477));
  assign n2095 = ~n500 & (n699 | (n405 & n1478));
  assign n2096 = ~n679 & n1159;
  assign n2097 = (n1805 | n489) & (n2096 | n498);
  assign n2098 = (n492 | ~n1053) & (n490 | n1468);
  assign n2099 = ~n763 & n1162;
  assign n2100 = ~n501 & n796;
  assign n2101 = (n2100 | n1124) & (n2087 | n781);
  assign n2102 = n755 & n1482;
  assign n2103 = (n1769 | n945) & (n2102 | n1228);
  assign n2104 = n2101 & n2103 & (n1165 | n1153);
  assign n2105 = n1164 & n1483;
  assign n2106 = (~n379 | n412) & (n1149 | n2105);
  assign n2107 = n1165 & n796 & n488;
  assign n2108 = (~n273 | n485) & (n1224 | n2107);
  assign n2109 = (n463 | n1400) & (~n385 | n1398);
  assign n2110 = (n243 | n401) & (n484 | ~n679);
  assign n2111 = (~n368 | n589) & (n755 | n756);
  assign n2112 = n494 & n2111 & (~n539 | n1136);
  assign n2113 = n1495 & n1013 & n140 & n476 & n450 & n1511 & n1488 & n1485;
  assign n2114 = n416 & n413 & n409 & n406 & n398 & n402 & n429 & n440;
  assign n2115 = n1385 & (n456 | (n1390 & n1280));
  assign n2116 = (n1134 | n2057) & (n535 | ~n546);
  assign n2117 = (~n815 | n1150) & (n1229 | n2066);
  assign n2118 = ~n212 | n1215;
  assign n2119 = n1221 & (n1164 | (n1390 & n1353));
  assign n2120 = n2119 & (n243 | (n653 & n990));
  assign n2121 = (n229 | n2061) & (n1482 | n727);
  assign n2122 = n247 & n1519;
  assign n2123 = (n2122 | n346) & (n2052 | n1143);
  assign n2124 = (~n503 | n1516) & (n232 | n1462);
  assign n2125 = (n1202 | n2012) & (~n818 | n1392);
  assign n2126 = (~n421 | n1105) & (n1280 | n2059);
  assign n2127 = n1398 & n456 & n684;
  assign n2128 = n2125 & n2126 & (n2127 | n1261);
  assign n2129 = (n1519 | n1127) & (n2063 | n245);
  assign n2130 = (n2102 | n1229) & (n2064 | n570);
  assign n2131 = n1098 | n1154;
  assign n2132 = ~n925 & n755 & ~n679 & ~n368 & n456;
  assign n2133 = (n994 | n2132) & (~n879 | n1152);
  assign n2134 = (n2092 | n535) & (n1156 | n1781);
  assign n2135 = ~n368 | n651;
  assign n2136 = n2289 | n469;
  assign n2137 = n651 | n469;
  assign n2138 = ~n368 | n1612;
  assign n2139 = n608 | n469;
  assign n2140 = n469 | n776;
  assign n2141 = n536 & n544 & n666 & n1589 & n606 & n612 & n476 & n448;
  assign n2142 = ~n220 | n645;
  assign n2143 = n456 | n572;
  assign n2144 = n620 | n456;
  assign n2145 = n1612 | n456;
  assign n2146 = n2289 | n456;
  assign n2147 = n1442 & n1330 & n327 & n1552 & n649 & n1511;
  assign n2148 = n1150 & n304;
  assign n2149 = n993 | n349;
  assign n2150 = n349 | n613;
  assign n2151 = ~n430 | n1634;
  assign n2152 = (~n421 | n741) & (~n430 | n739);
  assign n2153 = n266 & (~n142 | n261);
  assign n2154 = n622 | n243;
  assign n2155 = n1358 & n1848 & n1319 & n1966 & n1355 & n358 & n1847 & n1318;
  assign n2156 = n2166 | n405;
  assign n2157 = n1612 | n405;
  assign n2158 = n2292 | n405;
  assign n2159 = n620 | n405;
  assign n2160 = ~n277 | n748;
  assign n2161 = ~n381 | n1614;
  assign n2162 = n1936 & n1956;
  assign n2163 = n813 | ~n818;
  assign n2164 = n1925 & (n615 | (~n379 & ~n818));
  assign n2165 = n2166 | n850;
  assign n2166 = n1197 & n725 & n988;
  assign n2167 = (~n379 | n725) & (~n818 | n2166);
  assign n2168 = n2135 & n1981 & n1944 & n1978 & n1364 & n1415 & n1421 & n1816;
  assign n2169 = n1283 & n1341 & n2039 & n1235 & n1434 & n1977 & n1501 & n785;
  assign n2170 = n1801 & n1871 & n1313 & n1868 & n1288 & n1917 & n2002 & n2033;
  assign n2171 = ~n379 & n1152;
  assign n2172 = n242 & ~n709;
  assign n2173 = (~n368 | n572) & (~n818 | n1395);
  assign n2174 = n1504 & n1173;
  assign n2175 = n1812 & n2143 & n1962 & n2137 & n1410 & n1637 & n1238 & n2174;
  assign n2176 = n2072 & n2075 & n1475;
  assign n2177 = n1800 & (n349 | n632);
  assign n2178 = ~n220 | n825;
  assign n2179 = n453 & n647 & n1572 & n1601 & n735 & n576 & n1223 & n2178;
  assign n2180 = n1903 & n1887 & n2146 & n1814 & n1893 & n1815 & n1828;
  assign n2181 = n1476 & n1265 & n1407 & n1959 & n263 & n1408 & n786;
  assign n2182 = n1350 & n1804 & n1862 & n1431 & n1437 & n1976 & n2030;
  assign n2183 = (n1537 | n405) & (n469 | n463);
  assign n2184 = n464 & (n478 | n894);
  assign n2185 = n1874 & n1957 & n1937 & n2073 & n1418 & n1813;
  assign n2186 = n1348 & n1328 & n1436 & n1819 & n1349 & n1295;
  assign n2187 = n2082 & n1443 & n1831 & n2032 & n1832 & n1905 & n2186;
  assign n2188 = ~n867 & (n478 | (n242 & n477));
  assign n2189 = (n1994 | n781) & (n1400 | n792);
  assign n2190 = n2189 & (n1537 | n1477);
  assign n2191 = (n352 | n850) & (n353 | ~n1051);
  assign n2192 = n1438 & n1958 & n1938 & n1277 & n1939 & n1369;
  assign n2193 = n796 | n613;
  assign n2194 = n1140 & n2150 & n2027 & n2193 & n1796 & n1169 & n2192;
  assign n2195 = n2149 & n1428 & n1342 & n1286 & ~n116 & n1272;
  assign n2196 = n993 | n419;
  assign n2197 = (n405 | n589) & (n349 | n412);
  assign n2198 = n1589 & n637 & n413;
  assign n2199 = n1170 & n1413 & n1142;
  assign n2200 = n624 | n796;
  assign n2201 = n1256 & n1490 & n1193;
  assign n2202 = n1864 & n1861 & n1454 & n1894 & n2077 & n1822 & n1865 & n2201;
  assign n2203 = n1472 & n1895 & n1381;
  assign n2204 = (n895 | n265) & (n469 | n699);
  assign n2205 = n1859 & n1373 & n1294 & n1327 & n1372 & n1439 & n1890;
  assign n2206 = ~n818 | n993;
  assign n2207 = n1880 & n2206 & n1270 & n1079 & n1402 & n1924;
  assign n2208 = n2054 & n1491 & n1255 & n1192;
  assign n2209 = ~n213 & (n613 | (n850 & n1152));
  assign n2210 = n2209 & (~n539 | (n589 & n688));
  assign n2211 = n636 & n897;
  assign n2212 = n1889 & n1823 & n1370 & n1888 & n1422 & n1898 & n1141;
  assign n2213 = ~n539 | n624;
  assign n2214 = n1923 & n1290 & n1268 & n1324 & n1879 & n1269 & n2078;
  assign n2215 = n1234 & (n1574 | (~n539 & n850));
  assign n2216 = ~n907 & (~n368 | (n874 & n1755));
  assign n2217 = (n1400 | n1548) & (n1397 | n1281);
  assign n2218 = (~n277 | n746) & (~n212 | n528);
  assign n2219 = (n1152 | n738) & (n1164 | n747);
  assign n2220 = (n374 | ~n1051) & (n652 | n1398);
  assign n2221 = n265 | n242;
  assign n2222 = n2211 | n349;
  assign n2223 = n1136 & n236 & n397 & n1215 & n532 & n1307;
  assign n2224 = n1762 & ~n918 & n845 & n780 & n636 & n667;
  assign n2225 = (n1992 | n615) & (n225 | n613);
  assign n2226 = n620 | n419;
  assign n2227 = n2157 & n1948 & n1826 & n1362 & n1331 & n1275;
  assign n2228 = n1419 & n1901 & n1809 & n2145 & n1810 & n1883 & n1884 & n2227;
  assign n2229 = n1363 & n1332 & n1297 & n1856 & n1855 & n1298;
  assign n2230 = n1902 & n1417 & n1892 & n1827 & n731 & n2138 & n1885 & n1818;
  assign n2231 = ~n539 | n620;
  assign n2232 = n1185 & n1998 & n1300 & n1852 & n1500 & n828 & n2231;
  assign n2233 = (~n709 | n1112) & (~n220 | n776);
  assign n2234 = n2233 & n453 & n1541 & n1633 & n1585 & n621;
  assign n2235 = n1509 & n1867 & n1866 & n1821 & n1878 & n1549;
  assign n2236 = n796 | ~n1027;
  assign n2237 = n1571 & n1333 & n1817 & n830 & n1420 & n2139 & n2236 & n2235;
  assign n2238 = n1470 & n1838 & n1447 & n1190 & n1453 & n1380;
  assign n2239 = (n946 | n469) & (n685 | n684);
  assign n2240 = n1781 & ~n764 & n944;
  assign n2241 = (n2240 | n1161) & (n488 | n941);
  assign n2242 = n1180 & n1245 & (n992 | n796);
  assign n2243 = ~n979 | n982;
  assign n2244 = (~n172 | ~n1119) & (n1513 | n1790);
  assign n2245 = n516 & n969;
  assign n2246 = (n1083 | n122) & (n2245 | n990);
  assign n2247 = (n122 | ~n1119) & (n304 | n2245);
  assign n2248 = (n1230 | n2245) & (n122 | ~n173);
  assign n2249 = n1083 & n1790;
  assign n2250 = ~n159 & (~n222 | n1512 | n2249);
  assign n2251 = n1935 & n1917 & n2206;
  assign n2252 = n361 & n1965 & (n996 | n225);
  assign n2253 = (n610 | ~n815) & (~n818 | n991);
  assign n2254 = ~n1028 & (~n501 | (~n385 & n1780));
  assign n2255 = n2254 & (n1026 | n850);
  assign n2256 = (n2066 | n1230) & (n247 | n652);
  assign n2257 = ~n1050 & (n2092 | (n543 & n1340));
  assign n2258 = ~n1055 & (n990 | (~n381 & n1393));
  assign n2259 = (n1160 | n945) & (n2099 | n985);
  assign n2260 = (~n503 | n1047) & (n1478 | n1481);
  assign n2261 = (n615 | n1043) & (~n281 | n1465);
  assign n2262 = (~n815 | n1480) & (n645 | n1155);
  assign n2263 = (n1338 | n2100) & (~n1027 | n1477);
  assign n2264 = (n726 | n1165) & (n524 | ~n679);
  assign n2265 = (n1769 | n605) & (n2102 | n1230);
  assign n2266 = (n2105 | n304) & (n2066 | n776);
  assign n2267 = (n247 | n1466) & (n622 | n419);
  assign n2268 = (~n381 | n401) & (~n421 | n628);
  assign n2269 = (n488 | n1467) & (n1164 | n1111);
  assign n2270 = (n1398 | n652) & (n1156 | n1133);
  assign n2271 = (n456 | n632) & (~n110 | n463);
  assign n2272 = n796 | n1045;
  assign n2273 = n2270 & n2271 & n2272 & n450 & n554 & n526;
  assign n2274 = n1146 & (n1156 | (n1806 & n1134));
  assign n2275 = n2274 & (n484 | (n225 & ~n421));
  assign n2276 = ~n1065 & (n244 | (n1393 & n1807));
  assign n2277 = (n228 | n2061) & (~n110 | n778);
  assign n2278 = n2277 & (n1394 | n2059);
  assign n2279 = (n2122 | n345) & (n2052 | n1217);
  assign n2280 = ~n1066 & ~n1067 & (n1110 | n2100);
  assign n2281 = (n2127 | n1308) & (n1519 | n1208);
  assign n2282 = (n2063 | n1216) & (n2105 | n1150);
  assign n2283 = (n2064 | n269) & (n247 | n231);
  assign n2284 = (n2132 | n1199) & (n1210 | n243);
  assign n2285 = (~n503 | n1097) & (n1354 | n2092);
  assign n2286 = (n1135 | n2107) & (~n381 | n1202);
  assign n2287 = (~n430 | n1045) & (n405 | n652);
  assign n2288 = i_2_ | ~i_0_ | i_1_;
  assign n2289 = n610 & n1537;
  assign n2290 = n226 & n1110 & n1111;
  assign n2291 = n401 & n237 & n1204;
  assign n2292 = n642 & n353;
  assign n2293 = n226 & n401 & n1124;
  assign n2294 = n1123 & n1098;
  assign n2295 = n1219 & n1213;
  assign n2296 = n1198 & n459;
  assign n2297 = n636 & n348;
  assign n2298 = ~n879 & n1307;
endmodule


