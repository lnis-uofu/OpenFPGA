*****************************
*     FPGA SPICE Netlist    *
* Description: Connection Block Y-channel  [0][1] in FPGA *
*    Author: Xifan TANG     *
* Organization: EPFL/IC/LSI *
* Date: Thu Nov 15 14:26:08 2018
 *
*****************************
.subckt cby[0][1] 
+ chany[0][1]_midout[0] 
+ chany[0][1]_midout[1] 
+ chany[0][1]_midout[2] 
+ chany[0][1]_midout[3] 
+ chany[0][1]_midout[4] 
+ chany[0][1]_midout[5] 
+ chany[0][1]_midout[6] 
+ chany[0][1]_midout[7] 
+ chany[0][1]_midout[8] 
+ chany[0][1]_midout[9] 
+ chany[0][1]_midout[10] 
+ chany[0][1]_midout[11] 
+ chany[0][1]_midout[12] 
+ chany[0][1]_midout[13] 
+ chany[0][1]_midout[14] 
+ chany[0][1]_midout[15] 
+ chany[0][1]_midout[16] 
+ chany[0][1]_midout[17] 
+ chany[0][1]_midout[18] 
+ chany[0][1]_midout[19] 
+ chany[0][1]_midout[20] 
+ chany[0][1]_midout[21] 
+ chany[0][1]_midout[22] 
+ chany[0][1]_midout[23] 
+ chany[0][1]_midout[24] 
+ chany[0][1]_midout[25] 
+ chany[0][1]_midout[26] 
+ chany[0][1]_midout[27] 
+ chany[0][1]_midout[28] 
+ chany[0][1]_midout[29] 
+ chany[0][1]_midout[30] 
+ chany[0][1]_midout[31] 
+ chany[0][1]_midout[32] 
+ chany[0][1]_midout[33] 
+ chany[0][1]_midout[34] 
+ chany[0][1]_midout[35] 
+ chany[0][1]_midout[36] 
+ chany[0][1]_midout[37] 
+ chany[0][1]_midout[38] 
+ chany[0][1]_midout[39] 
+ chany[0][1]_midout[40] 
+ chany[0][1]_midout[41] 
+ chany[0][1]_midout[42] 
+ chany[0][1]_midout[43] 
+ chany[0][1]_midout[44] 
+ chany[0][1]_midout[45] 
+ chany[0][1]_midout[46] 
+ chany[0][1]_midout[47] 
+ chany[0][1]_midout[48] 
+ chany[0][1]_midout[49] 
+ chany[0][1]_midout[50] 
+ chany[0][1]_midout[51] 
+ chany[0][1]_midout[52] 
+ chany[0][1]_midout[53] 
+ chany[0][1]_midout[54] 
+ chany[0][1]_midout[55] 
+ chany[0][1]_midout[56] 
+ chany[0][1]_midout[57] 
+ chany[0][1]_midout[58] 
+ chany[0][1]_midout[59] 
+ chany[0][1]_midout[60] 
+ chany[0][1]_midout[61] 
+ chany[0][1]_midout[62] 
+ chany[0][1]_midout[63] 
+ chany[0][1]_midout[64] 
+ chany[0][1]_midout[65] 
+ chany[0][1]_midout[66] 
+ chany[0][1]_midout[67] 
+ chany[0][1]_midout[68] 
+ chany[0][1]_midout[69] 
+ chany[0][1]_midout[70] 
+ chany[0][1]_midout[71] 
+ chany[0][1]_midout[72] 
+ chany[0][1]_midout[73] 
+ chany[0][1]_midout[74] 
+ chany[0][1]_midout[75] 
+ chany[0][1]_midout[76] 
+ chany[0][1]_midout[77] 
+ chany[0][1]_midout[78] 
+ chany[0][1]_midout[79] 
+ chany[0][1]_midout[80] 
+ chany[0][1]_midout[81] 
+ chany[0][1]_midout[82] 
+ chany[0][1]_midout[83] 
+ chany[0][1]_midout[84] 
+ chany[0][1]_midout[85] 
+ chany[0][1]_midout[86] 
+ chany[0][1]_midout[87] 
+ chany[0][1]_midout[88] 
+ chany[0][1]_midout[89] 
+ chany[0][1]_midout[90] 
+ chany[0][1]_midout[91] 
+ chany[0][1]_midout[92] 
+ chany[0][1]_midout[93] 
+ chany[0][1]_midout[94] 
+ chany[0][1]_midout[95] 
+ chany[0][1]_midout[96] 
+ chany[0][1]_midout[97] 
+ chany[0][1]_midout[98] 
+ chany[0][1]_midout[99] 
+ grid[1][1]_pin[0][3][3] 
+ grid[1][1]_pin[0][3][7] 
+ grid[1][1]_pin[0][3][11] 
+ grid[1][1]_pin[0][3][15] 
+ grid[1][1]_pin[0][3][19] 
+ grid[1][1]_pin[0][3][23] 
+ grid[1][1]_pin[0][3][27] 
+ grid[1][1]_pin[0][3][31] 
+ grid[1][1]_pin[0][3][35] 
+ grid[1][1]_pin[0][3][39] 
+ grid[0][1]_pin[0][1][0] 
+ grid[0][1]_pin[0][1][2] 
+ grid[0][1]_pin[0][1][4] 
+ grid[0][1]_pin[0][1][6] 
+ grid[0][1]_pin[0][1][8] 
+ grid[0][1]_pin[0][1][10] 
+ grid[0][1]_pin[0][1][12] 
+ grid[0][1]_pin[0][1][14] 
+ svdd sgnd
Xmux_2level_tapbuf_size16[36] chany[0][1]_midout[0] chany[0][1]_midout[1] chany[0][1]_midout[12] chany[0][1]_midout[13] chany[0][1]_midout[24] chany[0][1]_midout[25] chany[0][1]_midout[38] chany[0][1]_midout[39] chany[0][1]_midout[50] chany[0][1]_midout[51] chany[0][1]_midout[62] chany[0][1]_midout[63] chany[0][1]_midout[74] chany[0][1]_midout[75] chany[0][1]_midout[88] chany[0][1]_midout[89] grid[1][1]_pin[0][3][3] sram[2370]->outb sram[2370]->out sram[2371]->out sram[2371]->outb sram[2372]->out sram[2372]->outb sram[2373]->out sram[2373]->outb sram[2374]->outb sram[2374]->out sram[2375]->out sram[2375]->outb sram[2376]->out sram[2376]->outb sram[2377]->out sram[2377]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[36], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2370] sram->in sram[2370]->out sram[2370]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2370]->out) 0
.nodeset V(sram[2370]->outb) vsp
Xsram[2371] sram->in sram[2371]->out sram[2371]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2371]->out) 0
.nodeset V(sram[2371]->outb) vsp
Xsram[2372] sram->in sram[2372]->out sram[2372]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2372]->out) 0
.nodeset V(sram[2372]->outb) vsp
Xsram[2373] sram->in sram[2373]->out sram[2373]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2373]->out) 0
.nodeset V(sram[2373]->outb) vsp
Xsram[2374] sram->in sram[2374]->out sram[2374]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2374]->out) 0
.nodeset V(sram[2374]->outb) vsp
Xsram[2375] sram->in sram[2375]->out sram[2375]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2375]->out) 0
.nodeset V(sram[2375]->outb) vsp
Xsram[2376] sram->in sram[2376]->out sram[2376]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2376]->out) 0
.nodeset V(sram[2376]->outb) vsp
Xsram[2377] sram->in sram[2377]->out sram[2377]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2377]->out) 0
.nodeset V(sram[2377]->outb) vsp
Xmux_2level_tapbuf_size16[37] chany[0][1]_midout[2] chany[0][1]_midout[3] chany[0][1]_midout[14] chany[0][1]_midout[15] chany[0][1]_midout[26] chany[0][1]_midout[27] chany[0][1]_midout[38] chany[0][1]_midout[39] chany[0][1]_midout[52] chany[0][1]_midout[53] chany[0][1]_midout[64] chany[0][1]_midout[65] chany[0][1]_midout[76] chany[0][1]_midout[77] chany[0][1]_midout[88] chany[0][1]_midout[89] grid[1][1]_pin[0][3][7] sram[2378]->outb sram[2378]->out sram[2379]->out sram[2379]->outb sram[2380]->out sram[2380]->outb sram[2381]->out sram[2381]->outb sram[2382]->outb sram[2382]->out sram[2383]->out sram[2383]->outb sram[2384]->out sram[2384]->outb sram[2385]->out sram[2385]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[37], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2378] sram->in sram[2378]->out sram[2378]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2378]->out) 0
.nodeset V(sram[2378]->outb) vsp
Xsram[2379] sram->in sram[2379]->out sram[2379]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2379]->out) 0
.nodeset V(sram[2379]->outb) vsp
Xsram[2380] sram->in sram[2380]->out sram[2380]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2380]->out) 0
.nodeset V(sram[2380]->outb) vsp
Xsram[2381] sram->in sram[2381]->out sram[2381]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2381]->out) 0
.nodeset V(sram[2381]->outb) vsp
Xsram[2382] sram->in sram[2382]->out sram[2382]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2382]->out) 0
.nodeset V(sram[2382]->outb) vsp
Xsram[2383] sram->in sram[2383]->out sram[2383]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2383]->out) 0
.nodeset V(sram[2383]->outb) vsp
Xsram[2384] sram->in sram[2384]->out sram[2384]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2384]->out) 0
.nodeset V(sram[2384]->outb) vsp
Xsram[2385] sram->in sram[2385]->out sram[2385]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2385]->out) 0
.nodeset V(sram[2385]->outb) vsp
Xmux_2level_tapbuf_size16[38] chany[0][1]_midout[2] chany[0][1]_midout[3] chany[0][1]_midout[14] chany[0][1]_midout[15] chany[0][1]_midout[28] chany[0][1]_midout[29] chany[0][1]_midout[40] chany[0][1]_midout[41] chany[0][1]_midout[52] chany[0][1]_midout[53] chany[0][1]_midout[64] chany[0][1]_midout[65] chany[0][1]_midout[78] chany[0][1]_midout[79] chany[0][1]_midout[90] chany[0][1]_midout[91] grid[1][1]_pin[0][3][11] sram[2386]->outb sram[2386]->out sram[2387]->out sram[2387]->outb sram[2388]->out sram[2388]->outb sram[2389]->out sram[2389]->outb sram[2390]->outb sram[2390]->out sram[2391]->out sram[2391]->outb sram[2392]->out sram[2392]->outb sram[2393]->out sram[2393]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[38], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2386] sram->in sram[2386]->out sram[2386]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2386]->out) 0
.nodeset V(sram[2386]->outb) vsp
Xsram[2387] sram->in sram[2387]->out sram[2387]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2387]->out) 0
.nodeset V(sram[2387]->outb) vsp
Xsram[2388] sram->in sram[2388]->out sram[2388]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2388]->out) 0
.nodeset V(sram[2388]->outb) vsp
Xsram[2389] sram->in sram[2389]->out sram[2389]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2389]->out) 0
.nodeset V(sram[2389]->outb) vsp
Xsram[2390] sram->in sram[2390]->out sram[2390]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2390]->out) 0
.nodeset V(sram[2390]->outb) vsp
Xsram[2391] sram->in sram[2391]->out sram[2391]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2391]->out) 0
.nodeset V(sram[2391]->outb) vsp
Xsram[2392] sram->in sram[2392]->out sram[2392]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2392]->out) 0
.nodeset V(sram[2392]->outb) vsp
Xsram[2393] sram->in sram[2393]->out sram[2393]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2393]->out) 0
.nodeset V(sram[2393]->outb) vsp
Xmux_2level_tapbuf_size16[39] chany[0][1]_midout[4] chany[0][1]_midout[5] chany[0][1]_midout[16] chany[0][1]_midout[17] chany[0][1]_midout[28] chany[0][1]_midout[29] chany[0][1]_midout[42] chany[0][1]_midout[43] chany[0][1]_midout[54] chany[0][1]_midout[55] chany[0][1]_midout[66] chany[0][1]_midout[67] chany[0][1]_midout[78] chany[0][1]_midout[79] chany[0][1]_midout[92] chany[0][1]_midout[93] grid[1][1]_pin[0][3][15] sram[2394]->outb sram[2394]->out sram[2395]->out sram[2395]->outb sram[2396]->out sram[2396]->outb sram[2397]->out sram[2397]->outb sram[2398]->outb sram[2398]->out sram[2399]->out sram[2399]->outb sram[2400]->out sram[2400]->outb sram[2401]->out sram[2401]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[39], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2394] sram->in sram[2394]->out sram[2394]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2394]->out) 0
.nodeset V(sram[2394]->outb) vsp
Xsram[2395] sram->in sram[2395]->out sram[2395]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2395]->out) 0
.nodeset V(sram[2395]->outb) vsp
Xsram[2396] sram->in sram[2396]->out sram[2396]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2396]->out) 0
.nodeset V(sram[2396]->outb) vsp
Xsram[2397] sram->in sram[2397]->out sram[2397]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2397]->out) 0
.nodeset V(sram[2397]->outb) vsp
Xsram[2398] sram->in sram[2398]->out sram[2398]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2398]->out) 0
.nodeset V(sram[2398]->outb) vsp
Xsram[2399] sram->in sram[2399]->out sram[2399]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2399]->out) 0
.nodeset V(sram[2399]->outb) vsp
Xsram[2400] sram->in sram[2400]->out sram[2400]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2400]->out) 0
.nodeset V(sram[2400]->outb) vsp
Xsram[2401] sram->in sram[2401]->out sram[2401]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2401]->out) 0
.nodeset V(sram[2401]->outb) vsp
Xmux_2level_tapbuf_size16[40] chany[0][1]_midout[4] chany[0][1]_midout[5] chany[0][1]_midout[18] chany[0][1]_midout[19] chany[0][1]_midout[30] chany[0][1]_midout[31] chany[0][1]_midout[42] chany[0][1]_midout[43] chany[0][1]_midout[54] chany[0][1]_midout[55] chany[0][1]_midout[68] chany[0][1]_midout[69] chany[0][1]_midout[80] chany[0][1]_midout[81] chany[0][1]_midout[92] chany[0][1]_midout[93] grid[1][1]_pin[0][3][19] sram[2402]->outb sram[2402]->out sram[2403]->out sram[2403]->outb sram[2404]->out sram[2404]->outb sram[2405]->out sram[2405]->outb sram[2406]->outb sram[2406]->out sram[2407]->out sram[2407]->outb sram[2408]->out sram[2408]->outb sram[2409]->out sram[2409]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[40], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2402] sram->in sram[2402]->out sram[2402]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2402]->out) 0
.nodeset V(sram[2402]->outb) vsp
Xsram[2403] sram->in sram[2403]->out sram[2403]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2403]->out) 0
.nodeset V(sram[2403]->outb) vsp
Xsram[2404] sram->in sram[2404]->out sram[2404]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2404]->out) 0
.nodeset V(sram[2404]->outb) vsp
Xsram[2405] sram->in sram[2405]->out sram[2405]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2405]->out) 0
.nodeset V(sram[2405]->outb) vsp
Xsram[2406] sram->in sram[2406]->out sram[2406]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2406]->out) 0
.nodeset V(sram[2406]->outb) vsp
Xsram[2407] sram->in sram[2407]->out sram[2407]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2407]->out) 0
.nodeset V(sram[2407]->outb) vsp
Xsram[2408] sram->in sram[2408]->out sram[2408]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2408]->out) 0
.nodeset V(sram[2408]->outb) vsp
Xsram[2409] sram->in sram[2409]->out sram[2409]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2409]->out) 0
.nodeset V(sram[2409]->outb) vsp
Xmux_2level_tapbuf_size16[41] chany[0][1]_midout[6] chany[0][1]_midout[7] chany[0][1]_midout[18] chany[0][1]_midout[19] chany[0][1]_midout[32] chany[0][1]_midout[33] chany[0][1]_midout[44] chany[0][1]_midout[45] chany[0][1]_midout[56] chany[0][1]_midout[57] chany[0][1]_midout[68] chany[0][1]_midout[69] chany[0][1]_midout[82] chany[0][1]_midout[83] chany[0][1]_midout[94] chany[0][1]_midout[95] grid[1][1]_pin[0][3][23] sram[2410]->outb sram[2410]->out sram[2411]->out sram[2411]->outb sram[2412]->out sram[2412]->outb sram[2413]->out sram[2413]->outb sram[2414]->outb sram[2414]->out sram[2415]->out sram[2415]->outb sram[2416]->out sram[2416]->outb sram[2417]->out sram[2417]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[41], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2410] sram->in sram[2410]->out sram[2410]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2410]->out) 0
.nodeset V(sram[2410]->outb) vsp
Xsram[2411] sram->in sram[2411]->out sram[2411]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2411]->out) 0
.nodeset V(sram[2411]->outb) vsp
Xsram[2412] sram->in sram[2412]->out sram[2412]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2412]->out) 0
.nodeset V(sram[2412]->outb) vsp
Xsram[2413] sram->in sram[2413]->out sram[2413]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2413]->out) 0
.nodeset V(sram[2413]->outb) vsp
Xsram[2414] sram->in sram[2414]->out sram[2414]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2414]->out) 0
.nodeset V(sram[2414]->outb) vsp
Xsram[2415] sram->in sram[2415]->out sram[2415]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2415]->out) 0
.nodeset V(sram[2415]->outb) vsp
Xsram[2416] sram->in sram[2416]->out sram[2416]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2416]->out) 0
.nodeset V(sram[2416]->outb) vsp
Xsram[2417] sram->in sram[2417]->out sram[2417]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2417]->out) 0
.nodeset V(sram[2417]->outb) vsp
Xmux_2level_tapbuf_size16[42] chany[0][1]_midout[8] chany[0][1]_midout[9] chany[0][1]_midout[20] chany[0][1]_midout[21] chany[0][1]_midout[32] chany[0][1]_midout[33] chany[0][1]_midout[44] chany[0][1]_midout[45] chany[0][1]_midout[58] chany[0][1]_midout[59] chany[0][1]_midout[70] chany[0][1]_midout[71] chany[0][1]_midout[82] chany[0][1]_midout[83] chany[0][1]_midout[94] chany[0][1]_midout[95] grid[1][1]_pin[0][3][27] sram[2418]->outb sram[2418]->out sram[2419]->out sram[2419]->outb sram[2420]->out sram[2420]->outb sram[2421]->out sram[2421]->outb sram[2422]->outb sram[2422]->out sram[2423]->out sram[2423]->outb sram[2424]->out sram[2424]->outb sram[2425]->out sram[2425]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[42], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2418] sram->in sram[2418]->out sram[2418]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2418]->out) 0
.nodeset V(sram[2418]->outb) vsp
Xsram[2419] sram->in sram[2419]->out sram[2419]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2419]->out) 0
.nodeset V(sram[2419]->outb) vsp
Xsram[2420] sram->in sram[2420]->out sram[2420]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2420]->out) 0
.nodeset V(sram[2420]->outb) vsp
Xsram[2421] sram->in sram[2421]->out sram[2421]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2421]->out) 0
.nodeset V(sram[2421]->outb) vsp
Xsram[2422] sram->in sram[2422]->out sram[2422]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2422]->out) 0
.nodeset V(sram[2422]->outb) vsp
Xsram[2423] sram->in sram[2423]->out sram[2423]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2423]->out) 0
.nodeset V(sram[2423]->outb) vsp
Xsram[2424] sram->in sram[2424]->out sram[2424]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2424]->out) 0
.nodeset V(sram[2424]->outb) vsp
Xsram[2425] sram->in sram[2425]->out sram[2425]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2425]->out) 0
.nodeset V(sram[2425]->outb) vsp
Xmux_2level_tapbuf_size16[43] chany[0][1]_midout[8] chany[0][1]_midout[9] chany[0][1]_midout[22] chany[0][1]_midout[23] chany[0][1]_midout[34] chany[0][1]_midout[35] chany[0][1]_midout[46] chany[0][1]_midout[47] chany[0][1]_midout[58] chany[0][1]_midout[59] chany[0][1]_midout[72] chany[0][1]_midout[73] chany[0][1]_midout[84] chany[0][1]_midout[85] chany[0][1]_midout[96] chany[0][1]_midout[97] grid[1][1]_pin[0][3][31] sram[2426]->outb sram[2426]->out sram[2427]->out sram[2427]->outb sram[2428]->out sram[2428]->outb sram[2429]->out sram[2429]->outb sram[2430]->outb sram[2430]->out sram[2431]->out sram[2431]->outb sram[2432]->out sram[2432]->outb sram[2433]->out sram[2433]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[43], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2426] sram->in sram[2426]->out sram[2426]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2426]->out) 0
.nodeset V(sram[2426]->outb) vsp
Xsram[2427] sram->in sram[2427]->out sram[2427]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2427]->out) 0
.nodeset V(sram[2427]->outb) vsp
Xsram[2428] sram->in sram[2428]->out sram[2428]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2428]->out) 0
.nodeset V(sram[2428]->outb) vsp
Xsram[2429] sram->in sram[2429]->out sram[2429]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2429]->out) 0
.nodeset V(sram[2429]->outb) vsp
Xsram[2430] sram->in sram[2430]->out sram[2430]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2430]->out) 0
.nodeset V(sram[2430]->outb) vsp
Xsram[2431] sram->in sram[2431]->out sram[2431]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2431]->out) 0
.nodeset V(sram[2431]->outb) vsp
Xsram[2432] sram->in sram[2432]->out sram[2432]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2432]->out) 0
.nodeset V(sram[2432]->outb) vsp
Xsram[2433] sram->in sram[2433]->out sram[2433]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2433]->out) 0
.nodeset V(sram[2433]->outb) vsp
Xmux_2level_tapbuf_size16[44] chany[0][1]_midout[10] chany[0][1]_midout[11] chany[0][1]_midout[22] chany[0][1]_midout[23] chany[0][1]_midout[34] chany[0][1]_midout[35] chany[0][1]_midout[48] chany[0][1]_midout[49] chany[0][1]_midout[60] chany[0][1]_midout[61] chany[0][1]_midout[72] chany[0][1]_midout[73] chany[0][1]_midout[84] chany[0][1]_midout[85] chany[0][1]_midout[98] chany[0][1]_midout[99] grid[1][1]_pin[0][3][35] sram[2434]->outb sram[2434]->out sram[2435]->out sram[2435]->outb sram[2436]->out sram[2436]->outb sram[2437]->out sram[2437]->outb sram[2438]->outb sram[2438]->out sram[2439]->out sram[2439]->outb sram[2440]->out sram[2440]->outb sram[2441]->out sram[2441]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[44], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2434] sram->in sram[2434]->out sram[2434]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2434]->out) 0
.nodeset V(sram[2434]->outb) vsp
Xsram[2435] sram->in sram[2435]->out sram[2435]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2435]->out) 0
.nodeset V(sram[2435]->outb) vsp
Xsram[2436] sram->in sram[2436]->out sram[2436]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2436]->out) 0
.nodeset V(sram[2436]->outb) vsp
Xsram[2437] sram->in sram[2437]->out sram[2437]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2437]->out) 0
.nodeset V(sram[2437]->outb) vsp
Xsram[2438] sram->in sram[2438]->out sram[2438]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2438]->out) 0
.nodeset V(sram[2438]->outb) vsp
Xsram[2439] sram->in sram[2439]->out sram[2439]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2439]->out) 0
.nodeset V(sram[2439]->outb) vsp
Xsram[2440] sram->in sram[2440]->out sram[2440]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2440]->out) 0
.nodeset V(sram[2440]->outb) vsp
Xsram[2441] sram->in sram[2441]->out sram[2441]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2441]->out) 0
.nodeset V(sram[2441]->outb) vsp
Xmux_2level_tapbuf_size16[45] chany[0][1]_midout[12] chany[0][1]_midout[13] chany[0][1]_midout[24] chany[0][1]_midout[25] chany[0][1]_midout[36] chany[0][1]_midout[37] chany[0][1]_midout[48] chany[0][1]_midout[49] chany[0][1]_midout[62] chany[0][1]_midout[63] chany[0][1]_midout[74] chany[0][1]_midout[75] chany[0][1]_midout[86] chany[0][1]_midout[87] chany[0][1]_midout[98] chany[0][1]_midout[99] grid[1][1]_pin[0][3][39] sram[2442]->outb sram[2442]->out sram[2443]->out sram[2443]->outb sram[2444]->out sram[2444]->outb sram[2445]->out sram[2445]->outb sram[2446]->outb sram[2446]->out sram[2447]->out sram[2447]->outb sram[2448]->out sram[2448]->outb sram[2449]->out sram[2449]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[45], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2442] sram->in sram[2442]->out sram[2442]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2442]->out) 0
.nodeset V(sram[2442]->outb) vsp
Xsram[2443] sram->in sram[2443]->out sram[2443]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2443]->out) 0
.nodeset V(sram[2443]->outb) vsp
Xsram[2444] sram->in sram[2444]->out sram[2444]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2444]->out) 0
.nodeset V(sram[2444]->outb) vsp
Xsram[2445] sram->in sram[2445]->out sram[2445]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2445]->out) 0
.nodeset V(sram[2445]->outb) vsp
Xsram[2446] sram->in sram[2446]->out sram[2446]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2446]->out) 0
.nodeset V(sram[2446]->outb) vsp
Xsram[2447] sram->in sram[2447]->out sram[2447]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2447]->out) 0
.nodeset V(sram[2447]->outb) vsp
Xsram[2448] sram->in sram[2448]->out sram[2448]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2448]->out) 0
.nodeset V(sram[2448]->outb) vsp
Xsram[2449] sram->in sram[2449]->out sram[2449]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2449]->out) 0
.nodeset V(sram[2449]->outb) vsp
Xmux_2level_tapbuf_size16[46] chany[0][1]_midout[0] chany[0][1]_midout[1] chany[0][1]_midout[12] chany[0][1]_midout[13] chany[0][1]_midout[24] chany[0][1]_midout[25] chany[0][1]_midout[36] chany[0][1]_midout[37] chany[0][1]_midout[50] chany[0][1]_midout[51] chany[0][1]_midout[62] chany[0][1]_midout[63] chany[0][1]_midout[74] chany[0][1]_midout[75] chany[0][1]_midout[86] chany[0][1]_midout[87] grid[0][1]_pin[0][1][0] sram[2450]->outb sram[2450]->out sram[2451]->out sram[2451]->outb sram[2452]->out sram[2452]->outb sram[2453]->out sram[2453]->outb sram[2454]->outb sram[2454]->out sram[2455]->out sram[2455]->outb sram[2456]->out sram[2456]->outb sram[2457]->out sram[2457]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[46], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2450] sram->in sram[2450]->out sram[2450]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2450]->out) 0
.nodeset V(sram[2450]->outb) vsp
Xsram[2451] sram->in sram[2451]->out sram[2451]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2451]->out) 0
.nodeset V(sram[2451]->outb) vsp
Xsram[2452] sram->in sram[2452]->out sram[2452]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2452]->out) 0
.nodeset V(sram[2452]->outb) vsp
Xsram[2453] sram->in sram[2453]->out sram[2453]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2453]->out) 0
.nodeset V(sram[2453]->outb) vsp
Xsram[2454] sram->in sram[2454]->out sram[2454]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2454]->out) 0
.nodeset V(sram[2454]->outb) vsp
Xsram[2455] sram->in sram[2455]->out sram[2455]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2455]->out) 0
.nodeset V(sram[2455]->outb) vsp
Xsram[2456] sram->in sram[2456]->out sram[2456]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2456]->out) 0
.nodeset V(sram[2456]->outb) vsp
Xsram[2457] sram->in sram[2457]->out sram[2457]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2457]->out) 0
.nodeset V(sram[2457]->outb) vsp
Xmux_2level_tapbuf_size16[47] chany[0][1]_midout[0] chany[0][1]_midout[1] chany[0][1]_midout[14] chany[0][1]_midout[15] chany[0][1]_midout[26] chany[0][1]_midout[27] chany[0][1]_midout[38] chany[0][1]_midout[39] chany[0][1]_midout[50] chany[0][1]_midout[51] chany[0][1]_midout[64] chany[0][1]_midout[65] chany[0][1]_midout[76] chany[0][1]_midout[77] chany[0][1]_midout[88] chany[0][1]_midout[89] grid[0][1]_pin[0][1][2] sram[2458]->outb sram[2458]->out sram[2459]->out sram[2459]->outb sram[2460]->out sram[2460]->outb sram[2461]->out sram[2461]->outb sram[2462]->outb sram[2462]->out sram[2463]->out sram[2463]->outb sram[2464]->out sram[2464]->outb sram[2465]->out sram[2465]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[47], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2458] sram->in sram[2458]->out sram[2458]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2458]->out) 0
.nodeset V(sram[2458]->outb) vsp
Xsram[2459] sram->in sram[2459]->out sram[2459]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2459]->out) 0
.nodeset V(sram[2459]->outb) vsp
Xsram[2460] sram->in sram[2460]->out sram[2460]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2460]->out) 0
.nodeset V(sram[2460]->outb) vsp
Xsram[2461] sram->in sram[2461]->out sram[2461]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2461]->out) 0
.nodeset V(sram[2461]->outb) vsp
Xsram[2462] sram->in sram[2462]->out sram[2462]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2462]->out) 0
.nodeset V(sram[2462]->outb) vsp
Xsram[2463] sram->in sram[2463]->out sram[2463]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2463]->out) 0
.nodeset V(sram[2463]->outb) vsp
Xsram[2464] sram->in sram[2464]->out sram[2464]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2464]->out) 0
.nodeset V(sram[2464]->outb) vsp
Xsram[2465] sram->in sram[2465]->out sram[2465]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2465]->out) 0
.nodeset V(sram[2465]->outb) vsp
Xmux_2level_tapbuf_size16[48] chany[0][1]_midout[2] chany[0][1]_midout[3] chany[0][1]_midout[16] chany[0][1]_midout[17] chany[0][1]_midout[28] chany[0][1]_midout[29] chany[0][1]_midout[40] chany[0][1]_midout[41] chany[0][1]_midout[52] chany[0][1]_midout[53] chany[0][1]_midout[66] chany[0][1]_midout[67] chany[0][1]_midout[78] chany[0][1]_midout[79] chany[0][1]_midout[90] chany[0][1]_midout[91] grid[0][1]_pin[0][1][4] sram[2466]->outb sram[2466]->out sram[2467]->out sram[2467]->outb sram[2468]->out sram[2468]->outb sram[2469]->out sram[2469]->outb sram[2470]->outb sram[2470]->out sram[2471]->out sram[2471]->outb sram[2472]->out sram[2472]->outb sram[2473]->out sram[2473]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[48], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2466] sram->in sram[2466]->out sram[2466]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2466]->out) 0
.nodeset V(sram[2466]->outb) vsp
Xsram[2467] sram->in sram[2467]->out sram[2467]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2467]->out) 0
.nodeset V(sram[2467]->outb) vsp
Xsram[2468] sram->in sram[2468]->out sram[2468]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2468]->out) 0
.nodeset V(sram[2468]->outb) vsp
Xsram[2469] sram->in sram[2469]->out sram[2469]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2469]->out) 0
.nodeset V(sram[2469]->outb) vsp
Xsram[2470] sram->in sram[2470]->out sram[2470]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2470]->out) 0
.nodeset V(sram[2470]->outb) vsp
Xsram[2471] sram->in sram[2471]->out sram[2471]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2471]->out) 0
.nodeset V(sram[2471]->outb) vsp
Xsram[2472] sram->in sram[2472]->out sram[2472]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2472]->out) 0
.nodeset V(sram[2472]->outb) vsp
Xsram[2473] sram->in sram[2473]->out sram[2473]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2473]->out) 0
.nodeset V(sram[2473]->outb) vsp
Xmux_2level_tapbuf_size16[49] chany[0][1]_midout[4] chany[0][1]_midout[5] chany[0][1]_midout[16] chany[0][1]_midout[17] chany[0][1]_midout[30] chany[0][1]_midout[31] chany[0][1]_midout[42] chany[0][1]_midout[43] chany[0][1]_midout[54] chany[0][1]_midout[55] chany[0][1]_midout[66] chany[0][1]_midout[67] chany[0][1]_midout[80] chany[0][1]_midout[81] chany[0][1]_midout[92] chany[0][1]_midout[93] grid[0][1]_pin[0][1][6] sram[2474]->outb sram[2474]->out sram[2475]->out sram[2475]->outb sram[2476]->out sram[2476]->outb sram[2477]->out sram[2477]->outb sram[2478]->outb sram[2478]->out sram[2479]->out sram[2479]->outb sram[2480]->out sram[2480]->outb sram[2481]->out sram[2481]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[49], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2474] sram->in sram[2474]->out sram[2474]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2474]->out) 0
.nodeset V(sram[2474]->outb) vsp
Xsram[2475] sram->in sram[2475]->out sram[2475]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2475]->out) 0
.nodeset V(sram[2475]->outb) vsp
Xsram[2476] sram->in sram[2476]->out sram[2476]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2476]->out) 0
.nodeset V(sram[2476]->outb) vsp
Xsram[2477] sram->in sram[2477]->out sram[2477]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2477]->out) 0
.nodeset V(sram[2477]->outb) vsp
Xsram[2478] sram->in sram[2478]->out sram[2478]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2478]->out) 0
.nodeset V(sram[2478]->outb) vsp
Xsram[2479] sram->in sram[2479]->out sram[2479]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2479]->out) 0
.nodeset V(sram[2479]->outb) vsp
Xsram[2480] sram->in sram[2480]->out sram[2480]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2480]->out) 0
.nodeset V(sram[2480]->outb) vsp
Xsram[2481] sram->in sram[2481]->out sram[2481]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2481]->out) 0
.nodeset V(sram[2481]->outb) vsp
Xmux_2level_tapbuf_size16[50] chany[0][1]_midout[6] chany[0][1]_midout[7] chany[0][1]_midout[18] chany[0][1]_midout[19] chany[0][1]_midout[30] chany[0][1]_midout[31] chany[0][1]_midout[44] chany[0][1]_midout[45] chany[0][1]_midout[56] chany[0][1]_midout[57] chany[0][1]_midout[68] chany[0][1]_midout[69] chany[0][1]_midout[80] chany[0][1]_midout[81] chany[0][1]_midout[94] chany[0][1]_midout[95] grid[0][1]_pin[0][1][8] sram[2482]->outb sram[2482]->out sram[2483]->out sram[2483]->outb sram[2484]->out sram[2484]->outb sram[2485]->out sram[2485]->outb sram[2486]->outb sram[2486]->out sram[2487]->out sram[2487]->outb sram[2488]->out sram[2488]->outb sram[2489]->out sram[2489]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[50], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2482] sram->in sram[2482]->out sram[2482]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2482]->out) 0
.nodeset V(sram[2482]->outb) vsp
Xsram[2483] sram->in sram[2483]->out sram[2483]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2483]->out) 0
.nodeset V(sram[2483]->outb) vsp
Xsram[2484] sram->in sram[2484]->out sram[2484]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2484]->out) 0
.nodeset V(sram[2484]->outb) vsp
Xsram[2485] sram->in sram[2485]->out sram[2485]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2485]->out) 0
.nodeset V(sram[2485]->outb) vsp
Xsram[2486] sram->in sram[2486]->out sram[2486]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2486]->out) 0
.nodeset V(sram[2486]->outb) vsp
Xsram[2487] sram->in sram[2487]->out sram[2487]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2487]->out) 0
.nodeset V(sram[2487]->outb) vsp
Xsram[2488] sram->in sram[2488]->out sram[2488]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2488]->out) 0
.nodeset V(sram[2488]->outb) vsp
Xsram[2489] sram->in sram[2489]->out sram[2489]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2489]->out) 0
.nodeset V(sram[2489]->outb) vsp
Xmux_2level_tapbuf_size16[51] chany[0][1]_midout[8] chany[0][1]_midout[9] chany[0][1]_midout[20] chany[0][1]_midout[21] chany[0][1]_midout[32] chany[0][1]_midout[33] chany[0][1]_midout[44] chany[0][1]_midout[45] chany[0][1]_midout[58] chany[0][1]_midout[59] chany[0][1]_midout[70] chany[0][1]_midout[71] chany[0][1]_midout[82] chany[0][1]_midout[83] chany[0][1]_midout[94] chany[0][1]_midout[95] grid[0][1]_pin[0][1][10] sram[2490]->outb sram[2490]->out sram[2491]->out sram[2491]->outb sram[2492]->out sram[2492]->outb sram[2493]->out sram[2493]->outb sram[2494]->outb sram[2494]->out sram[2495]->out sram[2495]->outb sram[2496]->out sram[2496]->outb sram[2497]->out sram[2497]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[51], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2490] sram->in sram[2490]->out sram[2490]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2490]->out) 0
.nodeset V(sram[2490]->outb) vsp
Xsram[2491] sram->in sram[2491]->out sram[2491]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2491]->out) 0
.nodeset V(sram[2491]->outb) vsp
Xsram[2492] sram->in sram[2492]->out sram[2492]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2492]->out) 0
.nodeset V(sram[2492]->outb) vsp
Xsram[2493] sram->in sram[2493]->out sram[2493]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2493]->out) 0
.nodeset V(sram[2493]->outb) vsp
Xsram[2494] sram->in sram[2494]->out sram[2494]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2494]->out) 0
.nodeset V(sram[2494]->outb) vsp
Xsram[2495] sram->in sram[2495]->out sram[2495]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2495]->out) 0
.nodeset V(sram[2495]->outb) vsp
Xsram[2496] sram->in sram[2496]->out sram[2496]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2496]->out) 0
.nodeset V(sram[2496]->outb) vsp
Xsram[2497] sram->in sram[2497]->out sram[2497]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2497]->out) 0
.nodeset V(sram[2497]->outb) vsp
Xmux_2level_tapbuf_size16[52] chany[0][1]_midout[8] chany[0][1]_midout[9] chany[0][1]_midout[22] chany[0][1]_midout[23] chany[0][1]_midout[34] chany[0][1]_midout[35] chany[0][1]_midout[46] chany[0][1]_midout[47] chany[0][1]_midout[58] chany[0][1]_midout[59] chany[0][1]_midout[72] chany[0][1]_midout[73] chany[0][1]_midout[84] chany[0][1]_midout[85] chany[0][1]_midout[96] chany[0][1]_midout[97] grid[0][1]_pin[0][1][12] sram[2498]->outb sram[2498]->out sram[2499]->out sram[2499]->outb sram[2500]->out sram[2500]->outb sram[2501]->out sram[2501]->outb sram[2502]->outb sram[2502]->out sram[2503]->out sram[2503]->outb sram[2504]->out sram[2504]->outb sram[2505]->out sram[2505]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[52], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2498] sram->in sram[2498]->out sram[2498]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2498]->out) 0
.nodeset V(sram[2498]->outb) vsp
Xsram[2499] sram->in sram[2499]->out sram[2499]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2499]->out) 0
.nodeset V(sram[2499]->outb) vsp
Xsram[2500] sram->in sram[2500]->out sram[2500]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2500]->out) 0
.nodeset V(sram[2500]->outb) vsp
Xsram[2501] sram->in sram[2501]->out sram[2501]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2501]->out) 0
.nodeset V(sram[2501]->outb) vsp
Xsram[2502] sram->in sram[2502]->out sram[2502]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2502]->out) 0
.nodeset V(sram[2502]->outb) vsp
Xsram[2503] sram->in sram[2503]->out sram[2503]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2503]->out) 0
.nodeset V(sram[2503]->outb) vsp
Xsram[2504] sram->in sram[2504]->out sram[2504]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2504]->out) 0
.nodeset V(sram[2504]->outb) vsp
Xsram[2505] sram->in sram[2505]->out sram[2505]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2505]->out) 0
.nodeset V(sram[2505]->outb) vsp
Xmux_2level_tapbuf_size16[53] chany[0][1]_midout[10] chany[0][1]_midout[11] chany[0][1]_midout[22] chany[0][1]_midout[23] chany[0][1]_midout[36] chany[0][1]_midout[37] chany[0][1]_midout[48] chany[0][1]_midout[49] chany[0][1]_midout[60] chany[0][1]_midout[61] chany[0][1]_midout[72] chany[0][1]_midout[73] chany[0][1]_midout[86] chany[0][1]_midout[87] chany[0][1]_midout[98] chany[0][1]_midout[99] grid[0][1]_pin[0][1][14] sram[2506]->outb sram[2506]->out sram[2507]->out sram[2507]->outb sram[2508]->out sram[2508]->outb sram[2509]->out sram[2509]->outb sram[2510]->outb sram[2510]->out sram[2511]->out sram[2511]->outb sram[2512]->out sram[2512]->outb sram[2513]->out sram[2513]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[53], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2506] sram->in sram[2506]->out sram[2506]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2506]->out) 0
.nodeset V(sram[2506]->outb) vsp
Xsram[2507] sram->in sram[2507]->out sram[2507]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2507]->out) 0
.nodeset V(sram[2507]->outb) vsp
Xsram[2508] sram->in sram[2508]->out sram[2508]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2508]->out) 0
.nodeset V(sram[2508]->outb) vsp
Xsram[2509] sram->in sram[2509]->out sram[2509]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2509]->out) 0
.nodeset V(sram[2509]->outb) vsp
Xsram[2510] sram->in sram[2510]->out sram[2510]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2510]->out) 0
.nodeset V(sram[2510]->outb) vsp
Xsram[2511] sram->in sram[2511]->out sram[2511]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2511]->out) 0
.nodeset V(sram[2511]->outb) vsp
Xsram[2512] sram->in sram[2512]->out sram[2512]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2512]->out) 0
.nodeset V(sram[2512]->outb) vsp
Xsram[2513] sram->in sram[2513]->out sram[2513]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2513]->out) 0
.nodeset V(sram[2513]->outb) vsp
.eom
