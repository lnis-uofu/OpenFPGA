// Benchmark "TOP" written by ABC on Mon Feb  4 17:33:19 2019

module pdc ( 
    i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_,
    i_11_, i_12_, i_13_, i_14_, i_15_,
    o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_,
    o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_,
    o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_,
    o_31_, o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_  );
  input  i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_,
    i_10_, i_11_, i_12_, i_13_, i_14_, i_15_;
  output o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_,
    o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_,
    o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_,
    o_31_, o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_;
  wire n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
    n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
    n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
    n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
    n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
    n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
    n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
    n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
    n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
    n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
    n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
    n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
    n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
    n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
    n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
    n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
    n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
    n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
    n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
    n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
    n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
    n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
    n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
    n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
    n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
    n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
    n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
    n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
    n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
    n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
    n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
    n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
    n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
    n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
    n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
    n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
    n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
    n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
    n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
    n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
    n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
    n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
    n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
    n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
    n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
    n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
    n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
    n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
    n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
    n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
    n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
    n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
    n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
    n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
    n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
    n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
    n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
    n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
    n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
    n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
    n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
    n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
    n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
    n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
    n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
    n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
    n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
    n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
    n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
    n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
    n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
    n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
    n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
    n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
    n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
    n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
    n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
    n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
    n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
    n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
    n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
    n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
    n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
    n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
    n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
    n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
    n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
    n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
    n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
    n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
    n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
    n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
    n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
    n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
    n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
    n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
    n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
    n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
    n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
    n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
    n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
    n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
    n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
    n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
    n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
    n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
    n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
    n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
    n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
    n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
    n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
    n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
    n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
    n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
    n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
    n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
    n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
    n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
    n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
    n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
    n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
    n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
    n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
    n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
    n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
    n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
    n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
    n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
    n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
    n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
    n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
    n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
    n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
    n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
    n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
    n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
    n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
    n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
    n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
    n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
    n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
    n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
    n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
    n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
    n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
    n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
    n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
    n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
    n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
    n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
    n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
    n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
    n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
    n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
    n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
    n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
    n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
    n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
    n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
    n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
    n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
    n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
    n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
    n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
    n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
    n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
    n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
    n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
    n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
    n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
    n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
    n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
    n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
    n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
    n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
    n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
    n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
    n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
    n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
    n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
    n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
    n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
    n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
    n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
    n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
    n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
    n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
    n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
    n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
    n2376, n2377, n2378, n2379, n2380, n2381;
  assign o_0_ = ~n126 & (n124 | n161);
  assign o_1_ = ~n126 & (n160 | ~n1042 | ~n1612);
  assign o_2_ = ~n126 & (n158 | n159 | ~n714);
  assign o_3_ = ~n126 & (~n2261 | ~n2266);
  assign o_4_ = ~n126 & (~n2241 | ~n2250 | ~n2252);
  assign o_5_ = ~n2380;
  assign o_6_ = ~n157;
  assign o_7_ = ~n126 & (n156 | ~n1365 | ~n1370);
  assign o_8_ = ~n2379;
  assign o_9_ = ~n126 & (n155 | ~n1984 | ~n1986);
  assign o_10_ = ~n154;
  assign o_11_ = ~n995;
  assign o_12_ = ~n1187;
  assign o_13_ = ~n1174;
  assign o_14_ = ~n1353;
  assign o_15_ = ~n152;
  assign o_16_ = ~n126 & (~n2359 | ~n2361 | ~n2363);
  assign o_17_ = ~n126 & (~n2347 | ~n2349 | ~n2351);
  assign o_18_ = ~n126 & (~n2332 | ~n2334 | ~n2336);
  assign o_19_ = ~n126 & (~n2318 | ~n2319 | ~n2320);
  assign o_20_ = ~n126 & (~n2302 | ~n2304);
  assign o_21_ = ~n151;
  assign o_22_ = ~n927 | ~n1431 | n148 | n149;
  assign o_23_ = ~n147;
  assign o_24_ = ~n145;
  assign o_25_ = ~n144;
  assign o_26_ = ~n142;
  assign o_27_ = n136 & ~n126 & n135;
  assign o_28_ = ~n2378;
  assign o_29_ = ~n126 & (~n866 | ~n2284 | ~n2285);
  assign o_30_ = ~n134;
  assign o_31_ = n132 | n130 | n131;
  assign o_32_ = ~n129;
  assign o_33_ = ~n2377;
  assign o_34_ = ~n126 & (~n2280 | ~n2282);
  assign o_35_ = ~n126 & (~n1622 | ~n1625 | ~n2278);
  assign o_36_ = ~n128;
  assign o_37_ = ~n126 & (n123 | n124 | n125);
  assign o_38_ = n121 & ~n1251;
  assign o_39_ = n121 & n122;
  assign n96 = n1239 & n1264;
  assign n97 = n1239 & n177;
  assign n98 = n1228 & n1239;
  assign n99 = ~n361 | ~n1373;
  assign n100 = n98 & (n99 | ~n617);
  assign n101 = n96 & (~n564 | ~n926);
  assign n102 = ~n617 | ~n1176;
  assign n103 = n96 & (n102 | ~n361);
  assign n104 = n1252 & n1256;
  assign n105 = ~n597 | ~n1377;
  assign n106 = n104 & (n105 | ~n500);
  assign n107 = n1256 & n1264;
  assign n108 = n107 & (~n336 | ~n1334);
  assign n109 = ~n305 | ~n653;
  assign n110 = n107 & (n109 | ~n685);
  assign n111 = n107 & (~n426 | ~n1378);
  assign n112 = n107 & (~n777 | ~n1795);
  assign n113 = ~n1214 & n1256;
  assign n114 = n113 & (~n1330 | ~n1418);
  assign n115 = n113 & (~n774 | ~n1795);
  assign n116 = n1228 & n1231;
  assign n117 = n116 & (~n653 | ~n1378);
  assign n118 = n113 & (~n266 | ~n1175);
  assign n119 = ~n226 | ~n845;
  assign n120 = n116 & (n119 | ~n472);
  assign n121 = n172 & (n173 | n174);
  assign n122 = i_6_ & ~i_7_;
  assign n123 = n178 & n1228;
  assign n124 = ~n1365 | ~n1370 | n159 | ~n714;
  assign n125 = n2267 | n1647 | n717;
  assign n126 = ~n1988 | ~n1989 | n184 | n185 | ~n157 | n175 | n180 | n182;
  assign n127 = ~n2277 & n1618 & n1617 & n923 & n748 & n817;
  assign n128 = n126 | n127;
  assign n129 = n895 & n896 & (~n136 | ~n1237);
  assign n130 = ~n481 & (n897 | n898);
  assign n131 = n899 & (n900 | n901);
  assign n132 = n1646 | n1647;
  assign n133 = n1990 & n1648 & n1365 & n904 & n895 & n863 & ~n159 & n460;
  assign n134 = n126 | n133;
  assign n135 = ~i_2_ & i_0_ & i_1_;
  assign n136 = i_6_ & i_7_;
  assign n137 = n907 | n777;
  assign n138 = n916 & n917 & (n918 | n911);
  assign n139 = n1654 & n1653 & n1652 & n1651 & ~n915 & n1650;
  assign n140 = n1658 & n1657 & n1656 & n1655 & ~n913 & n914;
  assign n141 = n1661 & n1660 & n1659 & n912 & ~n171 & n909;
  assign n142 = n141 & n140 & n139 & n137 & n138;
  assign n143 = n2288 & n919 & n1617 & n815 & n740 & n1457 & n747 & n746;
  assign n144 = n126 | n143;
  assign n145 = n923 & (~n161 | n924);
  assign n146 = n748 & n817 & n727 & n889 & n1622 & n862;
  assign n147 = n126 | n146;
  assign n148 = n929 & (~n984 | ~n1141);
  assign n149 = n928 & (~n677 | ~n1663);
  assign n150 = n978 & n977 & n976 & n938 & n975 & n974 & n972 & n973;
  assign n151 = n126 | n150;
  assign n152 = n187 & (~i_0_ | i_1_ | i_2_);
  assign n153 = n1859 & n927 & n1644 & n769 & n1537 & n1617 & n1618;
  assign n154 = n126 | n153;
  assign n155 = ~n1973 | ~n1977 | ~n358 | n1972 | n347 | n350 | n352 | n355;
  assign n156 = n1213 & ~n1214;
  assign n157 = (~i_3_ | n186) & (n187 | n188);
  assign n158 = n1213 & n176;
  assign n159 = n1215 & ~n1353;
  assign n160 = ~n481 & ~n1235;
  assign n161 = n158 | n156;
  assign n162 = n98 & (~n362 | ~n495);
  assign n163 = n1239 & n1252;
  assign n164 = n163 & (~n216 | ~n316);
  assign n165 = ~n1233 & n1253;
  assign n166 = n165 & (~n654 | ~n1012);
  assign n167 = n176 & n1231;
  assign n168 = n167 & (~n1176 | ~n1373);
  assign n169 = n107 & (~n329 | ~n1416);
  assign n170 = n167 & (~n709 | ~n1335);
  assign n171 = ~n907 & (~n879 | ~n979);
  assign n172 = ~i_2_ & ~i_0_ & i_1_;
  assign n173 = i_3_ & i_5_ & i_4_;
  assign n174 = ~i_5_ & i_3_ & i_4_;
  assign n175 = ~n2381 & (n156 | n158);
  assign n176 = n122 & i_8_;
  assign n177 = i_8_ & n136;
  assign n178 = n172 & n1215;
  assign n179 = n172 & n1216;
  assign n180 = (n176 | n177) & (n178 | n179);
  assign n181 = n1228 & n179;
  assign n182 = (~n1227 | ~n1987) & (n123 | n181);
  assign n183 = n1216 | ~n1229 | i_3_ | ~n1212;
  assign n184 = n135 & n183;
  assign n185 = ~n1235 & (~n1227 | (i_12_ & ~n943));
  assign n186 = i_0_ | i_1_ | i_2_;
  assign n187 = i_0_ | ~i_2_;
  assign n188 = i_1_ | ~i_3_;
  assign n189 = ~n98 | n316;
  assign n190 = n1240 | n1245;
  assign n191 = n1240 | n1243;
  assign n192 = n189 & (~n98 | (n190 & n191));
  assign n193 = ~n98 | n317;
  assign n194 = ~n98 | n287;
  assign n195 = n1245 | n1260;
  assign n196 = n193 & n194 & (~n98 | n195);
  assign n197 = ~n98 | n979;
  assign n198 = n264 & n1207;
  assign n199 = n197 & (~n98 | n198);
  assign n200 = ~n98 | n1105;
  assign n201 = n329 & n444;
  assign n202 = n200 & (~n98 | n201);
  assign n203 = ~n98 | n1262;
  assign n204 = n1238 | n1245;
  assign n205 = n203 & (~n98 | n204);
  assign n206 = n1198 | n1263;
  assign n207 = n205 & (~n98 | n206);
  assign n208 = ~n98 | n527;
  assign n209 = n330 & n442;
  assign n210 = n208 & (~n98 | n209);
  assign n211 = ~n97 | n284;
  assign n212 = n313 & n226;
  assign n213 = n211 & (~n97 | n212);
  assign n214 = ~n97 | n191;
  assign n215 = n214 & (~n97 | n190);
  assign n216 = n1198 | n1206;
  assign n217 = n215 & (~n97 | n216);
  assign n218 = ~n97 | n287;
  assign n219 = n195 & n356;
  assign n220 = n218 & (~n97 | n219);
  assign n221 = ~n97 | n1105;
  assign n222 = n221 & (~n97 | n201);
  assign n223 = ~n97 | n527;
  assign n224 = n223 & (~n97 | n209);
  assign n225 = ~n167 | n444;
  assign n226 = n1198 | n1201;
  assign n227 = n1217 | n1220;
  assign n228 = n225 & (~n167 | (n226 & n227));
  assign n229 = n113 & (~n331 | ~n334);
  assign n230 = n107 & (~n474 | ~n1207);
  assign n231 = ~n96 | n216;
  assign n232 = ~n96 | n251;
  assign n233 = ~n96 | n316;
  assign n234 = ~n96 | n1157;
  assign n235 = ~n96 | n1248;
  assign n236 = n834 & n1475 & n1928 & n1546 & n860 & n827;
  assign n237 = n1930 & n1932 & n1681 & n933 & n934 & n1715 & n955 & n1931;
  assign n238 = n1941 & n1943 & n1944 & n1948 & n1947 & n1838 & n1945 & n1946;
  assign n239 = n238 & n237 & n236 & n235 & n234 & n233 & n231 & n232;
  assign n240 = ~n96 | n1247;
  assign n241 = ~n96 | n204;
  assign n242 = ~n96 | n195;
  assign n243 = ~n278 | n617;
  assign n244 = ~n96 | n264;
  assign n245 = n1927 & (~n278 | (n204 & n306));
  assign n246 = ~n268 | n2036;
  assign n247 = (~n107 | n195) & (n263 | n907);
  assign n248 = n247 & n246 & n245 & n244 & n243 & n242 & n240 & n241;
  assign n249 = ~n167 | n316;
  assign n250 = ~n96 | n317;
  assign n251 = n1220 | n1238;
  assign n252 = n249 & n250 & (~n107 | n251);
  assign n253 = n278 | n107;
  assign n254 = ~n755 & (n97 | n253);
  assign n255 = ~n96 | n331;
  assign n256 = ~n113 | n1250;
  assign n257 = (~n107 | n1295) & (~n633 | n1866);
  assign n258 = (~n96 | n190) & (~n97 | n749);
  assign n259 = (~n167 | ~n268) & (n924 | n1968);
  assign n260 = n252 & n248 & n239 & n1282 & n1286 & n1054 & n217 & n220;
  assign n261 = n1962 & n1964 & n1967 & n1966 & n1965 & n1800 & n1842 & n1818;
  assign n262 = n261 & n260 & n259 & n258 & n257 & n256 & ~n254 & n255;
  assign n263 = n195 & n305;
  assign n264 = n1219 | n1245;
  assign n265 = ~i_15_ | n1218;
  assign n266 = n1197 | n1204;
  assign n267 = n266 & n265 & n263 & n264;
  assign n268 = ~n190 | ~n617;
  assign n269 = ~n327 & (~n263 | n268);
  assign n270 = ~n167 | n604;
  assign n271 = ~n167 | n204;
  assign n272 = n1923 & (n1924 | n313);
  assign n273 = (~n107 | n597) & (~n167 | n330);
  assign n274 = n1926 & (~n348 | n604);
  assign n275 = n1712 & n1502 & n1706 & n1750 & n1674 & n1680;
  assign n276 = n1594 & n1860 & n1548 & n1602 & n1568 & n1573;
  assign n277 = n276 & n275 & n274 & n273 & n272 & n271 & ~n269 & n270;
  assign n278 = ~n1214 & n1253;
  assign n279 = n278 & (~n284 | ~n287);
  assign n280 = n191 | ~n353;
  assign n281 = n116 & (~n287 | ~n979);
  assign n282 = n1105 & n309;
  assign n283 = ~n104 | n282;
  assign n284 = n1217 | n1243;
  assign n285 = ~n104 & ~n116;
  assign n286 = n284 | n285;
  assign n287 = n1243 | n1260;
  assign n288 = n1204 | n1238;
  assign n289 = n191 & n536 & n926;
  assign n290 = n289 & n287 & n288;
  assign n291 = ~n571 & n1292;
  assign n292 = ~n381 & n1291;
  assign n293 = n292 & n291 & ~n113 & ~n163;
  assign n294 = n113 | n571;
  assign n295 = n165 | n107;
  assign n296 = ~n674 & (n167 | n294 | n295);
  assign n297 = n1300 & n1299 & n1298 & n1297 & n1296 & n286 & ~n281 & n283;
  assign n298 = n563 & n561 & n497;
  assign n299 = (~n107 | n508) & (~n278 | n288);
  assign n300 = (n292 | n879) & (~n96 | n926);
  assign n301 = (n290 | ~n404) & (~n253 | n1293);
  assign n302 = n1910 & n1909 & n1400 & n1398 & n1396 & n559 & ~n296 & n483;
  assign n303 = n302 & n301 & n300 & n299 & n297 & n298;
  assign n304 = n610 & n604;
  assign n305 = n1204 | n1265;
  assign n306 = n1204 | n1263;
  assign n307 = n266 & n306 & n304 & n305;
  assign n308 = n1207 & n226;
  assign n309 = n1241 | n1243;
  assign n310 = n206 & n284 & n308 & n309;
  assign n311 = ~n98 | n227;
  assign n312 = ~n98 | n284;
  assign n313 = n1217 | n1245;
  assign n314 = n311 & n312 & (~n98 | n313);
  assign n315 = n314 & (~n98 | n226);
  assign n316 = n1220 | n1240;
  assign n317 = n1220 | n1260;
  assign n318 = n317 & n316 & n216;
  assign n319 = n316 & n474;
  assign n320 = ~n165 | n319;
  assign n321 = n571 | n104;
  assign n322 = n321 & (~n227 | ~n822 | ~n1157);
  assign n323 = ~n165 & ~n571;
  assign n324 = n317 | n323;
  assign n325 = n1308 & n1307 & n1306 & n1305 & n1304 & n1303 & n1301 & n1302;
  assign n326 = n487 & n494 & (n318 | ~n404);
  assign n327 = ~n294 & n1290;
  assign n328 = n325 & n326 & (n327 | n251);
  assign n329 = n1245 | n1249;
  assign n330 = n1245 | n1255;
  assign n331 = n1198 | n1255;
  assign n332 = n331 & n329 & n330;
  assign n333 = n1250 & n334;
  assign n334 = n1198 | n1217;
  assign n335 = (n291 | n333) & (~n98 | n334);
  assign n336 = n1247 & n1248;
  assign n337 = n336 & n316 & n204;
  assign n338 = n343 | n354;
  assign n339 = n338 & (~n755 | ~n924);
  assign n340 = n165 | ~n291;
  assign n341 = n340 & (~n921 | ~n1262);
  assign n342 = n294 & (~n287 | ~n474);
  assign n343 = n404 | n163;
  assign n344 = ~n327 | n348;
  assign n345 = ~n774 & (n343 | n344);
  assign n346 = n404 | n165;
  assign n347 = ~n1250 & (n96 | n346);
  assign n348 = n98 | n97;
  assign n349 = n113 | ~n291;
  assign n350 = ~n265 & (n348 | n349);
  assign n351 = n359 | n381 | n344;
  assign n352 = ~n597 & (n278 | n351);
  assign n353 = n1231 & n177;
  assign n354 = n98 | ~n327;
  assign n355 = ~n216 & (n353 | n354);
  assign n356 = n1198 | n1265;
  assign n357 = ~n98 & n1309;
  assign n358 = n356 | n357;
  assign n359 = n163 | n96;
  assign n360 = n359 & (~n265 | ~n604 | ~n1311);
  assign n361 = n1206 | n1221;
  assign n362 = n1197 | n1245;
  assign n363 = n361 & n362;
  assign n364 = ~n97 | n495;
  assign n365 = ~n97 | n566;
  assign n366 = ~n96 | n447;
  assign n367 = ~n96 | n426;
  assign n368 = ~n96 | n688;
  assign n369 = n1604 & n1701 & n2075 & n2076;
  assign n370 = n2081 & n947 & n1719 & n2080 & n2079 & n998 & n2077 & n2078;
  assign n371 = n2085 & n2086 & n1089 & n1846 & n1016 & n1007 & n1864 & n2087;
  assign n372 = n371 & n370 & n369 & n368 & n367 & n366 & n364 & n365;
  assign n373 = (~n116 | n1138) & (~n404 | n447);
  assign n374 = n2109 & (n361 | ~n381);
  assign n375 = n2108 & (~n165 | (n426 & n1331));
  assign n376 = n1131 & n1132 & n1078 & n2107;
  assign n377 = n2103 & n2106 & n916 & n1810 & n1785 & n1822 & n2104 & n2105;
  assign n378 = n2097 & n1709 & n2101 & n2100 & n2099 & n1697 & n2098 & n1687;
  assign n379 = n2091 & n1484 & n2094 & n1525 & n2093 & n1574 & n2092 & n1565;
  assign n380 = n379 & n378 & n377 & n376 & n375 & n374 & n373 & n372;
  assign n381 = n404 | n167;
  assign n382 = n163 | n107;
  assign n383 = ~n845 & (n381 | n382);
  assign n384 = ~n167 | n1331;
  assign n385 = ~n167 | n688;
  assign n386 = ~n278 | n1331;
  assign n387 = ~n96 | n845;
  assign n388 = n2110 & (~n107 | (n426 & n688));
  assign n389 = (~n163 | n361) & (~n167 | n426);
  assign n390 = n2111 & (~n348 | n1331);
  assign n391 = n390 & n380 & n389 & n388 & n387 & n386 & n384 & n385;
  assign n392 = i_15_ | n1332;
  assign n393 = n1243 | n1257;
  assign n394 = n392 & n393;
  assign n395 = ~n104 | n441;
  assign n396 = ~n104 | n393;
  assign n397 = (n394 | n911) & (~n253 | n1336);
  assign n398 = n1340 & n2071 & (~n116 | n441);
  assign n399 = n2069 & n1000 & n1805 & n1746 & n1747 & n2070;
  assign n400 = n2061 & n2065 & n1776 & n1786 & n1819 & n2066 & n1752 & n1830;
  assign n401 = n2049 & n2051 & n2054 & n2053 & n1694 & n2052 & n1710 & n1685;
  assign n402 = n2043 & n2037 & n770 & n2045 & n2044 & n733 & n1510 & n722;
  assign n403 = n402 & n401 & n400 & n399 & n398 & n397 & n395 & n396;
  assign n404 = n1231 & ~n1232;
  assign n405 = n404 & (~n430 | ~n529 | ~n709);
  assign n406 = ~n167 | n1334;
  assign n407 = ~n278 | n393;
  assign n408 = ~n96 | n441;
  assign n409 = n2073 & (~n278 | n429);
  assign n410 = (~n107 | n1334) & (~n167 | n471);
  assign n411 = n2074 & (~n348 | n393);
  assign n412 = n411 & n410 & n409 & n408 & n407 & n406 & n403 & ~n405;
  assign n413 = ~n107 | n1224;
  assign n414 = ~n113 | n1152;
  assign n415 = ~n113 | n1151;
  assign n416 = ~n107 | n1341;
  assign n417 = n990 & (n2036 | n1145);
  assign n418 = n1345 & n1344 & n1342 & n1343;
  assign n419 = n958 & n2035 & n1439 & n2034 & n2033 & n2032 & n2030 & n2031;
  assign n420 = n2028 & n2029 & n1419 & n1725 & n1471 & n1499 & n1729 & n782;
  assign n421 = n420 & n419 & n418 & n417 & n416 & n415 & n413 & n414;
  assign n422 = ~n96 | n1330;
  assign n423 = n1335 & n1330;
  assign n424 = n421 & n422 & (~n107 | n423);
  assign n425 = ~n97 | n471;
  assign n426 = n1245 | n1265;
  assign n427 = n425 & (~n97 | n426);
  assign n428 = n427 & (~n97 | n356);
  assign n429 = n709 & n473;
  assign n430 = n1221 | n1240;
  assign n431 = n429 & n430;
  assign n432 = ~n107 | n471;
  assign n433 = ~n107 | n1337;
  assign n434 = ~n107 | n472;
  assign n435 = (~n107 | n431) & (n907 | n908);
  assign n436 = ~n278 | n441;
  assign n437 = n2002 & n2001 & n2000 & n1999 & n1998 & n1997 & n989;
  assign n438 = n1993 & n1996 & n1995 & n1714 & n1600 & n1605 & n1994 & n1554;
  assign n439 = n438 & n437 & n436 & n435 & n434 & n433 & ~n170 & n432;
  assign n440 = n1220 | n1246;
  assign n441 = i_15_ | n1225;
  assign n442 = n1198 | n1258;
  assign n443 = n1224 & n1082;
  assign n444 = n1198 | n1257;
  assign n445 = n444 & n443 & n442 & n206 & n441 & n356 & n308 & n440;
  assign n446 = ~n98 | n473;
  assign n447 = n1245 | n1263;
  assign n448 = n446 & (~n98 | n447);
  assign n449 = (n119 | ~n206) & (n97 | n98);
  assign n450 = ~n216 | ~n564;
  assign n451 = ~n327 & (n450 | ~n1347);
  assign n452 = ~n361 & (n96 | n354);
  assign n453 = n163 | ~n292;
  assign n454 = ~n1224 & (n104 | n453);
  assign n455 = ~n291 & (~n316 | ~n685 | ~n1348);
  assign n456 = ~n1145 & (~n327 | n359 | n381);
  assign n457 = ~n1152 & (~n292 | n340 | n359);
  assign n458 = n1230 | n1251;
  assign n459 = n1230 | n1233;
  assign n460 = n458 & (n459 | ~n819);
  assign n461 = n1990 & n1624 & n1620;
  assign n462 = n444 & n508;
  assign n463 = n460 & n461 & (n462 | n459);
  assign n464 = n442 & n469;
  assign n465 = ~n450 & n464;
  assign n466 = (~n97 | n465) & (~n98 | n464);
  assign n467 = n393 & n1331;
  assign n468 = n426 & n845;
  assign n469 = n707 & n656;
  assign n470 = n709 & n362;
  assign n471 = n1243 | n1265;
  assign n472 = n1201 | n1243;
  assign n473 = n1243 | n1263;
  assign n474 = n1219 | n1220;
  assign n475 = n474 & n473 & n472 & n471 & n470 & n469 & n467 & n468;
  assign n476 = ~n362 & (n278 | n381);
  assign n477 = n1363 & n1362 & n1361 & n1360 & n766 & n239 & n439 & n428;
  assign n478 = n2117 & n1359 & n328 & n252;
  assign n479 = n2115 & n2113 & n1041 & n2114 & n2112 & n839 & n1385 & n869;
  assign n480 = n479 & n478 & n477 & n466 & n463 & n391 & n412 & n424;
  assign n481 = i_10_ | i_9_;
  assign n482 = n481 | ~n897;
  assign n483 = ~n98 | n508;
  assign n484 = n483 & (~n98 | n467);
  assign n485 = ~n96 | n227;
  assign n486 = n485 & (~n99 | ~n163);
  assign n487 = ~n163 | n227;
  assign n488 = ~n96 | n1372;
  assign n489 = n1221 | n1246;
  assign n490 = n487 & n488 & (~n96 | n489);
  assign n491 = ~n163 | n1372;
  assign n492 = n250 & n491 & (~n163 | n489);
  assign n493 = ~n96 | n1125;
  assign n494 = ~n163 | n474;
  assign n495 = ~i_15_ | n1223;
  assign n496 = n493 & n494 & (~n96 | n495);
  assign n497 = ~n98 | n1293;
  assign n498 = n497 & (~n98 | n469);
  assign n499 = n1258 | n1371;
  assign n500 = n1221 | n1258;
  assign n501 = n499 & n500;
  assign n502 = (n501 | ~n571) & (~n113 | n251);
  assign n503 = ~n96 | n288;
  assign n504 = n1238 | n1376;
  assign n505 = n422 & n503 & (~n96 | n504);
  assign n506 = n879 | n675;
  assign n507 = ~n107 | n499;
  assign n508 = n1204 | n1249;
  assign n509 = n1233 | ~n1239;
  assign n510 = n506 & n507 & (n508 | n509);
  assign n511 = ~n163 | n1375;
  assign n512 = ~n163 | n530;
  assign n513 = ~n98 | n1374;
  assign n514 = ~n98 | n951;
  assign n515 = n2185 & (~n929 | n984);
  assign n516 = n875 | n509;
  assign n517 = n516 & n515 & n514 & n513 & n511 & n512;
  assign n518 = n682 & n504;
  assign n519 = n1377 & n653;
  assign n520 = n979 & n1262;
  assign n521 = n1240 | n1371;
  assign n522 = n1238 | n1371;
  assign n523 = n1249 | n1376;
  assign n524 = n523 & n522 & n521 & n520 & n518 & n519;
  assign n525 = n430 & n926 & n1176;
  assign n526 = n1217 | n1376;
  assign n527 = n1243 | n1255;
  assign n528 = n1241 | n1376;
  assign n529 = n1221 | n1241;
  assign n530 = n1241 | n1371;
  assign n531 = n530 & n529 & n528 & n527 & n526 & n284 & n282 & n525;
  assign n532 = n107 & (~n1175 | ~n1381 | ~n2184);
  assign n533 = n528 & n1380;
  assign n534 = ~n532 & (~n104 | (n525 & n533));
  assign n535 = ~n278 | n529;
  assign n536 = n1204 | n1241;
  assign n537 = n535 & (~n278 | n536);
  assign n538 = ~n278 | n528;
  assign n539 = ~n453 & n1349;
  assign n540 = n1260 | n1371;
  assign n541 = n538 & n537 & (n539 | n540);
  assign n542 = n107 & (~n523 | ~n530 | ~n1382);
  assign n543 = (~n98 | n592) & (n567 | ~n929);
  assign n544 = (~n96 | n682) & (~n404 | n522);
  assign n545 = n2203 & n2204 & (~n346 | n1375);
  assign n546 = n944 & n765 & n541 & n534 & n517 & n510 & n1387 & n505;
  assign n547 = n2198 & n2199 & n2200 & n2201 & n2197 & n2195 & n2202 & n1283;
  assign n548 = n2191 & n2187 & n2188 & n200 & n2192 & n197 & n221 & n218;
  assign n549 = n548 & n547 & n546 & n545 & n543 & n544;
  assign n550 = n1395 & n1394 & n1393 & n1392 & n1391 & n1090 & n1389 & n1390;
  assign n551 = n1321 & n1320 & n1319 & n1318 & n1317 & n280 & ~n171 & ~n279;
  assign n552 = n2183 & (n1196 | ~n1388);
  assign n553 = (~n113 | n1374) & (n521 | n2036);
  assign n554 = n1843 & n2182 & (~n107 | n520);
  assign n555 = n2178 & n2181 & n1761 & n1061 & n1836 & n2180 & n1095 & n2179;
  assign n556 = n2172 & n1652 & n1659 & n2174 & n959 & n1682 & n2173 & n1728;
  assign n557 = n2171 & n1428 & n1453 & n1479 & n1468 & n1464 & n1534 & n1448;
  assign n558 = n557 & n556 & n555 & n554 & n553 & n552 & n550 & n551;
  assign n559 = ~n97 | n508;
  assign n560 = n559 & (~n97 | n467);
  assign n561 = ~n97 | n1293;
  assign n562 = n561 & (~n97 | n469);
  assign n563 = ~n97 | n926;
  assign n564 = n1337 & n1333;
  assign n565 = n563 & (~n97 | n564);
  assign n566 = ~i_15_ | n1332;
  assign n567 = n1257 | n1371;
  assign n568 = n566 & n567;
  assign n569 = (n568 | ~n571) & (~n113 | n474);
  assign n570 = ~n879 & (n116 | n165 | n381);
  assign n571 = ~n1233 & n1256;
  assign n572 = ~n1028 & (n346 | n571);
  assign n573 = (~n116 | n984) & (~n165 | n528);
  assign n574 = n1403 & n848 & n851 & n1402;
  assign n575 = (~n321 | n592) & (~n404 | n504);
  assign n576 = (n323 | n1125) & (~n253 | n1377);
  assign n577 = n2138 & n2137 & n2136 & n1743 & n1130 & ~n572 & n1079;
  assign n578 = n2134 & n1650 & n1852 & n1654 & n2135 & n1809 & n1824 & n1751;
  assign n579 = n2128 & n1741 & n1119 & n1733 & n2129 & n1688 & n1707 & n1708;
  assign n580 = n2121 & n2124 & n1542 & n1527 & n725 & n723 & n2122 & n2123;
  assign n581 = n580 & n579 & n578 & n577 & n576 & n575 & n573 & n574;
  assign n582 = ~n291 & (~n729 | ~n1405);
  assign n583 = n381 & (~n316 | ~n1377 | ~n1406);
  assign n584 = (n287 | ~n294) & (~n348 | n442);
  assign n585 = n2211 & (~n404 | n1756);
  assign n586 = n2208 & n2209 & (~n113 | n2210);
  assign n587 = n2206 & n2207 & n1071 & n1531 & n1691 & n1834 & n1792 & n1816;
  assign n588 = n2214 & n486 & n484 & n502 & n498 & n549 & n558 & n1414;
  assign n589 = n2213 & n581 & n1411 & n477 & n421 & n403;
  assign n590 = n589 & n588 & n587 & n586 & n584 & n585;
  assign n591 = ~n98 | n685;
  assign n592 = n1265 | n1371;
  assign n593 = n591 & (~n98 | n592);
  assign n594 = n593 & (~n98 | n305);
  assign n595 = ~n96 | n1377;
  assign n596 = ~n96 | n500;
  assign n597 = n1204 | n1258;
  assign n598 = n595 & n596 & (~n96 | n597);
  assign n599 = ~n163 | n1377;
  assign n600 = ~n163 | n500;
  assign n601 = n599 & n600 & (~n163 | n597);
  assign n602 = ~n96 | n523;
  assign n603 = ~n96 | n566;
  assign n604 = n1204 | n1257;
  assign n605 = n602 & n603 & (~n96 | n604);
  assign n606 = ~n163 | n523;
  assign n607 = ~n163 | n566;
  assign n608 = n606 & n607 & (~n163 | n604);
  assign n609 = ~n167 | n528;
  assign n610 = n1204 | n1246;
  assign n611 = n609 & (~n167 | n610);
  assign n612 = (~n167 | n1377) & (~n571 | n1141);
  assign n613 = n2227 & (~n343 | n652);
  assign n614 = n613 & n612 & n581;
  assign n615 = ~n97 | n361;
  assign n616 = ~n97 | n1373;
  assign n617 = n1204 | n1206;
  assign n618 = n615 & n616 & (~n97 | n617);
  assign n619 = ~n97 | n685;
  assign n620 = ~n97 | n592;
  assign n621 = n619 & n620 & (~n97 | n305);
  assign n622 = ~n96 | n526;
  assign n623 = ~n96 | n1138;
  assign n624 = n622 & n623 & (~n96 | n265);
  assign n625 = ~n96 | n653;
  assign n626 = n625 & (~n96 | n305);
  assign n627 = ~n113 | n777;
  assign n628 = n137 & n1461 & n1452;
  assign n629 = n489 & n1415;
  assign n630 = n627 & n628 & (~n107 | n629);
  assign n631 = n798 & n654 & n752;
  assign n632 = n631 & n264 & n204;
  assign n633 = n96 | n107;
  assign n634 = ~n738 & (n633 | ~n907);
  assign n635 = ~n96 | n2372;
  assign n636 = ~n96 | n629;
  assign n637 = ~n278 | n654;
  assign n638 = n1209 | ~n1388;
  assign n639 = ~n278 | n777;
  assign n640 = n2220 & n2219 & n2217 & n2218;
  assign n641 = n2216 & n2215 & n1519 & n1513 & n1497 & n1478 & ~n103 & n1467;
  assign n642 = n2225 & n2226 & n630 & n1420 & n1422 & n624 & n618 & n621;
  assign n643 = n642 & n641 & n640 & n639 & n638 & n637 & n635 & n636;
  assign n644 = ~n98 | n1138;
  assign n645 = ~n98 | n984;
  assign n646 = n644 & n645 & (~n98 | n265);
  assign n647 = ~n404 | n500;
  assign n648 = n647 & (~n105 | ~n404);
  assign n649 = n500 & n566;
  assign n650 = ~n571 | n649;
  assign n651 = n1258 | n1376;
  assign n652 = n1176 & n1373;
  assign n653 = n1260 | n1376;
  assign n654 = n1257 | n1376;
  assign n655 = n361 & n654 & n653 & n652 & n518 & n651;
  assign n656 = n1245 | n1258;
  assign n657 = n1415 & ~n1114 & n1331;
  assign n658 = n526 & n265;
  assign n659 = n658 & n657 & n656 & ~n105 & n362;
  assign n660 = n313 & n656 & n447 & n468 & n195 & n190;
  assign n661 = ~n98 | n684;
  assign n662 = ~n98 | n1028;
  assign n663 = n661 & n662 & (~n98 | n306);
  assign n664 = n597 & n610 & n306 & n265;
  assign n665 = ~n97 | n684;
  assign n666 = ~n97 | n1028;
  assign n667 = ~n97 | n984;
  assign n668 = n2027 & (~n97 | n664);
  assign n669 = n1427 & n1428;
  assign n670 = n1426 & n1425 & n1423 & n1424;
  assign n671 = ~n98 | n597;
  assign n672 = n671 & n670 & n669 & n663 & n668 & n667 & n665 & n666;
  assign n673 = n288 | n675;
  assign n674 = n1204 | n1260;
  assign n675 = n1214 | ~n1239;
  assign n676 = n673 & (n674 | n675);
  assign n677 = n592 & n1028;
  assign n678 = n507 & n676 & (n677 | ~n928);
  assign n679 = ~n738 & (n344 | n453);
  assign n680 = ~n359 & n911;
  assign n681 = n680 & ~n346 & ~n98 & n291;
  assign n682 = n1219 | n1376;
  assign n683 = n488 & n493 & (~n167 | n682);
  assign n684 = n1221 | n1263;
  assign n685 = n1221 | n1265;
  assign n686 = n684 & n685;
  assign n687 = n329 & n204 & n1247;
  assign n688 = n1245 | n1246;
  assign n689 = n330 & n688 & n687 & n264;
  assign n690 = n359 & (~n190 | ~n1429);
  assign n691 = n165 & (~n523 | ~n1377);
  assign n692 = n107 & (~n500 | ~n1247);
  assign n693 = ~n292 & (~n362 | ~n752 | ~n1382);
  assign n694 = (~n96 | n521) & (~n253 | n910);
  assign n695 = n2253 & (~n278 | n1378);
  assign n696 = n425 & n1005 & (~n113 | n1086);
  assign n697 = n696 & n695 & n439 & n694 & n683 & n558;
  assign n698 = n227 | n1234;
  assign n699 = n822 | n1234;
  assign n700 = n474 | n1234;
  assign n701 = n879 | n1234;
  assign n702 = n875 | n1234;
  assign n703 = n1207 | n1234;
  assign n704 = n226 | n1234;
  assign n705 = n1645 & (n462 | n1234);
  assign n706 = n705 & n704 & n703 & n702 & n701 & n700 & n698 & n699;
  assign n707 = n1243 | n1258;
  assign n708 = n441 & n393 & n473 & n707 & n536;
  assign n709 = n1197 | n1243;
  assign n710 = n472 & n709;
  assign n711 = n227 | n713;
  assign n712 = ~n136 | ~n1213;
  assign n713 = ~n1213 | n1232;
  assign n714 = n711 & n712 & (n713 | ~n716);
  assign n715 = n178 & ~n1232;
  assign n716 = n819 | ~n481 | ~n757;
  assign n717 = n715 & (~n227 | n716);
  assign n718 = ~n98 | n1341;
  assign n719 = n2192 & n1276 & n1344;
  assign n720 = n755 & n793;
  assign n721 = n718 & n719 & (~n98 | n720);
  assign n722 = ~n98 | n392;
  assign n723 = ~n98 | n523;
  assign n724 = ~n98 | n566;
  assign n725 = ~n98 | n567;
  assign n726 = n202 & (~n98 | n604);
  assign n727 = n484 & n726 & n725 & n724 & n722 & n723;
  assign n728 = ~n98 | n536;
  assign n729 = n1334 & n688;
  assign n730 = n728 & (~n98 | n729);
  assign n731 = ~n97 | n879;
  assign n732 = n731 & (~n97 | n470);
  assign n733 = ~n97 | n1335;
  assign n734 = ~n97 | n682;
  assign n735 = n733 & n734 & (~n97 | n266);
  assign n736 = ~n98 | n266;
  assign n737 = ~n98 | n334;
  assign n738 = n1265 | n1376;
  assign n739 = n1198 | n1260;
  assign n740 = (~n98 | n739) & (~n348 | n738);
  assign n741 = ~n97 | n530;
  assign n742 = ~n98 | n1797;
  assign n743 = ~n97 | n440;
  assign n744 = n740 & (~n97 | n774);
  assign n745 = n1457 & n732;
  assign n746 = n1466 & n1465 & n1464 & n1462 & n1463;
  assign n747 = n737 & n1461 & n1460 & n1459 & n1458 & n1434 & n513;
  assign n748 = n747 & n746 & n745 & n730 & n744 & n743 & n741 & n742;
  assign n749 = n1198 | n1219;
  assign n750 = ~n348 | n749;
  assign n751 = n750 & n1435 & n1471 & n1470 & n1469 & n1467 & n1468;
  assign n752 = n1197 | n1376;
  assign n753 = n751 & (~n98 | n752);
  assign n754 = ~n98 | n651;
  assign n755 = n1198 | n1238;
  assign n756 = n514 & n754 & (~n97 | n755);
  assign n757 = n1446 & n822 & n462;
  assign n758 = n757 | ~n1473;
  assign n759 = n1151 & n1250;
  assign n760 = (~n96 | n759) & (~n163 | n752);
  assign n761 = n309 & n1247;
  assign n762 = n1262 & n204;
  assign n763 = n330 & n313 & n761 & n762;
  assign n764 = n1477 & n1476 & n1474 & n1475;
  assign n765 = n1383 & n208 & n872 & n869 & n223 & n870;
  assign n766 = n1352 & n1351 & ~n449 & n1350;
  assign n767 = n1340 & n314 & n298;
  assign n768 = n2271 & n205 & n215 & n1928 & n834 & n1955 & n1626 & n852;
  assign n769 = n768 & n767 & n766 & n466 & n765 & n574 & n764 & n672;
  assign n770 = ~n97 | n392;
  assign n771 = ~n97 | n523;
  assign n772 = n770 & n771 & (~n97 | n604);
  assign n773 = n98 & (~n610 | ~n777);
  assign n774 = n1198 | n1241;
  assign n775 = ~n98 | n774;
  assign n776 = ~n96 | n530;
  assign n777 = n1246 | n1376;
  assign n778 = n776 & (~n96 | (n440 & n777));
  assign n779 = ~n163 | n440;
  assign n780 = n779 & (~n163 | n777);
  assign n781 = ~n359 | n739;
  assign n782 = ~n96 | n1097;
  assign n783 = ~n96 | n540;
  assign n784 = (~n96 | n738) & (~n163 | n1097);
  assign n785 = n780 & n784 & n783 & n782 & n781 & n512;
  assign n786 = ~n163 | n1155;
  assign n787 = ~n163 | n951;
  assign n788 = n786 & n787 & (~n163 | n651);
  assign n789 = n1417 & n924;
  assign n790 = ~n98 | n789;
  assign n791 = ~n96 | n1341;
  assign n792 = ~n96 | n522;
  assign n793 = n1263 | n1376;
  assign n794 = n791 & n792 & (~n96 | n793);
  assign n795 = n163 & (~n1224 | ~n1506);
  assign n796 = n163 & (~n654 | ~n749 | ~n1507);
  assign n797 = ~n96 | n749;
  assign n798 = n1201 | n1376;
  assign n799 = n798 & n738 & n540 & n313 & ~n102 & n191;
  assign n800 = n359 & (~n190 | ~n1166);
  assign n801 = n1505 & n255 & n1073;
  assign n802 = n1532 & n1537 & n1526 & n1521 & n1518;
  assign n803 = n2270 & n1951 & n1516 & n1436 & n1278 & n1195 & ~n103 & ~n164;
  assign n804 = n2269 & n244 & n1915 & n1275 & n1959 & n1345 & n1313 & n1273;
  assign n805 = n2268 & n2154 & n2089 & n2038 & n1991 & n1891 & ~n101 & n231;
  assign n806 = n805 & n804 & n803 & n802 & n788 & n785 & n778 & n801;
  assign n807 = n1553 & n1552 & n1551 & n1550 & n1549 & n1547 & n1548;
  assign n808 = n1546 & n1545 & n366 & n232 & n241 & n1544;
  assign n809 = n505 & (~n96 | n1867);
  assign n810 = n1543 & n1542 & n1541 & n1540 & n1539 & n1538 & n1329 & n601;
  assign n811 = n810 & n809 & n807 & n808;
  assign n812 = n96 & (~n682 | ~n1415);
  assign n813 = n163 & (~n305 | ~n774 | ~n1415);
  assign n814 = n266 | ~n359;
  assign n815 = n1611 & n1610 & n1609 & n1596 & n806 & n1588 & n1578 & n836;
  assign n816 = i_7_ | i_6_;
  assign n817 = n815 & (n816 | ~n1608);
  assign n818 = n179 & ~n1232;
  assign n819 = ~n879 | ~n1207;
  assign n820 = n818 & (~n227 | ~n757 | n819);
  assign n821 = n227 | ~n1619;
  assign n822 = n1220 | n1249;
  assign n823 = n822 | ~n1628;
  assign n824 = n474 | ~n897;
  assign n825 = n902 & ~n1473;
  assign n826 = n700 & n824 & (n825 | n474);
  assign n827 = ~n97 | n317;
  assign n828 = n220 & (~n98 | n263);
  assign n829 = n1563 & n1562 & n1560 & n1561;
  assign n830 = n1559 & n1558 & n1557 & n621;
  assign n831 = n427 & n593 & n830 & n829 & n828 & n827 & n193 & n194;
  assign n832 = ~n97 | n536;
  assign n833 = n832 & (~n97 | n729);
  assign n834 = ~n97 | n1157;
  assign n835 = ~n97 | n1797;
  assign n836 = n1582 & n1581 & n1580 & n368 & n240 & n235 & n1579 & n234;
  assign n837 = n1578 & n2228 & (~n163 | n774);
  assign n838 = n837 & n836 & n833 & n835 & n636 & n491 & n488 & n834;
  assign n839 = ~n97 | n529;
  assign n840 = ~n97 | n528;
  assign n841 = n839 & n840 & (~n97 | n610);
  assign n842 = ~n96 | n1375;
  assign n843 = n842 & (~n96 | n759);
  assign n844 = n97 & (~n265 | ~n845);
  assign n845 = n1201 | n1245;
  assign n846 = ~n98 | n845;
  assign n847 = ~n97 | n1336;
  assign n848 = ~n97 | n1377;
  assign n849 = n847 & n848 & (~n97 | n597);
  assign n850 = ~n98 | n1336;
  assign n851 = ~n98 | n1377;
  assign n852 = ~n98 | n1261;
  assign n853 = n210 & (~n98 | n597);
  assign n854 = n562 & n498 & n670 & n849 & n853 & n852 & n850 & n851;
  assign n855 = n1453 & n1451 & n1452;
  assign n856 = n756 & n1472 & n1312;
  assign n857 = n721 & n1450 & (~n98 | n752);
  assign n858 = ~n97 | n2369;
  assign n859 = n508 | ~n897;
  assign n860 = ~n97 | n474;
  assign n861 = n1858 & n1616 & (n888 | n508);
  assign n862 = n861 & n860 & n859 & n858 & n857 & n856 & n751 & n855;
  assign n863 = ~n136 | n1441;
  assign n864 = ~n136 | n1364;
  assign n865 = (~n136 | ~n159) & (n459 | n875);
  assign n866 = n865 & n863 & n864;
  assign n867 = ~n122 | n1364;
  assign n868 = n867 & (~n122 | ~n159);
  assign n869 = ~n97 | n1330;
  assign n870 = ~n97 | n504;
  assign n871 = n869 & n870 & (~n97 | n306);
  assign n872 = ~n97 | n288;
  assign n873 = n473 & n447;
  assign n874 = n872 & (~n97 | n873);
  assign n875 = i_15_ | n1218;
  assign n876 = n875 | n825;
  assign n877 = n163 & (~n266 | ~n305 | ~n752);
  assign n878 = ~n481 & (n818 | ~n1234);
  assign n879 = n1204 | n1219;
  assign n880 = n459 & n902;
  assign n881 = n879 | n880;
  assign n882 = ~n159 | n1251;
  assign n883 = n1251 | n1364;
  assign n884 = n882 & n883 & (n226 | n459);
  assign n885 = n816 | n1364;
  assign n886 = n885 & (~n159 | n816);
  assign n887 = n444 | ~n897;
  assign n888 = n1235 & ~n1628;
  assign n889 = n887 & (n888 | n444);
  assign n890 = n1355 & n1442 & n2118;
  assign n891 = n704 & n890 & (n825 | n226);
  assign n892 = n703 & n1356 & n1444 & n1367 & n1613;
  assign n893 = (n880 | n1207) & (n1235 | n481);
  assign n894 = n893 & n891 & n889 & n884 & n892 & n886;
  assign n895 = n1645 & n712 & n1368;
  assign n896 = n458 & (~n1608 | (~n136 & n816));
  assign n897 = n1213 & ~n1233;
  assign n898 = ~n713 | n715;
  assign n899 = n2267 | n2276;
  assign n900 = i_9_ & ~i_10_;
  assign n901 = ~i_9_ & i_10_;
  assign n902 = n713 & ~n1619;
  assign n903 = ~n819 | n902;
  assign n904 = n826 & n903 & n1641 & n892;
  assign n905 = n868 & n2287 & (~n899 | ~n901);
  assign n906 = n905 & n904 & ~n132 & n886;
  assign n907 = ~n176 | ~n1239;
  assign n908 = n709 & n1335;
  assign n909 = n907 | n908;
  assign n910 = n1219 | n1371;
  assign n911 = n1232 | ~n1239;
  assign n912 = n910 | n911;
  assign n913 = ~n907 & (~n263 | ~n738);
  assign n914 = n738 | n911;
  assign n915 = ~n911 & (~n393 | ~n1102);
  assign n916 = n911 | n688;
  assign n917 = n2135 & n2104 & n2133;
  assign n918 = n777 & n1649;
  assign n919 = n741 & n743 & (~n97 | n774);
  assign n920 = ~n98 | n761;
  assign n921 = n264 & n979;
  assign n922 = ~n97 | n921;
  assign n923 = n1615 & n1614 & n1613 & n758;
  assign n924 = n1198 | n1240;
  assign n925 = n2289 & (n509 | (n1662 & n875));
  assign n926 = n1204 | n1240;
  assign n927 = n676 & n925 & (n926 | n675);
  assign n928 = n177 & n1256;
  assign n929 = n1228 & n1256;
  assign n930 = n165 | n278;
  assign n931 = n930 & (~n685 | ~n1378);
  assign n932 = ~n278 | n979;
  assign n933 = ~n278 | n1207;
  assign n934 = ~n278 | n474;
  assign n935 = n2143 & (~n165 | n474);
  assign n936 = n1196 | ~n1388;
  assign n937 = n2100 & n2157 & n2075 & n1996 & n1877 & n2052;
  assign n938 = n937 & n936 & n935 & n934 & n932 & n933;
  assign n939 = n656 & n1665;
  assign n940 = ~n165 | n939;
  assign n941 = ~i_11_ | ~n900;
  assign n942 = n941 | ~n1379;
  assign n943 = i_11_ | n1202;
  assign n944 = n943 | ~n1379;
  assign n945 = ~n278 | n984;
  assign n946 = ~n278 | n982;
  assign n947 = ~n278 | n845;
  assign n948 = n1995 & (~n278 | (n284 & n983));
  assign n949 = n948 & n947 & n945 & n946;
  assign n950 = ~n278 | n939;
  assign n951 = n1255 | n1371;
  assign n952 = n1162 & n1028 & n1330;
  assign n953 = n651 & n1029;
  assign n954 = n953 & n952 & n684 & n288 & n951;
  assign n955 = n251 | ~n278;
  assign n956 = ~n278 | n1262;
  assign n957 = ~n165 | n499;
  assign n958 = ~n278 | n1341;
  assign n959 = ~n278 | n522;
  assign n960 = n1670 & (~n165 | n954);
  assign n961 = n2291 & (~n278 | (n204 & n793));
  assign n962 = n2290 & n638 & n1949 & n1994 & n1931 & n1874 & n2050 & n2098;
  assign n963 = n962 & n961 & n960 & n959 & n958 & n957 & n955 & n956;
  assign n964 = n313 & n334;
  assign n965 = n682 & n653 & n263 & n1676;
  assign n966 = n739 & n789 & n964 & n965;
  assign n967 = n1125 & ~n450 & n979;
  assign n968 = n1335 & n1247 & n1373 & n1678 & n331 & n1102;
  assign n969 = n774 & n777;
  assign n970 = n329 & n317 & n495;
  assign n971 = n970 & n793 & n798 & n969 & n968 & n967 & n657 & n525;
  assign n972 = n1697 & n1696 & n1695 & n1694 & n1693 & n1692 & n1691 & n942;
  assign n973 = n944 & n1690 & n1689 & n1688 & n1687 & n1685 & n1686;
  assign n974 = n1705 & n1704 & n1703 & n1702 & n1701 & n1700 & n1698 & n1699;
  assign n975 = n1713 & n1712 & n1711 & n1710 & n1709 & n1708 & n1706 & n1707;
  assign n976 = n1721 & n1002 & n1730 & n1726;
  assign n977 = n2298 & n2296 & n1936 & n1914 & n1684 & n963 & ~n166 & n949;
  assign n978 = n2294 & n2295 & n1999 & n1913 & n2079 & n1998 & n1927 & n1937;
  assign n979 = n1219 | n1243;
  assign n980 = ~n116 | n979;
  assign n981 = ~n116 | n287;
  assign n982 = n798 & n1374 & n1224;
  assign n983 = n1666 & n875 & n441;
  assign n984 = n1201 | n1371;
  assign n985 = n984 & n284 & n982 & n983;
  assign n986 = ~n116 | n227;
  assign n987 = ~n120 & n986 & (~n116 | n985);
  assign n988 = ~n353 | n926;
  assign n989 = ~n353 | n430;
  assign n990 = ~n353 | ~n450;
  assign n991 = n2162 & n2077 & n2161;
  assign n992 = n1742 & n1741 & n1740 & n1739 & n1738 & n1737 & n1736 & n980;
  assign n993 = n1735 & n1734 & n1733 & n1732 & ~n117 & n981;
  assign n994 = (~n116 | n1144) & (~n353 | n1677);
  assign n995 = n987 & n994 & n993 & n992 & n991 & n990 & n988 & n989;
  assign n996 = ~n167 | n567;
  assign n997 = ~n167 | n1157;
  assign n998 = ~n167 | n566;
  assign n999 = ~n167 | n508;
  assign n1000 = ~n167 | n529;
  assign n1001 = n1744 & n270 & n1743;
  assign n1002 = n1722 & n537;
  assign n1003 = n384 & n1440 & (~n167 | n982);
  assign n1004 = n1003 & n1002 & n1001 & n1000 & n999 & n998 & n996 & n997;
  assign n1005 = ~n167 | n393;
  assign n1006 = ~n167 | n1139;
  assign n1007 = ~n167 | n1138;
  assign n1008 = ~n167 | n984;
  assign n1009 = (~n381 | n658) & (~n404 | n982);
  assign n1010 = n1969 & n1997 & n1919 & n2059 & n1878 & n1901 & n1117 & n1879;
  assign n1011 = n1010 & n1004 & n1009 & n1008 & n1007 & n1005 & n1006;
  assign n1012 = n1250 & n1104;
  assign n1013 = ~n404 | n1012;
  assign n1014 = ~n167 | n474;
  assign n1015 = ~n167 | n979;
  assign n1016 = ~n167 | n495;
  assign n1017 = ~n170 & (~n381 | n2297);
  assign n1018 = ~n404 | n654;
  assign n1019 = n1899 & n2062 & n1884 & n1939 & n2165 & n1882;
  assign n1020 = n1019 & n1018 & n1017 & n1016 & n1014 & n1015;
  assign n1021 = ~n167 | n442;
  assign n1022 = n1021 & (~n167 | (n330 & n527));
  assign n1023 = ~n167 | n707;
  assign n1024 = n2096 & n1905 & n2058;
  assign n1025 = n1023 & n1024 & (~n105 | ~n167);
  assign n1026 = n684 & n1418;
  assign n1027 = n288 & n873;
  assign n1028 = n1263 | n1371;
  assign n1029 = n1341 & n522;
  assign n1030 = n1029 & n1028 & n204 & n1027 & n1026 & n720;
  assign n1031 = n1748 & n1747 & n1745 & n1746;
  assign n1032 = n1754 & n1753 & n1752 & n1751 & n1749 & n1750;
  assign n1033 = n1956 & n1965 & (~n404 | n1030);
  assign n1034 = n1279 & n1342 & n2132;
  assign n1035 = n2299 & n1881 & n1933 & n1906 & n1880 & n2060;
  assign n1036 = n1035 & n1034 & n1033 & n1022 & n1032 & n1031 & n1025 & n648;
  assign n1037 = n381 & (~n964 | ~n1678);
  assign n1038 = ~n774 | ~n329 | ~n604;
  assign n1039 = n404 & (~n918 | n1038 | ~n1756);
  assign n1040 = ~n176 | n1230;
  assign n1041 = n1214 | n1230;
  assign n1042 = n1040 & n1041;
  assign n1043 = ~n105 & n1336;
  assign n1044 = ~n571 | n1043;
  assign n1045 = n107 & (~n500 | ~n1665);
  assign n1046 = n331 & n951 & n1155;
  assign n1047 = ~n104 | n1046;
  assign n1048 = ~n113 | n1080;
  assign n1049 = ~n278 | n610;
  assign n1050 = n778 & (~n107 | n2307);
  assign n1051 = n1050 & n1049 & n1048 & n919 & ~n115 & n538;
  assign n1052 = n346 & (~n1247 | ~n1415);
  assign n1053 = n1490 & n1489 & n1488 & n1487 & n1486 & n1485 & ~n773 & n1484;
  assign n1054 = n1289 & n1287 & n1288;
  assign n1055 = (~n404 | n2307) & (~n571 | n1795);
  assign n1056 = n2309 & (~n104 | (n529 & n1136));
  assign n1057 = n1804 & n1051 & n1802 & n838 & n138 & n1783 & n972;
  assign n1058 = n2308 & n2231 & n2167 & n2083 & n1722 & n1679 & n997 & ~n1052;
  assign n1059 = n1058 & n1057 & n1056 & n1055 & n1054 & n630 & n1053 & n730;
  assign n1060 = n104 & (~n447 | ~n1026 | ~n1381);
  assign n1061 = ~n107 | n522;
  assign n1062 = (~n104 | n953) & (n720 | n1292);
  assign n1063 = n1062 & n416 & n1061;
  assign n1064 = n104 & (~n1336 | ~n1664);
  assign n1065 = n113 & (~n331 | ~n755);
  assign n1066 = n571 & (~n651 | ~n755 | ~n951);
  assign n1067 = n571 & (~n206 | ~n952 | ~n1026);
  assign n1068 = n107 & (~n206 | ~n1027 | ~n1330);
  assign n1069 = ~n113 | n1043;
  assign n1070 = ~n107 | n1026;
  assign n1071 = ~n113 | n2374;
  assign n1072 = n1854 & n255 & (n1292 | n1162);
  assign n1073 = n1499 & n1497 & n1498;
  assign n1074 = ~n1067 & ~n1068 & (~n165 | n793);
  assign n1075 = n2306 & n1063 & n1169 & n1823 & n1180 & n1812;
  assign n1076 = n1075 & n1074 & n756 & n1073 & n1072 & n1071 & n1069 & n1070;
  assign n1077 = n738 & n739;
  assign n1078 = n489 | ~n571;
  assign n1079 = ~n571 | n1372;
  assign n1080 = n529 & n1415;
  assign n1081 = n1078 & n1079 & (~n571 | n1080);
  assign n1082 = n1221 | n1260;
  assign n1083 = n1082 & n287 & ~n109 & n219;
  assign n1084 = n471 & n674 & n426;
  assign n1085 = n263 & n653 & n356;
  assign n1086 = n287 & n1082;
  assign n1087 = n685 & n592;
  assign n1088 = n1087 & n1086 & n1085 & n1084 & n317;
  assign n1089 = ~n113 | n685;
  assign n1090 = ~n113 | n592;
  assign n1091 = ~n113 | n317;
  assign n1092 = (~n113 | n1083) & (~n571 | n1088);
  assign n1093 = n1957 & n2145 & n1280 & n2030 & n2180 & n2142;
  assign n1094 = n1093 & n1081 & n1092 & n1091 & n1089 & n1090;
  assign n1095 = ~n113 | n951;
  assign n1096 = n1095 & (~n113 | n651);
  assign n1097 = n1220 | n1265;
  assign n1098 = n739 & n1097 & n195;
  assign n1099 = ~n653 & (n381 | n930);
  assign n1100 = ~n107 | n470;
  assign n1101 = n1887 & n2068 & n2102;
  assign n1102 = n392 & n508;
  assign n1103 = ~n169 & n1101 & (~n107 | n1102);
  assign n1104 = n1151 & n1375;
  assign n1105 = n1243 | n1249;
  assign n1106 = n1105 & n1104 & n329 & n822 & n654;
  assign n1107 = ~n104 | n1331;
  assign n1108 = ~n104 | n444;
  assign n1109 = (~n104 | n1106) & (~n107 | n654);
  assign n1110 = n2136 & n1946 & n2230 & n2223 & n2311 & n1916 & n2166;
  assign n1111 = n1110 & n1103 & n1109 & n1108 & n396 & n1107;
  assign n1112 = n1105 & n201;
  assign n1113 = ~n1114 & n1112 & n467 & n1102;
  assign n1114 = ~n523 | ~n604;
  assign n1115 = n571 & (~n392 | ~n822 | n1114);
  assign n1116 = n329 & ~n1114;
  assign n1117 = ~n167 | n1105;
  assign n1118 = ~n167 | n329;
  assign n1119 = ~n278 | n523;
  assign n1120 = (~n346 | n1116) & (n1102 | n1290);
  assign n1121 = ~n166 & ((~n107 & ~n571) | n1104);
  assign n1122 = n1616 & n1430 & n2156 & n2081 & n1681 & n996 & n1680 & n998;
  assign n1123 = n2323 & n1111 & n1779 & n1181 & n139 & n1675 & n1001 & n973;
  assign n1124 = n1123 & n1122 & n1121 & n1120 & n1119 & n1118 & n225 & n1117;
  assign n1125 = n1197 | n1371;
  assign n1126 = n1125 & n1028;
  assign n1127 = n116 | n253;
  assign n1128 = (~n749 | ~n752) & (~n327 | n1127);
  assign n1129 = ~n682 & (n321 | n930);
  assign n1130 = ~n104 | n526;
  assign n1131 = ~n104 | n1138;
  assign n1132 = ~n104 | n845;
  assign n1133 = n1823 & (~n104 | (n875 & n1224));
  assign n1134 = n507 & n2168 & n2224 & n2144 & n1922 & n2137 & n1889 & n2067;
  assign n1135 = n1134 & n1133 & n1132 & n434 & n413 & n1131 & n395 & n1130;
  assign n1136 = n1797 & n1157 & n1796;
  assign n1137 = ~n571 | n1136;
  assign n1138 = ~i_15_ | n1225;
  assign n1139 = n472 & n875 & n845;
  assign n1140 = n1139 & n1138 & n984;
  assign n1141 = n499 & n567;
  assign n1142 = n226 & n526 & n1141 & n441;
  assign n1143 = n525 & ~n450 & n191 & ~n268;
  assign n1144 = n879 & n1147;
  assign n1145 = n1206 | n1220;
  assign n1146 = n361 & n1145 & n1144 & n658;
  assign n1147 = n313 & n1152 & n752 & n1731 & n263 & n1676;
  assign n1148 = n1147 & n658 & n685;
  assign n1149 = n1866 & n1224 & n1166 & n738 & ~n99 & n631;
  assign n1150 = n953 & n474 & n251 & n1149 & n1085 & n720;
  assign n1151 = n1220 | n1257;
  assign n1152 = n1197 | n1220;
  assign n1153 = n447 & n1152 & n1151 & n333 & n316 & n313;
  assign n1154 = n426 & n738;
  assign n1155 = n1220 | n1258;
  assign n1156 = n284 & n265 & n227;
  assign n1157 = n1220 | n1241;
  assign n1158 = n1248 & n1334 & n951;
  assign n1159 = n1158 & n1157 & n1156 & n1155 & n969 & n968 & n309 & ~n450;
  assign n1160 = n334 & n749;
  assign n1161 = n752 & n1507;
  assign n1162 = n251 & n762;
  assign n1163 = n1250 & n1374 & n610 & n688 & n489 & n313;
  assign n1164 = n1163 & n1162 & n1161 & n1160 & n798 & n979;
  assign n1165 = n1868 & n1867 & n1104 & n430 & n319 & ~n268 & n198 & n206;
  assign n1166 = n789 & n521 & n1145;
  assign n1167 = n1166 & n1165 & n873 & n195 & n361;
  assign n1168 = n1833 & n1832 & n1831 & n1830 & n1829 & n1828 & ~n110 & n1827;
  assign n1169 = n1826 & n1825 & ~n1060 & n1824;
  assign n1170 = n1853 & n1852 & n1851 & n1850 & n1849 & n1848 & n1847 & n1100;
  assign n1171 = n1063 & n1808 & n1802;
  assign n1172 = n534 & n1790 & (~n104 | n1159);
  assign n1173 = n2364 & n2365 & n2169 & n1267 & n1266 & n433 & n2087 & n1921;
  assign n1174 = n1173 & n1172 & n1171 & n1170 & n1135 & n1111 & n1168 & n1169;
  assign n1175 = n1335 & n682;
  assign n1176 = n1240 | n1376;
  assign n1177 = n227 & n1250 & n540;
  assign n1178 = n1507 & n952 & n967 & n969 & n1795 & n1165 & n1870 & n1869;
  assign n1179 = n1178 & n1177 & n926 & n504 & n1176 & n191 & n1175 & n1097;
  assign n1180 = n1818 & n1817 & n1816 & n1815 & n1814 & ~n114 & n1813;
  assign n1181 = n1839 & n1838 & n1837 & n1836 & n1835 & n1834 & n1096 & ~n1115;
  assign n1182 = n1865 & n1855 & n1137 & n1864 & n1863 & n1390;
  assign n1183 = n1846 & n1845 & n1844 & n1843 & n1842 & ~n118 & n414;
  assign n1184 = n1812 & n1794 & n569;
  assign n1185 = n2367 & (~n571 | n1179);
  assign n1186 = n2366 & n1958 & n1942 & n1409 & ~n115 & n1268;
  assign n1187 = n1186 & n1185 & n1184 & n1183 & n1182 & n1181 & n1094 & n1180;
  assign n1188 = ~n96 | n755;
  assign n1189 = ~n163 | n1341;
  assign n1190 = ~n163 | n522;
  assign n1191 = ~n163 | n288;
  assign n1192 = n1512 & n1511 & n1510 & n598 & n1508 & n1509;
  assign n1193 = ~n163 | (n306 & n720);
  assign n1194 = n2149 & n1860 & n1912 & n1954 & n2123 & n2088 & n2041 & n2122;
  assign n1195 = n1194 & n1193 & n794 & n1192 & n1191 & n1190 & n1188 & n1189;
  assign n1196 = i_11_ | ~n901;
  assign n1197 = ~i_15_ | n1196;
  assign n1198 = i_12_ | i_14_ | i_13_;
  assign n1199 = i_12_ | ~i_13_;
  assign n1200 = i_11_ | ~n900;
  assign n1201 = ~i_15_ | n1200;
  assign n1202 = ~i_9_ | ~i_10_;
  assign n1203 = n1202 & n941;
  assign n1204 = ~i_14_ | i_12_ | i_13_;
  assign n1205 = i_11_ | n481;
  assign n1206 = ~i_15_ | n1205;
  assign n1207 = n1197 | n1198;
  assign n1208 = ~i_12_ | n1196;
  assign n1209 = ~i_11_ | ~n901;
  assign n1210 = ~i_12_ | n1200;
  assign n1211 = n1199 & n1204 & n1210 & n1209 & n226 & n1208 & n1207 & n1203;
  assign n1212 = i_3_ | i_5_ | i_4_;
  assign n1213 = n172 & ~n1212;
  assign n1214 = ~i_8_ | n816;
  assign n1215 = i_5_ & ~i_3_ & ~i_4_;
  assign n1216 = i_5_ & ~i_3_ & i_4_;
  assign n1217 = i_15_ | n1200;
  assign n1218 = n1200 | n1204;
  assign n1219 = i_15_ | n1196;
  assign n1220 = i_14_ | n1199;
  assign n1221 = ~i_14_ | n1199;
  assign n1222 = n481 & n1202;
  assign n1223 = n1196 | n1221;
  assign n1224 = n1201 | n1220;
  assign n1225 = n1200 | n1221;
  assign n1226 = n266 & n1209 & n941 & n1208 & n265 & n1210;
  assign n1227 = n1226 & n1225 & n1224 & n1223 & n749 & n1152;
  assign n1228 = ~i_8_ & n136;
  assign n1229 = i_5_ | i_3_ | ~i_4_;
  assign n1230 = ~n172 | n1229;
  assign n1231 = ~n186 & ~n1212;
  assign n1232 = i_8_ | ~n122;
  assign n1233 = i_8_ | n816;
  assign n1234 = n1230 | n1232;
  assign n1235 = n1234 & n459;
  assign n1236 = ~i_5_ & i_3_ & ~i_4_;
  assign n1237 = n172 & n174;
  assign n1238 = i_15_ | n1209;
  assign n1239 = ~n186 & n1216;
  assign n1240 = i_15_ | n1205;
  assign n1241 = i_15_ | n941;
  assign n1242 = ~i_12_ | i_13_;
  assign n1243 = i_14_ | n1242;
  assign n1244 = ~i_12_ | ~i_13_;
  assign n1245 = i_14_ | n1244;
  assign n1246 = ~i_15_ | n941;
  assign n1247 = n1241 | n1245;
  assign n1248 = n1198 | n1246;
  assign n1249 = i_15_ | n943;
  assign n1250 = n1198 | n1249;
  assign n1251 = i_6_ | ~i_7_;
  assign n1252 = ~i_8_ & ~n1251;
  assign n1253 = ~n186 & n1215;
  assign n1254 = ~i_11_ | n1202;
  assign n1255 = i_15_ | n1254;
  assign n1256 = ~n186 & ~n1229;
  assign n1257 = ~i_15_ | n943;
  assign n1258 = ~i_15_ | n1254;
  assign n1259 = ~i_11_ | n481;
  assign n1260 = i_15_ | n1259;
  assign n1261 = n1220 | n1255;
  assign n1262 = n1238 | n1243;
  assign n1263 = ~i_15_ | n1209;
  assign n1264 = i_8_ & ~n1251;
  assign n1265 = ~i_15_ | n1259;
  assign n1266 = ~n107 | n226;
  assign n1267 = ~n107 | n227;
  assign n1268 = ~n113 | n227;
  assign n1269 = n1957 & n1815 & n1826 & n1956;
  assign n1270 = n1955 & n1476 & n1954 & n1953 & n1952 & n1951 & n1949 & n1950;
  assign n1271 = n1270 & n1269 & n1268 & n1267 & n1266 & n228;
  assign n1272 = ~n96 | n1207;
  assign n1273 = ~n96 | n474;
  assign n1274 = n1273 & ~n230 & n1272;
  assign n1275 = ~n96 | n334;
  assign n1276 = ~n97 | n331;
  assign n1277 = ~n97 | n334;
  assign n1278 = ~n96 | n313;
  assign n1279 = ~n167 | n331;
  assign n1280 = ~n113 | n1797;
  assign n1281 = n1958 & n1271 & n1118 & ~n229 & n222 & n224;
  assign n1282 = n1281 & n1280 & n1279 & n1278 & n1277 & n1276 & n485 & n1275;
  assign n1283 = ~n167 | n309;
  assign n1284 = ~n167 | n1247;
  assign n1285 = ~n167 | n1248;
  assign n1286 = n1285 & n1283 & n1284;
  assign n1287 = ~n278 | n309;
  assign n1288 = ~n278 | n1248;
  assign n1289 = ~n278 | n1247;
  assign n1290 = ~n104 & ~n165;
  assign n1291 = ~n116 & ~n278;
  assign n1292 = ~n104 & ~n107;
  assign n1293 = n1204 | n1255;
  assign n1294 = n1293 & n508;
  assign n1295 = n288 & n879;
  assign n1296 = n1908 & (n911 | n508);
  assign n1297 = n1828 & n1907 & n1788 & n1651 & n1753 & n1748;
  assign n1298 = n1904 & n1749 & n1906 & n1905 & n1692 & n1717 & n1671 & n1689;
  assign n1299 = n1892 & n731 & n1893 & n728 & n1626 & n1477 & n1482 & n1560;
  assign n1300 = n1896 & n1599 & n1898 & n1564 & n1589 & n1897 & n1577 & n1570;
  assign n1301 = n1789 & n1820 & n1829 & n1831 & n1888 & n1793 & n1806 & n1887;
  assign n1302 = n1889 & n1851 & n1850 & n1108 & n324 & ~n322 & ~n164 & n320;
  assign n1303 = n1737 & n1735 & n1021 & n986 & n1881 & n1880 & n1878 & n1879;
  assign n1304 = n1886 & n1885 & n1884 & n1883 & n1773 & n1882 & n1777 & n1784;
  assign n1305 = n1504 & n1501 & n1669 & n1875 & n1703 & n1874 & n1872 & n1873;
  assign n1306 = n1693 & n1695 & n1686 & n1877 & n1711 & n1690 & n1876 & n1673;
  assign n1307 = n852 & n1474 & n1871 & n1487 & n1509 & n1451 & n1547 & n1552;
  assign n1308 = n1529 & n1539 & n1590 & n1593 & n1571 & n1572 & n1567 & n1601;
  assign n1309 = ~n116 & ~n294;
  assign n1310 = n617 & n306 & n305;
  assign n1311 = n266 & n1310;
  assign n1312 = ~n98 | n331;
  assign n1313 = ~n163 | n331;
  assign n1314 = ~n571 | n2375;
  assign n1315 = n1890 & (~n165 | n331);
  assign n1316 = n1315 & n1314 & n1312 & n1313;
  assign n1317 = ~n107 | n191;
  assign n1318 = n1922 & n1117 & n1920 & n1921;
  assign n1319 = n1919 & n988 & n1769 & n1918 & n1917 & n1015 & n1825 & n1916;
  assign n1320 = n1912 & n1557 & n1911 & n1544 & n1579 & n1582 & n1585 & n1587;
  assign n1321 = n1603 & n1635 & n1555 & n1915 & n932 & n956 & n1913 & n1914;
  assign n1322 = ~n404 | n442;
  assign n1323 = n330 | ~n404;
  assign n1324 = ~n404 | n527;
  assign n1325 = n1324 & n1322 & n1323;
  assign n1326 = ~n163 | n330;
  assign n1327 = ~n163 | n527;
  assign n1328 = ~n163 | n1261;
  assign n1329 = n1328 & n1326 & n1327;
  assign n1330 = n1221 | n1238;
  assign n1331 = n1245 | n1257;
  assign n1332 = n1221 | n943;
  assign n1333 = n1206 | n1245;
  assign n1334 = n1243 | n1246;
  assign n1335 = i_15_ | n1223;
  assign n1336 = n1221 | n1255;
  assign n1337 = n1206 | n1243;
  assign n1338 = ~n97 | n441;
  assign n1339 = ~n98 | n1330;
  assign n1340 = n1339 & n847 & n850 & n1338;
  assign n1341 = n1220 | n1263;
  assign n1342 = ~n167 | n1155;
  assign n1343 = ~n113 | n1155;
  assign n1344 = ~n97 | n1155;
  assign n1345 = ~n96 | n1224;
  assign n1346 = n1248 & n729;
  assign n1347 = n423 & n1336 & n392;
  assign n1348 = n684 & n1151;
  assign n1349 = ~n165 & ~n321;
  assign n1350 = ~n97 | n472;
  assign n1351 = ~n98 | n472;
  assign n1352 = n448 & (~n97 | (n873 & n1346));
  assign n1353 = ~i_0_ | i_1_;
  assign n1354 = n1229 | n1353;
  assign n1355 = n1251 | n1354;
  assign n1356 = n816 | n1354;
  assign n1357 = ~n136 | n1354;
  assign n1358 = ~n122 | n1354;
  assign n1359 = n1358 & n1357 & n1355 & n1356;
  assign n1360 = n1271 & n2026 & (~n107 | n495);
  assign n1361 = n2024 & n2023 & n2022 & n2021 & ~n456 & ~n457;
  assign n1362 = n2018 & n2016 & n2020 & n1288 & n1791 & n2019 & n1732 & n1322;
  assign n1363 = n2013 & n2005 & n2006 & n1536 & n1857 & n1472 & n619 & n718;
  assign n1364 = n1212 | n1353;
  assign n1365 = n883 & n864 & n867 & n885;
  assign n1366 = n879 | ~n897;
  assign n1367 = ~n897 | n1207;
  assign n1368 = ~n1213 | n1251;
  assign n1369 = n887 & n859 & n1621 & n2118 & n1623 & n1631;
  assign n1370 = n1369 & n482 & n1368 & n1367 & n824 & n1366;
  assign n1371 = ~i_14_ | n1242;
  assign n1372 = n1246 | n1371;
  assign n1373 = n1206 | n1371;
  assign n1374 = n1217 | n1371;
  assign n1375 = n1249 | n1371;
  assign n1376 = ~i_14_ | n1244;
  assign n1377 = n1255 | n1376;
  assign n1378 = n1082 & n674;
  assign n1379 = n1252 & n1253;
  assign n1380 = n529 & n536;
  assign n1381 = n1330 & n288;
  assign n1382 = n526 & n653;
  assign n1383 = n840 & n211 & n839 & n832;
  assign n1384 = ~n98 | n1176;
  assign n1385 = ~n98 | n430;
  assign n1386 = ~n98 | n926;
  assign n1387 = n1386 & n1384 & n1385;
  assign n1388 = n1253 & n1264;
  assign n1389 = ~n107 | n1176;
  assign n1390 = ~n113 | n984;
  assign n1391 = ~n168 & n1845 & (~n278 | n518);
  assign n1392 = n2170 & n1661 & n1660 & n2169 & n2168 & n1008;
  assign n1393 = n1798 & n2165 & n1762 & n1658 & n1827 & n1656;
  assign n1394 = n1765 & n2167 & n1813 & n1848 & n1807 & n2166;
  assign n1395 = n2155 & n2159 & n996 & n2164 & n2163 & n2162 & n2160 & n2161;
  assign n1396 = ~n167 | n536;
  assign n1397 = n406 & n1396 & n385;
  assign n1398 = ~n96 | n875;
  assign n1399 = n387 & n408 & n1398;
  assign n1400 = ~n278 | n508;
  assign n1401 = n407 & n1400 & n386;
  assign n1402 = ~n97 | n526;
  assign n1403 = ~n98 | n504;
  assign n1404 = n447 & n649;
  assign n1405 = n1374 & n1375;
  assign n1406 = n521 & n910 & n653 & n191;
  assign n1407 = n523 & n592 & n984 & n1125 & n528;
  assign n1408 = n685 & n688 & n1138 & n566 & n495;
  assign n1409 = ~n571 | n2376;
  assign n1410 = n2139 & (n474 | ~n571);
  assign n1411 = n1410 & n1409 & n1401 & n1005 & n999 & ~n570 & n384 & n569;
  assign n1412 = n1397 & n2147 & (~n278 | n875);
  assign n1413 = n2141 & n2145 & n1817 & n2144 & n1844 & n2143 & n2142 & n1767;
  assign n1414 = n1413 & n1412 & n565 & n1399 & n562 & n560;
  assign n1415 = n610 & n528;
  assign n1416 = n566 & ~n1114;
  assign n1417 = n1206 | n1376;
  assign n1418 = n504 & n306;
  assign n1419 = ~n278 | n489;
  assign n1420 = n538 & n1419 & n1049;
  assign n1421 = ~n96 | n685;
  assign n1422 = n1421 & n626;
  assign n1423 = ~n98 | n499;
  assign n1424 = ~n98 | n500;
  assign n1425 = ~n97 | n499;
  assign n1426 = ~n97 | n500;
  assign n1427 = ~n97 | n489;
  assign n1428 = ~n97 | n1372;
  assign n1429 = n793 & n752;
  assign n1430 = n1293 | n509;
  assign n1431 = ~n929 | n1372;
  assign n1432 = (n509 | n536) & (n499 | ~n929);
  assign n1433 = n1432 & n1431 & n1430 & n678 & ~n679;
  assign n1434 = ~n98 | n798;
  assign n1435 = ~n98 | n654;
  assign n1436 = ~n163 | n1666;
  assign n1437 = (~n343 | n654) & (n327 | n798);
  assign n1438 = n1437 & n646 & n648 & n650 & n1436 & n1435 & n754 & n1434;
  assign n1439 = ~n167 | n489;
  assign n1440 = n1439 & n611;
  assign n1441 = ~n1216 | n1353;
  assign n1442 = n1251 | n1441;
  assign n1443 = ~n122 | n1441;
  assign n1444 = n816 | n1441;
  assign n1445 = n1444 & n1442 & n1443;
  assign n1446 = n474 & n226 & n875;
  assign n1447 = ~n97 | n793;
  assign n1448 = ~n97 | n522;
  assign n1449 = ~n97 | n1341;
  assign n1450 = n1449 & n1447 & n1448;
  assign n1451 = ~n98 | n822;
  assign n1452 = ~n97 | n651;
  assign n1453 = ~n97 | n951;
  assign n1454 = n1450 & n721;
  assign n1455 = n855 & n860 & n727 & n1454;
  assign n1456 = n2120 & n1953 & n2045 & n2119 & n2044 & n1893 & n1871 & n2148;
  assign n1457 = n1456 & n736 & n735 & n560 & n364 & n222 & ~n162 & n199;
  assign n1458 = ~n97 | n1145;
  assign n1459 = ~n97 | n924;
  assign n1460 = ~n98 | n1224;
  assign n1461 = ~n97 | n777;
  assign n1462 = ~n98 | n540;
  assign n1463 = ~n98 | n1097;
  assign n1464 = ~n97 | n540;
  assign n1465 = ~n97 | n1097;
  assign n1466 = ~n97 | n739;
  assign n1467 = ~n97 | n752;
  assign n1468 = ~n97 | n910;
  assign n1469 = ~n98 | n910;
  assign n1470 = ~n98 | n1152;
  assign n1471 = ~n97 | n1152;
  assign n1472 = ~n98 | n1155;
  assign n1473 = n179 & ~n1233;
  assign n1474 = ~n98 | n251;
  assign n1475 = ~n97 | n251;
  assign n1476 = ~n97 | n1261;
  assign n1477 = ~n98 | n288;
  assign n1478 = ~n97 | n654;
  assign n1479 = ~n97 | n1375;
  assign n1480 = ~n98 | n526;
  assign n1481 = ~n98 | n441;
  assign n1482 = ~n98 | n875;
  assign n1483 = n1482 & n1481 & n1480 & n775 & n1478 & n1479;
  assign n1484 = ~n98 | n489;
  assign n1485 = ~n98 | n440;
  assign n1486 = ~n98 | n1372;
  assign n1487 = ~n98 | n1157;
  assign n1488 = ~n98 | n530;
  assign n1489 = ~n98 | n528;
  assign n1490 = ~n98 | n529;
  assign n1491 = ~n97 | n1151;
  assign n1492 = ~n97 | n1250;
  assign n1493 = ~n97 | n567;
  assign n1494 = ~n98 | n1151;
  assign n1495 = ~n98 | n1250;
  assign n1496 = n772 & n1495 & n1494 & n365 & n1493 & n1491 & n1492;
  assign n1497 = ~n96 | n651;
  assign n1498 = ~n96 | n951;
  assign n1499 = ~n96 | n1155;
  assign n1500 = ~n163 | n393;
  assign n1501 = ~n163 | n444;
  assign n1502 = ~n163 | n329;
  assign n1503 = ~n163 | n1105;
  assign n1504 = ~n163 | n822;
  assign n1505 = n1504 & n1503 & n1502 & n1500 & n1501;
  assign n1506 = n334 & n1374;
  assign n1507 = n1152 & n910;
  assign n1508 = ~n96 | n707;
  assign n1509 = ~n96 | n442;
  assign n1510 = ~n96 | n1336;
  assign n1511 = ~n96 | n1293;
  assign n1512 = ~n96 | n656;
  assign n1513 = ~n96 | n654;
  assign n1514 = ~n163 | n1151;
  assign n1515 = ~n163 | n1250;
  assign n1516 = n1515 & n1513 & n1514;
  assign n1517 = ~n96 | n1161;
  assign n1518 = n1517 & n797 & n511 & ~n796;
  assign n1519 = ~n96 | n798;
  assign n1520 = ~n96 | n1374;
  assign n1521 = n1520 & ~n795 & n1519;
  assign n1522 = ~n163 | n567;
  assign n1523 = ~n163 | n392;
  assign n1524 = ~n163 | n508;
  assign n1525 = ~n163 | n1331;
  assign n1526 = n608 & n1525 & n1524 & n1522 & n1523;
  assign n1527 = ~n163 | n984;
  assign n1528 = ~n163 | n472;
  assign n1529 = ~n163 | n226;
  assign n1530 = ~n163 | n284;
  assign n1531 = ~n163 | n2371;
  assign n1532 = n1531 & n1530 & n1529 & n1527 & n1528;
  assign n1533 = ~n97 | n1417;
  assign n1534 = ~n97 | n521;
  assign n1535 = ~n98 | n521;
  assign n1536 = ~n98 | n1145;
  assign n1537 = n1536 & n1535 & n1277 & n790 & n1533 & n1534;
  assign n1538 = ~n163 | n707;
  assign n1539 = ~n163 | n442;
  assign n1540 = ~n163 | n1293;
  assign n1541 = ~n163 | n656;
  assign n1542 = ~n163 | n499;
  assign n1543 = ~n163 | n1336;
  assign n1544 = ~n96 | n1262;
  assign n1545 = ~n96 | n473;
  assign n1546 = ~n96 | n206;
  assign n1547 = ~n163 | n206;
  assign n1548 = ~n163 | n204;
  assign n1549 = ~n163 | n447;
  assign n1550 = ~n163 | n473;
  assign n1551 = ~n163 | n1262;
  assign n1552 = ~n163 | n251;
  assign n1553 = ~n96 | n1028;
  assign n1554 = ~n96 | n472;
  assign n1555 = ~n96 | n284;
  assign n1556 = n1399 & n1554 & n1555;
  assign n1557 = ~n97 | n674;
  assign n1558 = ~n97 | n653;
  assign n1559 = ~n97 | n1082;
  assign n1560 = ~n98 | n674;
  assign n1561 = ~n98 | n2368;
  assign n1562 = ~n98 | n653;
  assign n1563 = ~n98 | n1082;
  assign n1564 = ~n96 | n508;
  assign n1565 = ~n96 | n1331;
  assign n1566 = ~n96 | n393;
  assign n1567 = ~n96 | n444;
  assign n1568 = ~n96 | n329;
  assign n1569 = n1568 & n1567 & n1566 & n1564 & n1565;
  assign n1570 = ~n163 | n309;
  assign n1571 = ~n163 | n1157;
  assign n1572 = ~n163 | n1248;
  assign n1573 = ~n163 | n1247;
  assign n1574 = ~n163 | n688;
  assign n1575 = ~n163 | n1334;
  assign n1576 = ~n163 | n529;
  assign n1577 = ~n163 | n536;
  assign n1578 = n1577 & n1576 & n1575 & n1574 & n1573 & n1572 & n1570 & n1571;
  assign n1579 = ~n96 | n309;
  assign n1580 = ~n96 | n1334;
  assign n1581 = ~n96 | n529;
  assign n1582 = ~n96 | n536;
  assign n1583 = ~n96 | n471;
  assign n1584 = ~n96 | n1082;
  assign n1585 = ~n96 | n674;
  assign n1586 = ~n96 | n356;
  assign n1587 = ~n96 | n287;
  assign n1588 = n1587 & n242 & n1586 & n1585 & n1584 & n367 & n1583;
  assign n1589 = ~n163 | n287;
  assign n1590 = ~n163 | n317;
  assign n1591 = ~n96 | n592;
  assign n1592 = ~n163 | n471;
  assign n1593 = ~n163 | n356;
  assign n1594 = ~n163 | n195;
  assign n1595 = n2127 & n2090 & n2124 & n2093 & n2042 & n1897;
  assign n1596 = n1595 & n1594 & n1593 & n1592 & n1591 & n1589 & n1590;
  assign n1597 = n2150 & n2004 & n1992 & n1387 & ~n100 & n192;
  assign n1598 = n1597 & n1496 & n1053 & n1483 & n618 & n646;
  assign n1599 = ~n163 | n979;
  assign n1600 = ~n96 | n1335;
  assign n1601 = ~n163 | n1207;
  assign n1602 = ~n163 | n264;
  assign n1603 = ~n96 | n879;
  assign n1604 = ~n96 | n362;
  assign n1605 = ~n96 | n709;
  assign n1606 = n2046 & n2094 & n1898 & n2092 & n2126 & n2125 & n2047;
  assign n1607 = n1606 & n1605 & n1604 & n1603 & n1602 & n1601 & n1599 & n1600;
  assign n1608 = n172 & n173;
  assign n1609 = n1607 & n1598 & n769 & n760;
  assign n1610 = n2275 & n605 & n1556 & n594 & n830 & n811 & n829 & n1569;
  assign n1611 = n2274 & n2272 & n1629 & n1634 & n1633 & n1635 & n842 & n2152;
  assign n1612 = n706 & n1445 & n463 & n863 & n1359;
  assign n1613 = n1207 | ~n1473;
  assign n1614 = n227 | ~n1473;
  assign n1615 = n879 | ~n1473;
  assign n1616 = ~n98 | n1375;
  assign n1617 = n753 & n1616 & n856;
  assign n1618 = n858 & n1455;
  assign n1619 = n715 | n123 | n818 | n181;
  assign n1620 = n822 | n459;
  assign n1621 = n822 | ~n897;
  assign n1622 = n699 & n1621 & n1620 & n823;
  assign n1623 = n227 | ~n897;
  assign n1624 = n227 | n459;
  assign n1625 = n1624 & n1614 & n1623 & n821 & n711 & n698;
  assign n1626 = ~n97 | n875;
  assign n1627 = n1626 & n1402 & n1350 & n1338 & n213 & ~n844;
  assign n1628 = n898 | n1473 | n818;
  assign n1629 = ~n96 | n392;
  assign n1630 = n1569 & n1629 & n605;
  assign n1631 = n875 | ~n897;
  assign n1632 = n1357 & n1631 & n702 & n876;
  assign n1633 = ~n96 | n822;
  assign n1634 = ~n96 | n567;
  assign n1635 = ~n96 | n1105;
  assign n1636 = n1635 & n1634 & n1633 & n1630;
  assign n1637 = n493 & n494 & n635 & n1607;
  assign n1638 = n1422 & n250 & n1588 & n1596;
  assign n1639 = n666 & n1339 & n1403 & n224 & n665 & n1961;
  assign n1640 = n1639 & n663 & n448 & n207 & n871 & n764 & n874;
  assign n1641 = n701 & n1358 & n1615 & n1366 & n1443;
  assign n1642 = n2027 & n667 & n2152 & n1351 & n846 & n487 & n315 & n624;
  assign n1643 = n1642 & n841 & n843 & n1627 & n727 & n669 & n810 & n1556;
  assign n1644 = n831 & n1598 & n748;
  assign n1645 = ~n136 | n1230;
  assign n1646 = n1237 & ~n481 & ~n1214;
  assign n1647 = n1236 & ~n1214 & n172 & ~n481;
  assign n1648 = n891 & n1625 & n1632;
  assign n1649 = n1247 & n610;
  assign n1650 = n911 | n523;
  assign n1651 = n1105 | n911;
  assign n1652 = n907 | n1375;
  assign n1653 = n911 | n1375;
  assign n1654 = n911 | n567;
  assign n1655 = n907 | n426;
  assign n1656 = n907 | n592;
  assign n1657 = n907 | n685;
  assign n1658 = n907 | n653;
  assign n1659 = n907 | n910;
  assign n1660 = n907 | n1125;
  assign n1661 = n907 | n682;
  assign n1662 = n508 & n536;
  assign n1663 = n1373 & n1125;
  assign n1664 = n330 & n1293;
  assign n1665 = n1664 & n1043;
  assign n1666 = n1138 & n658;
  assign n1667 = ~n278 | n527;
  assign n1668 = ~n278 | n707;
  assign n1669 = ~n278 | n442;
  assign n1670 = n1669 & n1668 & n1667 & n950;
  assign n1671 = ~n278 | n1105;
  assign n1672 = ~n278 | n392;
  assign n1673 = ~n278 | n444;
  assign n1674 = ~n278 | n329;
  assign n1675 = n1401 & n1674 & n1673 & n1671 & n1672;
  assign n1676 = n1097 & n738 & n264 & n540 & n266;
  assign n1677 = n1166 & n316 & n191 & ~n268;
  assign n1678 = n965 & n1677 & n739 & n879 & n361;
  assign n1679 = ~n278 | n1334;
  assign n1680 = ~n278 | n604;
  assign n1681 = ~n278 | n822;
  assign n1682 = ~n278 | n530;
  assign n1683 = n2081 & n1932 & n2156;
  assign n1684 = n1683 & n1682 & n1681 & n1675 & n1054 & n1119 & n1679 & n1680;
  assign n1685 = ~n165 | n393;
  assign n1686 = ~n165 | n444;
  assign n1687 = ~n165 | n566;
  assign n1688 = ~n165 | n567;
  assign n1689 = ~n165 | n1105;
  assign n1690 = ~n165 | n822;
  assign n1691 = ~n165 | n1796;
  assign n1692 = ~n165 | n309;
  assign n1693 = ~n165 | n1157;
  assign n1694 = ~n165 | n529;
  assign n1695 = ~n165 | n1248;
  assign n1696 = ~n165 | n1372;
  assign n1697 = ~n165 | n489;
  assign n1698 = ~n165 | n1155;
  assign n1699 = n1254 | ~n1379;
  assign n1700 = ~n278 | n499;
  assign n1701 = ~n278 | n500;
  assign n1702 = ~n165 | n707;
  assign n1703 = ~n165 | n442;
  assign n1704 = ~n165 | n527;
  assign n1705 = n2174 & n2220 & n1872 & n940 & n2029 & n1963;
  assign n1706 = ~n165 | n265;
  assign n1707 = ~n165 | n526;
  assign n1708 = ~n165 | n984;
  assign n1709 = ~n165 | n1138;
  assign n1710 = ~n165 | n472;
  assign n1711 = ~n165 | n226;
  assign n1712 = ~n165 | n313;
  assign n1713 = n2010 & n2194 & n2101 & n1875 & n1895 & n2054 & n1894;
  assign n1714 = ~n278 | n471;
  assign n1715 = ~n278 | n356;
  assign n1716 = n2292 & (n1259 | ~n1388);
  assign n1717 = ~n165 | n287;
  assign n1718 = ~n278 | n592;
  assign n1719 = ~n278 | n426;
  assign n1720 = n2129 & n1929 & n2053 & n1873;
  assign n1721 = n1720 & n1719 & n1718 & n1717 & n1716 & n1715 & ~n931 & n1714;
  assign n1722 = ~n278 | n688;
  assign n1723 = ~n278 | n774;
  assign n1724 = ~n278 | n1372;
  assign n1725 = ~n278 | n440;
  assign n1726 = n1725 & n1724 & n1723 & n639;
  assign n1727 = ~n278 | n1250;
  assign n1728 = ~n278 | n1375;
  assign n1729 = ~n278 | n1151;
  assign n1730 = n1729 & n1728 & n1727 & n637;
  assign n1731 = n739 & n1160;
  assign n1732 = ~n116 | n2368;
  assign n1733 = ~n116 | n592;
  assign n1734 = ~n116 | n685;
  assign n1735 = ~n116 | n317;
  assign n1736 = ~n116 | n2373;
  assign n1737 = ~n116 | n474;
  assign n1738 = ~n116 | n910;
  assign n1739 = ~n116 | n682;
  assign n1740 = ~n116 | n1335;
  assign n1741 = ~n116 | n1125;
  assign n1742 = ~n116 | n495;
  assign n1743 = ~n167 | n523;
  assign n1744 = ~n167 | n392;
  assign n1745 = ~n404 | n656;
  assign n1746 = ~n404 | n707;
  assign n1747 = ~n404 | n1336;
  assign n1748 = ~n404 | n1293;
  assign n1749 = ~n167 | n1262;
  assign n1750 = ~n167 | n306;
  assign n1751 = ~n167 | n504;
  assign n1752 = ~n167 | n1330;
  assign n1753 = ~n167 | n288;
  assign n1754 = n2070 & n2106 & n1888 & n271;
  assign n1755 = n317 & n1373 & n287;
  assign n1756 = n1755 & n1408 & n1407 & n1380 & n1139 & n525 & ~n450 & n470;
  assign n1757 = ~n404 | n951;
  assign n1758 = ~n404 | n651;
  assign n1759 = ~n167 | n500;
  assign n1760 = ~n167 | n651;
  assign n1761 = ~n167 | n951;
  assign n1762 = ~n167 | n499;
  assign n1763 = n2015 & n1970;
  assign n1764 = n1763 & n1762 & n1761 & n1760 & n1759 & n1758 & n1757 & n1325;
  assign n1765 = ~n167 | n592;
  assign n1766 = ~n167 | n685;
  assign n1767 = ~n167 | n1084;
  assign n1768 = ~n167 | n356;
  assign n1769 = ~n167 | n287;
  assign n1770 = ~n167 | n317;
  assign n1771 = n2095 & n1902 & n2056 & n2002 & n2055 & n1885;
  assign n1772 = n1771 & n1770 & n1769 & n1768 & n1767 & n1765 & n1766;
  assign n1773 = ~n404 | n444;
  assign n1774 = ~n404 | n1105;
  assign n1775 = ~n404 | n1331;
  assign n1776 = n393 | ~n404;
  assign n1777 = ~n404 | n822;
  assign n1778 = n2219 & n1934 & n1966 & n2033 & n2130 & n2181 & n2064 & n1900;
  assign n1779 = n1778 & n1730 & n1013 & n1777 & n1776 & n1775 & n1773 & n1774;
  assign n1780 = ~n404 | n489;
  assign n1781 = n2020 & n1883 & n2202;
  assign n1782 = n2300 & n1967 & n2034 & n1903 & n1886 & n2063 & n2217 & n2131;
  assign n1783 = n1782 & n1781 & n1780 & n1000 & n1397 & n1286 & n611 & n1726;
  assign n1784 = ~n107 | n442;
  assign n1785 = ~n107 | n656;
  assign n1786 = ~n107 | n707;
  assign n1787 = n1786 & n1785 & ~n1045 & n1784;
  assign n1788 = ~n104 | n527;
  assign n1789 = ~n104 | n1261;
  assign n1790 = n1787 & n1788 & n1789;
  assign n1791 = ~n571 | n1155;
  assign n1792 = ~n571 | n2374;
  assign n1793 = ~n571 | n1261;
  assign n1794 = n1793 & n1792 & n1791 & n1044;
  assign n1795 = n440 & n530;
  assign n1796 = n536 & n729;
  assign n1797 = n309 & n336;
  assign n1798 = ~n107 | n1372;
  assign n1799 = ~n104 | n1372;
  assign n1800 = ~n107 | n774;
  assign n1801 = n2019 & n2196 & n1920 & n1945;
  assign n1802 = n1801 & n1800 & n1799 & n1798 & ~n108 & ~n112;
  assign n1803 = n1047 & n1876 & n1472 & n854 & n1316 & n788;
  assign n1804 = n1803 & n1794 & n1790 & n1764 & n974 & n1031;
  assign n1805 = ~n104 | n473;
  assign n1806 = ~n104 | n206;
  assign n1807 = ~n107 | n1028;
  assign n1808 = n1807 & n1805 & n1806;
  assign n1809 = ~n113 | n499;
  assign n1810 = ~n113 | n500;
  assign n1811 = n1343 & (~n294 | (n793 & n1029));
  assign n1812 = n1811 & n1810 & n1809 & ~n1066 & n502 & ~n1065;
  assign n1813 = ~n113 | n1028;
  assign n1814 = ~n113 | n684;
  assign n1815 = ~n113 | n1261;
  assign n1816 = ~n571 | n1027;
  assign n1817 = ~n113 | n1027;
  assign n1818 = ~n113 | n2370;
  assign n1819 = ~n104 | n707;
  assign n1820 = ~n104 | n442;
  assign n1821 = ~n104 | n499;
  assign n1822 = ~n104 | n656;
  assign n1823 = n1822 & n1821 & n1820 & n1819 & ~n106 & ~n1064;
  assign n1824 = ~n104 | n1028;
  assign n1825 = ~n107 | n527;
  assign n1826 = ~n107 | n1261;
  assign n1827 = ~n107 | n592;
  assign n1828 = ~n104 | n287;
  assign n1829 = ~n104 | n317;
  assign n1830 = ~n104 | n471;
  assign n1831 = ~n104 | n356;
  assign n1832 = n2105 & n2066 & n1907;
  assign n1833 = n2305 & n2179 & n2031 & n1947 & n1940 & n1917 & ~n111 & n432;
  assign n1834 = ~n571 | n2210;
  assign n1835 = ~n571 | n1112;
  assign n1836 = ~n113 | n1375;
  assign n1837 = n415 & n256;
  assign n1838 = ~n113 | n822;
  assign n1839 = ~n113 | n1113;
  assign n1840 = n495 & n1125;
  assign n1841 = n291 & ~n930;
  assign n1842 = ~n113 | n2369;
  assign n1843 = ~n113 | n910;
  assign n1844 = ~n113 | n2376;
  assign n1845 = ~n113 | n1125;
  assign n1846 = ~n113 | n495;
  assign n1847 = ~n104 | n362;
  assign n1848 = ~n107 | n1125;
  assign n1849 = ~n104 | n495;
  assign n1850 = ~n104 | n1207;
  assign n1851 = ~n104 | n474;
  assign n1852 = ~n104 | n1125;
  assign n1853 = ~n104 | n709;
  assign n1854 = ~n113 | n2375;
  assign n1855 = n1854 & n1069 & n1071;
  assign n1856 = ~n97 | n1374;
  assign n1857 = ~n97 | n1224;
  assign n1858 = ~n97 | n798;
  assign n1859 = n1858 & n1856 & n1857;
  assign n1860 = ~n96 | n330;
  assign n1861 = n1025 & n1684 & n1022 & n1859;
  assign n1862 = n1861 & n1670 & n1192 & n1810 & n1860 & n1809;
  assign n1863 = ~n571 | n1139;
  assign n1864 = ~n113 | n1138;
  assign n1865 = n2337 & n2082 & n2170 & n2107 & n2146 & n2138;
  assign n1866 = n739 & n749;
  assign n1867 = n684 & n306;
  assign n1868 = n266 & n495;
  assign n1869 = n441 & n658;
  assign n1870 = n284 & n212;
  assign n1871 = ~n98 | n474;
  assign n1872 = ~n165 | n1261;
  assign n1873 = ~n165 | n356;
  assign n1874 = ~n165 | n206;
  assign n1875 = ~n165 | n227;
  assign n1876 = ~n404 | n1261;
  assign n1877 = ~n165 | n1207;
  assign n1878 = n226 | ~n404;
  assign n1879 = n227 | ~n404;
  assign n1880 = n206 | ~n404;
  assign n1881 = n251 | ~n404;
  assign n1882 = ~n404 | n474;
  assign n1883 = ~n404 | n1157;
  assign n1884 = ~n404 | n1207;
  assign n1885 = n356 | ~n404;
  assign n1886 = ~n404 | n1248;
  assign n1887 = ~n107 | n444;
  assign n1888 = ~n167 | n206;
  assign n1889 = ~n104 | n226;
  assign n1890 = n331 | ~n571;
  assign n1891 = ~n163 | n926;
  assign n1892 = n1551 & n1191 & n1511 & n1530 & n1540 & n1891;
  assign n1893 = ~n98 | n879;
  assign n1894 = ~n165 | n875;
  assign n1895 = ~n165 | n284;
  assign n1896 = n1895 & n1503 & n1524 & n1894 & n1667 & n1704;
  assign n1897 = ~n163 | n674;
  assign n1898 = ~n163 | n879;
  assign n1899 = ~n404 | n979;
  assign n1900 = ~n404 | n508;
  assign n1901 = n284 | ~n404;
  assign n1902 = ~n404 | n674;
  assign n1903 = n309 | ~n404;
  assign n1904 = n1903 & n1902 & n1901 & n1774 & n1899 & n1900;
  assign n1905 = ~n167 | n1293;
  assign n1906 = ~n404 | n1262;
  assign n1907 = ~n104 | n674;
  assign n1908 = (~n163 | n191) & (~n167 | n527);
  assign n1909 = n999 & (n327 | (n1295 & n1294));
  assign n1910 = n293 | n875;
  assign n1911 = ~n96 | n191;
  assign n1912 = ~n96 | n527;
  assign n1913 = ~n278 | n926;
  assign n1914 = n191 | ~n278;
  assign n1915 = ~n96 | n979;
  assign n1916 = ~n107 | n1105;
  assign n1917 = ~n107 | n287;
  assign n1918 = ~n167 | n926;
  assign n1919 = ~n167 | n284;
  assign n1920 = ~n107 | n309;
  assign n1921 = ~n107 | n926;
  assign n1922 = ~n107 | n284;
  assign n1923 = (n1649 | n911) & (n292 | n267);
  assign n1924 = n291 & ~n453;
  assign n1925 = n327 & ~n404;
  assign n1926 = (n306 | n1925) & (n266 | ~n344);
  assign n1927 = n190 | ~n278;
  assign n1928 = ~n97 | n316;
  assign n1929 = ~n278 | n317;
  assign n1930 = n1929 & n1633 & n1586;
  assign n1931 = n206 | ~n278;
  assign n1932 = ~n278 | n1157;
  assign n1933 = ~n167 | n251;
  assign n1934 = ~n167 | n822;
  assign n1935 = ~n167 | n216;
  assign n1936 = ~n278 | n316;
  assign n1937 = n216 | ~n278;
  assign n1938 = n997 & n1937 & n1936 & n1935 & n1933 & n1934;
  assign n1939 = ~n167 | n1207;
  assign n1940 = ~n107 | n317;
  assign n1941 = n1938 & n1014 & n1940 & n1939 & n1770 & n1768;
  assign n1942 = ~n113 | n316;
  assign n1943 = n1091 & n1942 & (n316 | ~n353);
  assign n1944 = n1274 & (~n107 | n206);
  assign n1945 = ~n107 | n1157;
  assign n1946 = ~n107 | n822;
  assign n1947 = ~n107 | n356;
  assign n1948 = ~n107 | n216;
  assign n1949 = ~n278 | n1261;
  assign n1950 = n226 | ~n278;
  assign n1951 = ~n96 | n226;
  assign n1952 = n227 | ~n278;
  assign n1953 = ~n97 | n822;
  assign n1954 = ~n96 | n1261;
  assign n1955 = ~n97 | n227;
  assign n1956 = ~n167 | n1261;
  assign n1957 = ~n113 | n1157;
  assign n1958 = ~n113 | n1870;
  assign n1959 = ~n96 | n774;
  assign n1960 = n1959 & n1188;
  assign n1961 = ~n97 | n2370;
  assign n1962 = n1960 & n1961 & n835 & n1492 & n503 & n1466 & n1459 & n858;
  assign n1963 = ~n278 | n331;
  assign n1964 = n1963 & n1723 & n1727;
  assign n1965 = ~n167 | n755;
  assign n1966 = ~n167 | n1250;
  assign n1967 = ~n167 | n774;
  assign n1968 = ~n353 & ~n253 & ~n96 & ~n167;
  assign n1969 = ~n165 | n334;
  assign n1970 = n331 | ~n404;
  assign n1971 = n1386 & n872 & n742 & n832 & n1515 & n1495 & n1969 & n1970;
  assign n1972 = n339 | n341 | n342 | n345 | ~n1854 | ~n1971 | ~n1049 | ~n1835;
  assign n1973 = (n291 | n337) & (~n354 | n1866);
  assign n1974 = (n332 | n1292) & (~n453 | n1731);
  assign n1975 = ~n360 & n1974 & (~n116 | n308);
  assign n1976 = (n310 | ~n571) & (~n107 | n307);
  assign n1977 = n1975 & n1976 & (~n348 | n1310);
  assign n1978 = (n1291 | n674) & (n1925 | n604);
  assign n1979 = (n289 | n327) & (~n351 | n610);
  assign n1980 = (~n113 | n1112) & (~n346 | n687);
  assign n1981 = n1980 & (~n268 | ~n404);
  assign n1982 = (~n253 | n536) & (n330 | ~n930);
  assign n1983 = (~n163 | n190) & (~n167 | n191);
  assign n1984 = n1981 & n1978 & n1979 & n1982 & n1983 & n315 & n328 & n335;
  assign n1985 = n192 & n196 & n199 & n207 & n210 & n1329 & n202;
  assign n1986 = n1985 & n213 & n1325 & n262 & n303 & n1316 & n551 & n277;
  assign n1987 = n334 & n1222;
  assign n1988 = (n481 | n1042) & (~n116 | n1203);
  assign n1989 = (n1042 | n1211) & (~n899 | n1222);
  assign n1990 = n1446 | n459;
  assign n1991 = ~n96 | n430;
  assign n1992 = ~n97 | n430;
  assign n1993 = n1992 & n1559 & n1545 & n1991 & n1581 & n1580 & n1583 & n1584;
  assign n1994 = ~n278 | n1330;
  assign n1995 = ~n278 | n472;
  assign n1996 = ~n278 | n1335;
  assign n1997 = ~n167 | n441;
  assign n1998 = ~n278 | n1337;
  assign n1999 = ~n278 | n430;
  assign n2000 = ~n167 | n1337;
  assign n2001 = ~n167 | n430;
  assign n2002 = ~n167 | n1082;
  assign n2003 = n591 & n644 & n311;
  assign n2004 = ~n98 | ~n450;
  assign n2005 = n2003 & n193 & n1561 & n615 & n189 & n2004 & n661 & n1424;
  assign n2006 = n743 & n1460 & n1463 & n1485;
  assign n2007 = n607 & n603 & n1189 & n791;
  assign n2008 = n2007 & n1421 & n1328 & n600 & n1470 & n596;
  assign n2009 = n1494 & n786 & n779;
  assign n2010 = ~n165 | n1224;
  assign n2011 = ~n98 | n1346;
  assign n2012 = ~n97 | n2373;
  assign n2013 = n2008 & n2009 & n1514 & n623 & n2012 & n2011 & n1698 & n2010;
  assign n2014 = ~n165 | n440;
  assign n2015 = ~n404 | n1155;
  assign n2016 = n535 & n2014 & n2015;
  assign n2017 = ~n120 & (n1292 | (n489 & n1155));
  assign n2018 = n2017 & n1736 & n1285 & n647 & ~n455 & ~n454 & ~n451 & ~n452;
  assign n2019 = ~n104 | n440;
  assign n2020 = ~n404 | n440;
  assign n2021 = (n440 | ~n633) & (n1341 | n1925);
  assign n2022 = (~n349 | n1248) & (~n382 | n1138);
  assign n2023 = (~n294 | n445) & (n539 | n1097);
  assign n2024 = ~n96 | n1348;
  assign n2025 = (~n346 | n1151) & (~n348 | n444);
  assign n2026 = n2025 & (~n98 | n1207);
  assign n2027 = ~n97 | n1138;
  assign n2028 = n1426 & n665 & n2027 & n1427 & n1449 & n1458 & n1491 & n1465;
  assign n2029 = ~n278 | n1155;
  assign n2030 = ~n113 | n1097;
  assign n2031 = ~n107 | n1097;
  assign n2032 = ~n167 | n1341;
  assign n2033 = ~n167 | n1151;
  assign n2034 = ~n167 | n440;
  assign n2035 = ~n278 | n1145;
  assign n2036 = ~n107 & ~n353;
  assign n2037 = n1490 & n1563 & n1481;
  assign n2038 = ~n163 | n1337;
  assign n2039 = ~n163 | n430;
  assign n2040 = n2038 & n2039;
  assign n2041 = ~n163 | n1330;
  assign n2042 = ~n163 | n1082;
  assign n2043 = n2040 & n1528 & n2042 & n1543 & n1538 & n1550 & n2041 & n1508;
  assign n2044 = ~n98 | n709;
  assign n2045 = ~n98 | n1335;
  assign n2046 = ~n163 | n709;
  assign n2047 = ~n163 | n1335;
  assign n2048 = n2047 & n2046 & n1500 & n1523;
  assign n2049 = n2048 & n1629 & n1566 & n1575 & n1576 & n1592;
  assign n2050 = ~n165 | n473;
  assign n2051 = n1702 & n2050 & n1668;
  assign n2052 = ~n165 | n709;
  assign n2053 = ~n165 | n471;
  assign n2054 = ~n165 | n441;
  assign n2055 = ~n404 | n471;
  assign n2056 = ~n404 | n1082;
  assign n2057 = n2055 & n2056;
  assign n2058 = ~n167 | n1336;
  assign n2059 = ~n404 | n441;
  assign n2060 = ~n404 | n1330;
  assign n2061 = n2057 & n2060 & n2059 & n2058 & n1023 & n1740 & n1672 & n1679;
  assign n2062 = ~n404 | n1335;
  assign n2063 = ~n404 | n1334;
  assign n2064 = n392 | ~n404;
  assign n2065 = n2064 & n2062 & n2063;
  assign n2066 = ~n104 | n1082;
  assign n2067 = ~n104 | n472;
  assign n2068 = ~n107 | n393;
  assign n2069 = n2068 & n1853 & n2067 & n1744;
  assign n2070 = ~n167 | n473;
  assign n2071 = (~n107 | n392) & (~n404 | n473);
  assign n2072 = ~n96 & ~n404;
  assign n2073 = (~n295 | n1082) & (n1337 | n2072);
  assign n2074 = (~n381 | n472) & (~n382 | n441);
  assign n2075 = ~n278 | n495;
  assign n2076 = ~n278 | n684;
  assign n2077 = ~n353 | n361;
  assign n2078 = ~n167 | n684;
  assign n2079 = ~n278 | n1333;
  assign n2080 = ~n278 | n361;
  assign n2081 = ~n278 | n566;
  assign n2082 = ~n113 | n566;
  assign n2083 = ~n113 | n489;
  assign n2084 = ~n167 | n1333;
  assign n2085 = n2084 & n1657 & n1655 & n1814 & n2083 & n1759 & n2082 & n1766;
  assign n2086 = (~n107 | n363) & (~n278 | n1138);
  assign n2087 = ~n107 | n1333;
  assign n2088 = ~n163 | n684;
  assign n2089 = ~n163 | n1333;
  assign n2090 = ~n163 | n685;
  assign n2091 = n2090 & n1541 & n2089 & n724 & n1512 & n1549 & n2088;
  assign n2092 = ~n163 | n495;
  assign n2093 = ~n163 | n426;
  assign n2094 = ~n163 | n362;
  assign n2095 = ~n404 | n426;
  assign n2096 = ~n167 | n656;
  assign n2097 = n1742 & n1722 & n1734 & n1775 & n2095 & n2096;
  assign n2098 = ~n165 | n447;
  assign n2099 = ~n165 | n500;
  assign n2100 = ~n165 | n362;
  assign n2101 = ~n165 | n845;
  assign n2102 = ~n107 | n1331;
  assign n2103 = n2102 & n1745 & n1780 & n1107 & n1847 & n1849;
  assign n2104 = n911 | n489;
  assign n2105 = ~n104 | n426;
  assign n2106 = ~n167 | n447;
  assign n2107 = ~n571 | n1138;
  assign n2108 = ~n162 & (~n930 | (n656 & n685));
  assign n2109 = (n323 | n495) & (~n346 | n684);
  assign n2110 = ~n383 & (n447 | (~n113 & ~n278));
  assign n2111 = (~n404 | n1408) & (n1333 | n2072);
  assign n2112 = n485 & n1005 & (~n294 | n475);
  assign n2113 = ~n476 & (n327 | (n430 & n729));
  assign n2114 = (~n349 | n529) & (n291 | n1404);
  assign n2115 = n1291 | n1082;
  assign n2116 = (~n96 | n495) & (~n359 | n489);
  assign n2117 = n2116 & (n481 | n459);
  assign n2118 = n226 | ~n897;
  assign n2119 = ~n98 | n682;
  assign n2120 = ~n98 | n1125;
  assign n2121 = n734 & n2120 & n2119 & n1480 & n1562 & n771 & n1489;
  assign n2122 = ~n163 | n504;
  assign n2123 = ~n163 | n1028;
  assign n2124 = ~n163 | n592;
  assign n2125 = ~n163 | n682;
  assign n2126 = ~n163 | n1125;
  assign n2127 = ~n163 | n653;
  assign n2128 = n957 & n1486 & n1696 & n2127 & n2126 & n1522 & n2125;
  assign n2129 = ~n165 | n592;
  assign n2130 = ~n404 | n567;
  assign n2131 = ~n404 | n1372;
  assign n2132 = ~n404 | n499;
  assign n2133 = n911 | n1372;
  assign n2134 = n2133 & n1821 & n1799 & n1739 & n2132 & n2130 & n2131;
  assign n2135 = n911 | n528;
  assign n2136 = ~n104 | n567;
  assign n2137 = ~n104 | n984;
  assign n2138 = ~n571 | n984;
  assign n2139 = (~n381 | n682) & (n910 | n1841);
  assign n2140 = ~n278 | n1027;
  assign n2141 = n2140 & ~n101 & ~n111;
  assign n2142 = ~n113 | n1084;
  assign n2143 = ~n278 | n2376;
  assign n2144 = ~n107 | n2371;
  assign n2145 = ~n113 | n1796;
  assign n2146 = ~n113 | n1139;
  assign n2147 = n1006 & n2146 & (~n167 | n362);
  assign n2148 = ~n97 | n1125;
  assign n2149 = ~n96 | n499;
  assign n2150 = ~n97 | n1176;
  assign n2151 = n1493 & n1558 & n2150 & n1553 & n2148 & n2149;
  assign n2152 = ~n96 | n984;
  assign n2153 = ~n278 | n1028;
  assign n2154 = ~n96 | n1373;
  assign n2155 = n2151 & n1634 & n1591 & n2154 & n2153 & n2152 & n1700;
  assign n2156 = ~n278 | n567;
  assign n2157 = ~n278 | n1125;
  assign n2158 = ~n278 | n1373;
  assign n2159 = n2158 & n2157 & n1724 & n1718 & n2156 & n945;
  assign n2160 = ~n167 | n1028;
  assign n2161 = ~n353 | n1373;
  assign n2162 = ~n353 | n1176;
  assign n2163 = ~n278 | n1176;
  assign n2164 = ~n167 | n1372;
  assign n2165 = ~n167 | n1125;
  assign n2166 = ~n107 | n567;
  assign n2167 = ~n113 | n1372;
  assign n2168 = ~n107 | n984;
  assign n2169 = ~n107 | n1373;
  assign n2170 = ~n113 | n567;
  assign n2171 = n667 & n666 & n1425;
  assign n2172 = n783 & n1520 & n1498;
  assign n2173 = n1205 | ~n1388;
  assign n2174 = ~n278 | n951;
  assign n2175 = ~n167 | n530;
  assign n2176 = ~n278 | n521;
  assign n2177 = ~n167 | n522;
  assign n2178 = n2177 & n2175 & n2176;
  assign n2179 = ~n107 | n540;
  assign n2180 = ~n113 | n540;
  assign n2181 = ~n167 | n1375;
  assign n2182 = ~n928 | n1663;
  assign n2183 = (~n278 | n653) & (n675 | n926);
  assign n2184 = n533 & n879 & n504;
  assign n2185 = n1200 | ~n1379;
  assign n2186 = n620 & n194;
  assign n2187 = n2186 & n645 & n312 & n616 & n214 & n1423 & n203 & n662;
  assign n2188 = n1856 & n1535 & n1462 & n741;
  assign n2189 = n1616 & n1469 & n1488;
  assign n2190 = n1190 & n792 & n787 & n776 & n842 & n622 & n1287 & n1653;
  assign n2191 = n2190 & n2189 & n595 & n599 & n1327 & n625 & n606 & n602;
  assign n2192 = ~n98 | n522;
  assign n2193 = ~n165 | n530;
  assign n2194 = ~n165 | n1374;
  assign n2195 = n1738 & n2193 & n2194;
  assign n2196 = ~n104 | n530;
  assign n2197 = n2196 & n1324 & ~n117 & n609;
  assign n2198 = n1757 & (~n354 | (n191 & n1373));
  assign n2199 = ~n542 & (~n453 | (n526 & n1374));
  assign n2200 = (~n97 | n520) & (n680 | n910);
  assign n2201 = (n327 | n524) & (~n294 | n531);
  assign n2202 = ~n404 | n530;
  assign n2203 = (~n165 | n525) & (~n340 | n951);
  assign n2204 = (n309 | ~n348) & (~n359 | n528);
  assign n2205 = n1863 & (~n930 | (n1293 & n1378));
  assign n2206 = n2205 & (~n359 | (n521 & n1176));
  assign n2207 = ~n582 & (n1292 | (n1294 & n1404));
  assign n2208 = ~n583 & (~n571 | (n536 & n1084));
  assign n2209 = (n285 | n875) & (~n104 | n1295);
  assign n2210 = n508 & n467;
  assign n2211 = (n288 | ~n346) & (n251 | ~n340);
  assign n2212 = (~n97 | n216) & (~n165 | n508);
  assign n2213 = n297 & n2212 & n380 & n325;
  assign n2214 = n490 & n492 & n496;
  assign n2215 = n1533 & n1447;
  assign n2216 = ~n96 | n1026;
  assign n2217 = ~n167 | n777;
  assign n2218 = ~n167 | n793;
  assign n2219 = ~n167 | n654;
  assign n2220 = ~n278 | n651;
  assign n2221 = (~n107 | n632) & (n1417 | n1968);
  assign n2222 = ~n107 | n2372;
  assign n2223 = ~n107 | n651;
  assign n2224 = ~n107 | n1666;
  assign n2225 = n2224 & n2223 & n2222 & n2221 & n1760 & n1070 & ~n110 & ~n634;
  assign n2226 = (n1259 | ~n1388) & (~n253 | n793);
  assign n2227 = n491 & (~n404 | (n682 & n1407));
  assign n2228 = ~n163 | n629;
  assign n2229 = n2228 & n1699 & n1384 & n1326 & n1278 & n870 & ~n100 & n840;
  assign n2230 = ~n104 | n1416;
  assign n2231 = ~n104 | n629;
  assign n2232 = n2231 & n2230 & n1758 & n1323 & n1289 & n1284 & ~n106 & n1118;
  assign n2233 = (~n321 | n686) & (~n344 | n689);
  assign n2234 = ~n690 & (~n404 | (n687 & n793));
  assign n2235 = ~n691 & (~n163 | (n651 & n1311));
  assign n2236 = ~n692 & (n597 | (~n167 & ~n930));
  assign n2237 = ~n693 & (n468 | n1309) & n2236;
  assign n2238 = ~n344 & ~n353;
  assign n2239 = (n304 | ~n346) & (n1333 | n2238);
  assign n2240 = n2237 & n2239 & (~n354 | n1429);
  assign n2241 = n2240 & n2235 & n2234 & n2233 & n2232 & n2229 & ~n169 & n1858;
  assign n2242 = (n681 | n777) & (~n338 | n1417);
  assign n2243 = (~n294 | n659) & (~n348 | n660);
  assign n2244 = (~n268 | ~n381) & (n327 | n655);
  assign n2245 = (~n253 | n330) & (~n453 | n798);
  assign n2246 = (~n113 | n313) & (n291 | n447);
  assign n2247 = (~n97 | n362) & (~n98 | n610);
  assign n2248 = (~n104 | n265) & (n738 | n911);
  assign n2249 = n248 & (n941 | ~n1379);
  assign n2250 = n2242 & n2243 & n2244 & n2245 & n2246 & n2247 & n2249 & n2248;
  assign n2251 = n391 & n277 & n683 & n550 & n672 & n1433 & n1438 & n643;
  assign n2252 = n2251 & n594 & n598 & n601 & n1440 & n614 & n608 & n605;
  assign n2253 = (~n107 | n1405) & (~n167 | n1406);
  assign n2254 = (~n404 | n519) & (n710 | n1309);
  assign n2255 = n2254 & (n357 | n471);
  assign n2256 = ~n321 & ~n346;
  assign n2257 = (n2256 | n910) & (n2238 | n1337);
  assign n2258 = (~n294 | n708) & (~n571 | n1086);
  assign n2259 = (~n97 | n429) & (~n321 | n1405);
  assign n2260 = n2259 & (n327 | n1347);
  assign n2261 = n2260 & n2257 & n2258 & n2255 & n863 & n446 & n1351 & n1350;
  assign n2262 = (~n344 | n1334) & (~n348 | n707);
  assign n2263 = n1040 & n2262 & (~n343 | n521);
  assign n2264 = (~n96 | n1176) & (~n165 | n536);
  assign n2265 = n2264 & n2263 & (n481 | n1234);
  assign n2266 = n2265 & n697 & n1445 & n706 & n303 & n412 & n614 & n549;
  assign n2267 = n1236 & n172 & ~n1233;
  assign n2268 = n2039 & n1857 & n1856;
  assign n2269 = n1272 & n233 & n1911;
  assign n2270 = n486 & ~n800 & (~n163 | n799);
  assign n2271 = (~n97 | n763) & (~n98 | n330);
  assign n2272 = n1421 & n218 & n827;
  assign n2273 = n196 & (~n97 | n195);
  assign n2274 = n2273 & n814 & ~n813 & ~n812 & n496 & n492 & n428 & n490;
  assign n2275 = n626 & n624;
  assign n2276 = ~n1233 & n1237;
  assign n2277 = ~n1612 | n181 | n820 | n2276 | n1646 | ~n1858;
  assign n2278 = n826 & (n459 | (n481 & n474));
  assign n2279 = n565 & n217 & n881 & n806 & n808 & n807;
  assign n2280 = n2279 & n2216 & n1955 & n1928 & ~n878 & ~n877 & n422 & n503;
  assign n2281 = n854 & n862 & n866 & n1644 & n1643 & n838;
  assign n2282 = n2281 & n1641 & n868 & n1640 & n1636 & n1632 & n1637 & n1638;
  assign n2283 = n1251 & ~n122 & ~n136;
  assign n2284 = (~n899 | ~n900) & (~n1608 | n2283);
  assign n2285 = n1648 & ~n132 & n884;
  assign n2286 = ~n1237 | n2283;
  assign n2287 = n2286 & (n459 | (n474 & ~n819));
  assign n2288 = n731 & n728 & n2012 & n2011 & n920 & n1858 & n922 & n1455;
  assign n2289 = n506 & n1430;
  assign n2290 = n2099 & n2076 & n2153;
  assign n2291 = n2140 & (~n930 | (n755 & n1418));
  assign n2292 = (~n165 | n426) & (~n278 | n287);
  assign n2293 = n2185 & n2173 & n1952;
  assign n2294 = n2293 & n2158 & n1969 & n2193 & n2014 & n2035 & n2176 & n1950;
  assign n2295 = n2163 & n243 & n2080;
  assign n2296 = (~n165 | n971) & (~n278 | n966);
  assign n2297 = n749 & n1161;
  assign n2298 = n1420 & (~n930 | n2297);
  assign n2299 = n1876 & n2160 & n2078 & n2032 & n2177 & n2218;
  assign n2300 = n2175 & n2164 & n1439;
  assign n2301 = n2084 & n2001 & n1918;
  assign n2302 = n2301 & n2000 & n1935 & n1118 & ~n1039 & ~n1037 & ~n168 & n995;
  assign n2303 = n150 & n228 & (~n167 | n362);
  assign n2304 = n2303 & n1764 & n1036 & n1783 & n1011 & n1779 & n1020 & n1772;
  assign n2305 = (~n104 | n1087) & (~n107 | n1077);
  assign n2306 = n1640 & n1195 & n811 & n1808 & n1036 & n963;
  assign n2307 = n688 & n1380;
  assign n2308 = n742 & n1453 & n1959 & n1419 & n1932 & n1682 & n2014 & n2193;
  assign n2309 = n2256 | n969;
  assign n2310 = ~n1099 & (~n404 | (n287 & n1087));
  assign n2311 = ~n107 | n1046;
  assign n2312 = n2310 & n2311 & n2223;
  assign n2313 = (n292 | n1098) & (n1349 | n1097);
  assign n2314 = (~n104 | ~n109) & (~n354 | n739);
  assign n2315 = (~n165 | n263) & (~n571 | n1136);
  assign n2316 = (n317 | ~n346) & (n305 | ~n453);
  assign n2317 = (~n98 | n774) & (n195 | n1292);
  assign n2318 = n2312 & n2313 & n2314 & n2315 & n2316 & n2317 & n669 & n541;
  assign n2319 = n1454 & n1433 & n785 & n746 & n841 & n831 & n1638 & n140;
  assign n2320 = n993 & n1721 & n1096 & n1772 & n1168 & n1094 & n1076 & n1059;
  assign n2321 = (~n294 | n654) & (~n929 | n1141);
  assign n2322 = (~n165 | n1331) & (~n404 | n566);
  assign n2323 = n2321 & n2322 & n1496 & n1516 & n1636 & n1526;
  assign n2324 = n244 & n1478 & n1479 & n673 & n842 & n1915;
  assign n2325 = ~n1128 & (~n340 | (n921 & n1335));
  assign n2326 = ~n1129 & (~n571 | (n1207 & n1840));
  assign n2327 = n2326 & (n1152 | (~n116 & n1841));
  assign n2328 = (~n346 | n1840) & (~n928 | n1126);
  assign n2329 = (n362 | ~n381) & (n266 | n539);
  assign n2330 = (n291 | n1250) & (n292 | n264);
  assign n2331 = n2329 & n2330 & (n1292 | n879);
  assign n2332 = n2331 & n2327 & n2328 & n2324 & n2325 & n2082 & n2170 & n2222;
  assign n2333 = n510 & n1274 & (~n404 | n709);
  assign n2334 = n2333 & n1411 & n745 & n760 & n1618 & n1518 & n1505 & n753;
  assign n2335 = n938 & n1637 & n141;
  assign n2336 = n2335 & n1020 & n992 & n1170 & n1183 & n1124 & n1804 & n1076;
  assign n2337 = ~n113 | n1869;
  assign n2338 = n2149 & n1451 & n1460 & n957 & n2099 & n1912;
  assign n2339 = n1431 & (~n571 | n1142);
  assign n2340 = (~n404 | n1140) & (n313 | n1924);
  assign n2341 = (~n321 | n1156) & (n651 | n1349);
  assign n2342 = n2341 & (~n349 | n1374);
  assign n2343 = n2340 & n2342 & (n1662 | n509);
  assign n2344 = (~n382 | n798) & (n323 | n951);
  assign n2345 = n2344 & (~n294 | n1224);
  assign n2346 = n1282 & (n292 | n334);
  assign n2347 = n2343 & n2345 & n2346 & n2338 & n2339 & n1825 & n2145 & n2132;
  assign n2348 = n517 & n418 & n335 & n1483 & n560 & n1438;
  assign n2349 = n2348 & n1643 & n801 & n1532 & n780 & n1521;
  assign n2350 = n987 & n949 & n975;
  assign n2351 = n2350 & n1081 & n1011 & n1135 & n1182 & n1862 & n1059 & n1124;
  assign n2352 = n2311 & n1517 & n946 & ~n114 & ~n108 & ~n112;
  assign n2353 = ~n113 | n1143;
  assign n2354 = n2353 & n2352 & n2337 & n1839 & ~n118 & n506;
  assign n2355 = (~n97 | n1154) & (~n107 | n1153);
  assign n2356 = n2355 & (~n113 | n1150);
  assign n2357 = (~n167 | n1146) & (~n278 | n1148);
  assign n2358 = n2357 & (~n96 | n1145);
  assign n2359 = n2354 & n2356 & n2358 & n1414 & n678 & n424 & n372 & n262;
  assign n2360 = n735 & n697 & n643 & n794 & n732 & n772;
  assign n2361 = n2360 & n849 & n841 & n843 & n833 & n1627;
  assign n2362 = n1630 & n874 & n871;
  assign n2363 = n2362 & n1032 & n1004 & n1862 & n1855 & n1103 & n1787 & n1051;
  assign n2364 = n1389 & n1317 & n1948;
  assign n2365 = (~n107 | n1167) & (n1164 | n1292);
  assign n2366 = n2083 & n1314 & n2167 & n627 & n1890 & n1048;
  assign n2367 = n2353 & (~n294 | (n1149 & n1506));
  assign n2368 = n471 & n426 & n356;
  assign n2369 = n1207 & n921;
  assign n2370 = n206 & n762;
  assign n2371 = n845 & n875 & n441;
  assign n2372 = n682 & n266 & n495;
  assign n2373 = n1207 & n470;
  assign n2374 = n1293 & n469;
  assign n2375 = n527 & n209;
  assign n2376 = n879 & n470;
  assign n2377 = n894 | n126;
  assign n2378 = n906 | n126;
  assign n2379 = n480 | n126;
  assign n2380 = n590 | n126;
  assign n2381 = n1259 & n1211 & ~i_12_ & n216;
endmodule


