// Benchmark "top" written by ABC on Tue Mar  5 10:05:48 2019

module tseng ( clock, 
    tin_pv10_4_4_, tin_pv11_4_4_, tin_pv6_7_7_, tin_pv2_0_0_,
    tin_pv10_3_3_, tin_pv1_2_2_, tin_pv11_3_3_, tin_pv4_3_3_,
    tin_pv10_2_2_, tin_pv11_2_2_, tin_pv6_0_0_, tin_pv2_1_1_,
    tin_pv10_1_1_, tin_pv1_3_3_, preset_0_0_, tin_pv11_1_1_, tin_pv4_4_4_,
    tin_pready_0_0_, tin_pv10_0_0_, tin_pv11_0_0_, tin_pv6_1_1_,
    tin_pv2_2_2_, tin_pv1_4_4_, tin_pv4_5_5_, tin_pv6_2_2_, tin_pv2_3_3_,
    tin_pv1_5_5_, tin_pv4_6_6_, tin_pv6_3_3_, tin_pv2_4_4_, tin_pv1_6_6_,
    tin_pv4_7_7_, tin_pv6_4_4_, tin_pv2_5_5_, tin_pv1_7_7_,
    tin_pv4_0_0_, tin_pv6_5_5_, tin_pv2_6_6_, tin_pv10_7_7_, tin_pv1_0_0_,
    tin_pv11_7_7_, tin_pv4_1_1_, tin_pv10_6_6_, tin_pv11_6_6_,
    tin_pv6_6_6_, tin_pv2_7_7_, preset, tin_pv10_5_5_, tin_pv1_1_1_,
    tin_pv11_5_5_, tin_pv4_2_2_,
    pv14_2_2_, pv12_3_3_, pv10_4_4_, pv7_5_5_, pv3_6_6_, pv15_2_2_,
    pv13_3_3_, pv11_4_4_, pv6_7_7_, pv2_0_0_, pv14_1_1_, pv12_2_2_,
    pv10_3_3_, pv9_0_0_, pv5_1_1_, pv1_2_2_, pv15_1_1_, pv13_2_2_,
    pv11_3_3_, pv8_2_2_, pv4_3_3_, pv14_0_0_, pv12_1_1_, pv10_2_2_,
    pv7_6_6_, pv3_7_7_, pv15_0_0_, pv13_1_1_, pv11_2_2_, pv6_0_0_,
    pv2_1_1_, pv12_0_0_, pv10_1_1_, pv9_1_1_, pv5_2_2_, pv1_3_3_,
    pv13_0_0_, pv11_1_1_, pv8_3_3_, pv4_4_4_, pready_0_0_, pv10_0_0_,
    pv7_7_7_, pv3_0_0_, pv11_0_0_, pv6_1_1_, pv2_2_2_, pv9_2_2_, pv5_3_3_,
    pv1_4_4_, pv8_4_4_, pv4_5_5_, pv7_0_0_, pv3_1_1_, pv6_2_2_, pv2_3_3_,
    pv9_3_3_, pv5_4_4_, pv1_5_5_, pv8_5_5_, pv4_6_6_, pv7_1_1_, pv3_2_2_,
    pv6_3_3_, pv2_4_4_, pv9_4_4_, pv5_5_5_, pv1_6_6_, pv8_6_6_, pv4_7_7_,
    pv7_2_2_, pv3_3_3_, pv6_4_4_, pv2_5_5_, pv14_7_7_, pv9_5_5_, pv5_6_6_,
    pv1_7_7_, pv15_7_7_, pv8_7_7_, pv4_0_0_, pv14_6_6_, pv12_7_7_,
    pv7_3_3_, pv3_4_4_, pv15_6_6_, pv13_7_7_, pv6_5_5_, pv2_6_6_, pdn,
    pv14_5_5_, pv12_6_6_, pv10_7_7_, pv9_6_6_, pv5_7_7_, pv1_0_0_,
    pv15_5_5_, pv13_6_6_, pv11_7_7_, pv8_0_0_, pv4_1_1_, pv14_4_4_,
    pv12_5_5_, pv10_6_6_, pv7_4_4_, pv3_5_5_, pv15_4_4_, pv13_5_5_,
    pv11_6_6_, pv6_6_6_, pv2_7_7_, pv14_3_3_, pv12_4_4_, pv10_5_5_,
    pv9_7_7_, pv5_0_0_, pv1_1_1_, pv15_3_3_, pv13_4_4_, pv11_5_5_,
    pv8_1_1_, pv4_2_2_  );
  input  tin_pv10_4_4_, tin_pv11_4_4_, tin_pv6_7_7_, tin_pv2_0_0_,
    tin_pv10_3_3_, tin_pv1_2_2_, tin_pv11_3_3_, tin_pv4_3_3_,
    tin_pv10_2_2_, tin_pv11_2_2_, tin_pv6_0_0_, tin_pv2_1_1_,
    tin_pv10_1_1_, tin_pv1_3_3_, preset_0_0_, tin_pv11_1_1_, tin_pv4_4_4_,
    tin_pready_0_0_, tin_pv10_0_0_, tin_pv11_0_0_, tin_pv6_1_1_,
    tin_pv2_2_2_, tin_pv1_4_4_, tin_pv4_5_5_, tin_pv6_2_2_, tin_pv2_3_3_,
    tin_pv1_5_5_, tin_pv4_6_6_, tin_pv6_3_3_, tin_pv2_4_4_, tin_pv1_6_6_,
    clock, tin_pv4_7_7_, tin_pv6_4_4_, tin_pv2_5_5_, tin_pv1_7_7_,
    tin_pv4_0_0_, tin_pv6_5_5_, tin_pv2_6_6_, tin_pv10_7_7_, tin_pv1_0_0_,
    tin_pv11_7_7_, tin_pv4_1_1_, tin_pv10_6_6_, tin_pv11_6_6_,
    tin_pv6_6_6_, tin_pv2_7_7_, preset, tin_pv10_5_5_, tin_pv1_1_1_,
    tin_pv11_5_5_, tin_pv4_2_2_;
  output pv14_2_2_, pv12_3_3_, pv10_4_4_, pv7_5_5_, pv3_6_6_, pv15_2_2_,
    pv13_3_3_, pv11_4_4_, pv6_7_7_, pv2_0_0_, pv14_1_1_, pv12_2_2_,
    pv10_3_3_, pv9_0_0_, pv5_1_1_, pv1_2_2_, pv15_1_1_, pv13_2_2_,
    pv11_3_3_, pv8_2_2_, pv4_3_3_, pv14_0_0_, pv12_1_1_, pv10_2_2_,
    pv7_6_6_, pv3_7_7_, pv15_0_0_, pv13_1_1_, pv11_2_2_, pv6_0_0_,
    pv2_1_1_, pv12_0_0_, pv10_1_1_, pv9_1_1_, pv5_2_2_, pv1_3_3_,
    pv13_0_0_, pv11_1_1_, pv8_3_3_, pv4_4_4_, pready_0_0_, pv10_0_0_,
    pv7_7_7_, pv3_0_0_, pv11_0_0_, pv6_1_1_, pv2_2_2_, pv9_2_2_, pv5_3_3_,
    pv1_4_4_, pv8_4_4_, pv4_5_5_, pv7_0_0_, pv3_1_1_, pv6_2_2_, pv2_3_3_,
    pv9_3_3_, pv5_4_4_, pv1_5_5_, pv8_5_5_, pv4_6_6_, pv7_1_1_, pv3_2_2_,
    pv6_3_3_, pv2_4_4_, pv9_4_4_, pv5_5_5_, pv1_6_6_, pv8_6_6_, pv4_7_7_,
    pv7_2_2_, pv3_3_3_, pv6_4_4_, pv2_5_5_, pv14_7_7_, pv9_5_5_, pv5_6_6_,
    pv1_7_7_, pv15_7_7_, pv8_7_7_, pv4_0_0_, pv14_6_6_, pv12_7_7_,
    pv7_3_3_, pv3_4_4_, pv15_6_6_, pv13_7_7_, pv6_5_5_, pv2_6_6_, pdn,
    pv14_5_5_, pv12_6_6_, pv10_7_7_, pv9_6_6_, pv5_7_7_, pv1_0_0_,
    pv15_5_5_, pv13_6_6_, pv11_7_7_, pv8_0_0_, pv4_1_1_, pv14_4_4_,
    pv12_5_5_, pv10_6_6_, pv7_4_4_, pv3_5_5_, pv15_4_4_, pv13_5_5_,
    pv11_6_6_, pv6_6_6_, pv2_7_7_, pv14_3_3_, pv12_4_4_, pv10_5_5_,
    pv9_7_7_, pv5_0_0_, pv1_1_1_, pv15_3_3_, pv13_4_4_, pv11_5_5_,
    pv8_1_1_, pv4_2_2_;
  reg n_n4142, n_n3936, n_n3574, n_n3008, n_n3726, n_n3604, n_n3144,
    n_n3782, n_n3067, n_n4258, n_n3225, n_n3180, n_n3274, n_n3475, n_n3687,
    n_n3381, n_n3098, n_n4108, n_n3497, n_n3793, n_n4316, n_n4349, n_n3029,
    n_n3619, n_n3264, n_n3780, ndn3_4, n_n4114, n_n3146, n_n3511, n_n3152,
    n_n3833, n_n4282, n_n3305, n_n4392, n_n4224, n_n3198, n_n3204, n_n3024,
    n_n4139, ndn3_15, n_n3133, n_n4074, n_n3270, n_n3858, n_n3456, n_n3521,
    n_n3081, n_n4381, n_n3670, n_n4211, n_n3493, n_n3495, n_n3916, n_n3195,
    n_n3525, n_n3729, n_n3876, ndn3_5, n_n3549, n_n3489, n_n3764, n_n3281,
    n_n3707, n_n3517, n_n4160, n_n4222, n_n3012, n_n4071, n_n3372, n_n3344,
    n_n3688, n_n3079, n_n3313, n_n3411, n_n3231, n_n3396, n_n3432, n_n3606,
    n_n3733, n_n3556, n_n4040, n_n3120, n_n3221, n_n3173, n_n3851, n_n3113,
    n_n3242, n_n3118, n_n3376, n_n4089, n_n3044, n_n3627, n_n3035, n_n3111,
    n_n3321, n_n3443, n_n3215, ndn3_10, n_n4172, nlc1_2, n_n3590, n_n4110,
    nlc3_3, n_n3576, n_n4129, n_n4189, n_n4286, n_n4383, pdn, n_n3567,
    n_n3892, n_n3075, n_n3354, n_n3465, ndn3_6, n_n3617, n_n4162, n_n3207,
    n_n4120, n_n3065, n_n4005, n_n3266, n_n4337, n_n3600, n_n3415, n_n4243,
    n_n3872, n_n3648, n_n3358, n_n3350, ndn3_7, n_n3116, n_n3583, n_n3906,
    n_n4131, n_n3316, n_n3061, n_n3048, n_n3886, n_n3919, n_n3128, n_n3995,
    n_n4213, n_n3761, ndn3_8, n_n3252, n_n4366, n_n3328, n_n3988, n_n3348,
    n_n3544, n_n3101, n_n4279, n_n3896, n_n3736, n_n4251, n_n3650, n_n3307,
    n_n4294, n_n4334, n_n3955, n_n4164, n_n3155, n_n3749, n_n4233, n_n4347,
    n_n3826, n_n3360, n_n3458, n_n3093, n_n3157, n_n3506, n_n3161, n_n3319,
    n_n3429, n_n3971, n_n3449, n_n4270, n_n4288, n_n3183, n_n3130, nlak4_2,
    n_n4047, n_n3978, n_n3239, n_n4145, n_n3890, n_n4003, n_n3091, n_n3985,
    n_n3326, n_n4052, nsr4_2, n_n4099, n_n4375, n_n4067, n_n4290, n_n3898,
    n_n4122, n_n3774, n_n3014, n_n4241, n_n3952, n_n3237, n_n3968, n_n3922,
    n_n3551, n_n3379, n_n4275, n_n3570, n_n3854, n_n4057, n_n3451, n_n4037,
    n_n3408, n_n4229, n_n4201, n_n3339, n_n4362, n_n3483, n_n3557, n_n4185,
    n_n3069, n_n3643, n_n3404, n_n3057, n_n3020, n_n3828, n_n3631, n_n3138,
    nsr1_2, n_n4065, n_n3679, n_n3287, n_n4351, n_n4059, n_n3436, nen3_10,
    n_n3461, n_n4012, n_n3051, n_n3073, n_n3777, n_n3709, n_n3946, n_n3085,
    n_n3259, n_n3504, n_n4045, n_n3954, n_n3136, n_n4372, n_n4236, n_n3040,
    n_n3874, n_n3999, n_n3223, ndn1_34, n_n3743, n_n3657, n_n3213, n_n3095,
    n_n3663, n_n3724, n_n3038, n_n3370, n_n3624, n_n3578, n_n3713, n_n3089,
    n_n3211, n_n3367, n_n3434, n_n3126, n_n4192, n_n4136, n_n3053, n_n3938,
    n_n3769, n_n4390, nsr3_17, n_n3903, n_n3658, nrq3_11, n_n3818, n_n3533,
    n_n3463, n_n3175, n_n3055, n_n3202, n_n3385, n_n4077, n_n3142, n_n3901,
    n_n3934, n_n3823, n_n3722, n_n4309, n_n4159, n_n4330, n_n3836, n_n3470,
    n_n3331, n_n3883, n_n4299, n_n4157, ndn3_9, n_n3208, n_n3190, n_n4029,
    n_n3042, nsr3_14, n_n4151, n_n3188, n_n4303, n_n3250, n_n3170, n_n3758,
    n_n3910, n_n3108, n_n3150, n_n4320, n_n4360, n_n4247, n_n4199, n_n3966,
    n_n3766, n_n4021, n_n4062, n_n3514, n_n3572, n_n4166, n_n3976, n_n3394,
    n_n4095, n_n3863, n_n3720, ngfdn_3, n_n3756, n_n3667, n_n3342, n_n3529,
    n_n4209, n_n4324, n_n3337, n_n4227, n_n4153, n_n3831, n_n3233, n_n4263,
    n_n3413, n_n4182, n_n3841, n_n3441, n_n4026, n_n4342, n_n4102, n_n3277,
    n_n4180, n_n3878, n_n3931, n_n3845, n_n3865, n_n3486, n_n4056, n_n3674,
    n_n3959, n_n3608, n_n4080, n_n4018, n_n4354, n_n3797, n_n3739, n_n3646,
    n_n3099, n_n3537, n_n3806, n_n3087, n_n4105, n_n3262, n_n4125, n_n3814,
    n_n4093, nsr3_3;
  wire n1835, n1836, n1837, n1838_1, n1839, n1840, n1841, n1842, n1843_1,
    n1844, n1845, n1846, n1847, n1848_1, n1849, n1850, n1851, n1852,
    n1853_1, n1854, n1855, n1856, n1857, n1858_1, n1859, n1860, n1861,
    n1862, n1863_1, n1864, n1865, n1866, n1867, n1868_1, n1869, n1870,
    n1871, n1872, n1873_1, n1874, n1875, n1876, n1877, n1878_1, n1879,
    n1880, n1881, n1882, n1883_1, n1884, n1885, n1886, n1887, n1888_1,
    n1889, n1890, n1891, n1892, n1893_1, n1894, n1895, n1896, n1897,
    n1898_1, n1899, n1900, n1901, n1902, n1903_1, n1904, n1905, n1906,
    n1907, n1908_1, n1909, n1910, n1911, n1912, n1913_1, n1914, n1915,
    n1916, n1917, n1918_1, n1919, n1920, n1921, n1922, n1923_1, n1924,
    n1925, n1926, n1927, n1928_1, n1929, n1930, n1931, n1932, n1933_1,
    n1934, n1935, n1936, n1937, n1938_1, n1939, n1940, n1941, n1942,
    n1943_1, n1944, n1945, n1946, n1947, n1948_1, n1949, n1950, n1951,
    n1952, n1953_1, n1954, n1955, n1956, n1957, n1958_1, n1959, n1960,
    n1961, n1962, n1963_1, n1964, n1965, n1966, n1967, n1968_1, n1969,
    n1970, n1971, n1972, n1973_1, n1974, n1975, n1976, n1977, n1978_1,
    n1979, n1980, n1981, n1982, n1983_1, n1984, n1985, n1986, n1987,
    n1988_1, n1989, n1990, n1991, n1992, n1993_1, n1994, n1995, n1996,
    n1997, n1998_1, n1999, n2000, n2001, n2002, n2003_1, n2004, n2005,
    n2006, n2007, n2008_1, n2009, n2010, n2011, n2012, n2013_1, n2014,
    n2015, n2016, n2017, n2018_1, n2019, n2020, n2021, n2022, n2023_1,
    n2024, n2025, n2026, n2027, n2028_1, n2029, n2030, n2031, n2032,
    n2033_1, n2034, n2035, n2036, n2037, n2038_1, n2039, n2040, n2041,
    n2042, n2043_1, n2044, n2045, n2046, n2047, n2048_1, n2049, n2050,
    n2051, n2052, n2053_1, n2054, n2055, n2056, n2057, n2058_1, n2059,
    n2060, n2061, n2062, n2063_1, n2064, n2065, n2066, n2067, n2068_1,
    n2069, n2070, n2071, n2072, n2073_1, n2074, n2075, n2076, n2077,
    n2078_1, n2079, n2080, n2081, n2082, n2083_1, n2084, n2085, n2086,
    n2087, n2088_1, n2089, n2090, n2091, n2092, n2093_1, n2094, n2095,
    n2096, n2097, n2098_1, n2099, n2100, n2101, n2102, n2103_1, n2104,
    n2105, n2106, n2107, n2108_1, n2109, n2110, n2111, n2112, n2113_1,
    n2114, n2115, n2116, n2117, n2118_1, n2119, n2120, n2121, n2122,
    n2123_1, n2124, n2125, n2126, n2127, n2128_1, n2129, n2130, n2131,
    n2132, n2133_1, n2134, n2135, n2136, n2137, n2138_1, n2139, n2140,
    n2141, n2142, n2143_1, n2144, n2145, n2146, n2147, n2148_1, n2149,
    n2150, n2151, n2152, n2153_1, n2154, n2155, n2156, n2157, n2158_1,
    n2159, n2160, n2161, n2162, n2163_1, n2164, n2165, n2166, n2167,
    n2168_1, n2169, n2170, n2171, n2172, n2173_1, n2174, n2175, n2176,
    n2177, n2178_1, n2179, n2180, n2181, n2182, n2183_1, n2184, n2185,
    n2186, n2187, n2188_1, n2189, n2190, n2191, n2192, n2193_1, n2194,
    n2195, n2196, n2197, n2198_1, n2199, n2200, n2201, n2202, n2203_1,
    n2204, n2205, n2206, n2207, n2208_1, n2209, n2210, n2211, n2212,
    n2213_1, n2214, n2215, n2216, n2217, n2218_1, n2219, n2220, n2221,
    n2222, n2223_1, n2224, n2225, n2226, n2227, n2228_1, n2229, n2230,
    n2231, n2232, n2233_1, n2234, n2235, n2236, n2237, n2238_1, n2239,
    n2240, n2241, n2242, n2243_1, n2244, n2245, n2246, n2247, n2248_1,
    n2249, n2250, n2251, n2252, n2253_1, n2254, n2255, n2256, n2257,
    n2258_1, n2259, n2260, n2261, n2262, n2263_1, n2264, n2265, n2266,
    n2267, n2268_1, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
    n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
    n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
    n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
    n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
    n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
    n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
    n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
    n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
    n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
    n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n349, n354,
    n359, n364, n369, n374, n379, n384, n389, n394, n399, n404, n409, n414,
    n419, n424, n429, n434, n439, n444, n449, n454, n459, n464, n469, n474,
    n479, n484, n489, n494, n499, n504, n509, n514, n519, n524, n529, n534,
    n539, n544, n549, n554, n559, n564, n569, n574, n579, n584, n589, n594,
    n599, n604, n609, n614, n619, n624, n629, n634, n639, n644, n649, n654,
    n659, n664, n669, n674, n679, n684, n689, n694, n699, n704, n709, n714,
    n719, n724, n729, n734, n739, n744, n749, n754, n759, n764, n769, n774,
    n779, n784, n789, n794, n799, n804, n809, n814, n819, n824, n829, n834,
    n839, n844, n849, n854, n859, n864, n869, n874, n879, n884, n889, n894,
    n898, n903, n908, n913, n918, n923, n928, n933, n938, n943, n948, n953,
    n958, n963, n968, n973, n978, n983, n988, n993, n998, n1003, n1008,
    n1013, n1018, n1023, n1028, n1033, n1038, n1043, n1048, n1053, n1058,
    n1063, n1068, n1073, n1078, n1083, n1088, n1093, n1098, n1103, n1108,
    n1113, n1118, n1123, n1128, n1133, n1138, n1143, n1148, n1153, n1158,
    n1163, n1168, n1173, n1178, n1183, n1188, n1193, n1198, n1203, n1208,
    n1213, n1218, n1223, n1228, n1233, n1238, n1243, n1248, n1253, n1258,
    n1263, n1268, n1273, n1278, n1283, n1288, n1293, n1298, n1303, n1308,
    n1313, n1318, n1323, n1328, n1333, n1338, n1343, n1348, n1353, n1358,
    n1363, n1368, n1373, n1378, n1383, n1388, n1393, n1398, n1403, n1408,
    n1413, n1418, n1423, n1428, n1433, n1438, n1443, n1448, n1453, n1458,
    n1463, n1468, n1473, n1478, n1483, n1488, n1493, n1498, n1503, n1508,
    n1513, n1518, n1523, n1528, n1533, n1538, n1543, n1548, n1553, n1558,
    n1563, n1568, n1573, n1578, n1583, n1588, n1593, n1598, n1603, n1608,
    n1613, n1618, n1623, n1628, n1633, n1638, n1643, n1648, n1653, n1658,
    n1663, n1668, n1673, n1678, n1683, n1688, n1693, n1698, n1703, n1708,
    n1713, n1718, n1723, n1728, n1733, n1738, n1743, n1748, n1753, n1758,
    n1763, n1768, n1773, n1778, n1783, n1788, n1793, n1798, n1803, n1808,
    n1813, n1818, n1823, n1828, n1833, n1838, n1843, n1848, n1853, n1858,
    n1863, n1868, n1873, n1878, n1883, n1888, n1893, n1898, n1903, n1908,
    n1913, n1918, n1923, n1928, n1933, n1938, n1943, n1948, n1953, n1958,
    n1963, n1968, n1973, n1978, n1983, n1988, n1993, n1998, n2003, n2008,
    n2013, n2018, n2023, n2028, n2033, n2038, n2043, n2048, n2053, n2058,
    n2063, n2068, n2073, n2078, n2083, n2088, n2093, n2098, n2103, n2108,
    n2113, n2118, n2123, n2128, n2133, n2138, n2143, n2148, n2153, n2158,
    n2163, n2168, n2173, n2178, n2183, n2188, n2193, n2198, n2203, n2208,
    n2213, n2218, n2223, n2228, n2233, n2238, n2243, n2248, n2253, n2258,
    n2263, n2268;
  assign pv14_2_2_ = n_n3358 & n_n4153;
  assign pv12_3_3_ = n_n3631 & n_n3367;
  assign pv10_4_4_ = n_n3042 ? n_n4136 : tin_pv10_4_4_;
  assign pv7_5_5_ = n_n3130 & n_n3679;
  assign pv3_6_6_ = n_n3252 & n_n3057;
  assign pv15_2_2_ = n_n3113 & n_n4037;
  assign pv13_3_3_ = n_n3600 & n_n3404;
  assign pv11_4_4_ = n_n4120 ? n_n3966 : tin_pv11_4_4_;
  assign pv6_7_7_ = n_n4164 ? n_n3370 : tin_pv6_7_7_;
  assign pv2_0_0_ = n_n3211 ? n_n3910 : tin_pv2_0_0_;
  assign pv14_1_1_ = n_n3012 & n_n3038;
  assign pv12_2_2_ = n_n3067 & n_n3576;
  assign pv10_3_3_ = n_n4129 ? n_n3213 : tin_pv10_3_3_;
  assign pv9_0_0_ = n_n3128 & n_n3890;
  assign pv5_1_1_ = n_n3443 & n_n3287;
  assign pv1_2_2_ = n_n3470 ? n_n3537 : tin_pv1_2_2_;
  assign pv15_1_1_ = n_n3606 & n_n3108;
  assign pv13_2_2_ = n_n3379 & n_n3463;
  assign pv11_3_3_ = n_n3432 ? n_n3583 : tin_pv11_3_3_;
  assign pv8_2_2_ = n_n3456 & n_n3055;
  assign pv4_3_3_ = n_n3489 ? n_n4309 : tin_pv4_3_3_;
  assign pv14_0_0_ = n_n3761 & n_n3903;
  assign pv12_1_1_ = n_n3264 & n_n4390;
  assign pv10_2_2_ = n_n3065 ? n_n3549 : tin_pv10_2_2_;
  assign pv7_6_6_ = n_n3670 & n_n3617;
  assign pv3_7_7_ = n_n3590 & n_n4102;
  assign pv15_0_0_ = n_n4003 & n_n3188;
  assign pv13_1_1_ = n_n3221 & n_n3150;
  assign pv11_2_2_ = n_n3152 ? n_n3823 : tin_pv11_2_2_;
  assign pv6_0_0_ = n_n3029 ? n_n3506 : tin_pv6_0_0_;
  assign pv2_1_1_ = n_n3999 ? n_n3646 : tin_pv2_1_1_;
  assign pv12_0_0_ = n_n3098 & n_n3339;
  assign pv10_1_1_ = n_n3872 ? n_n3270 : tin_pv10_1_1_;
  assign pv9_1_1_ = n_n3024 & n_n3044;
  assign pv5_2_2_ = n_n4286 & n_n3350;
  assign pv1_3_3_ = n_n3441 ? n_n4180 : tin_pv1_3_3_;
  assign pv13_0_0_ = n_n3061 & n_n3434;
  assign pv11_1_1_ = n_n4185 ? n_n4142 : tin_pv11_1_1_;
  assign pv8_3_3_ = n_n3146 & n_n3091;
  assign pv4_4_4_ = n_n4110 ? n_n3627 : tin_pv4_4_4_;
  assign pready_0_0_ = n_n4108 ? n_n3354 : tin_pready_0_0_;
  assign pv10_0_0_ = n_n4282 ? n_n4209 : tin_pv10_0_0_;
  assign pv7_7_7_ = n_n3136 & n_n4077;
  assign pv3_0_0_ = n_n3173 & n_n3828;
  assign pv11_0_0_ = n_n3233 ? n_n3514 : tin_pv11_0_0_;
  assign pv6_1_1_ = n_n3144 ? n_n3952 : tin_pv6_1_1_;
  assign pv2_2_2_ = n_n4354 ? n_n3202 : tin_pv2_2_2_;
  assign pv9_2_2_ = n_n3736 & n_n3157;
  assign pv5_3_3_ = n_n3321 & n_n4236;
  assign pv1_4_4_ = n_n3863 ? n_n3806 : tin_pv1_4_4_;
  assign pv8_4_4_ = n_n3344 & n_n3095;
  assign pv4_5_5_ = n_n3087 ? n_n3733 : tin_pv4_5_5_;
  assign pv7_0_0_ = n_n3161 & n_n3069;
  assign pv3_1_1_ = n_n3048 & n_n3461;
  assign pv6_2_2_ = n_n3307 ? n_n3138 : tin_pv6_2_2_;
  assign pv2_3_3_ = n_n3874 ? n_n3465 : tin_pv2_3_3_;
  assign pv9_3_3_ = n_n3906 & n_n3749;
  assign pv5_4_4_ = n_n3793 & n_n4213;
  assign pv1_5_5_ = n_n3101 ? n_n3313 : tin_pv1_5_5_;
  assign pv8_5_5_ = n_n3116 & n_n3331;
  assign pv4_6_6_ = n_n3774 ? n_n3413 : tin_pv4_6_6_;
  assign pv7_1_1_ = n_n3415 & n_n3971;
  assign pv3_2_2_ = n_n3190 & n_n3739;
  assign pv6_3_3_ = n_n3204 ? n_n3486 : tin_pv6_3_3_;
  assign pv2_4_4_ = n_n3643 ? n_n3133 : tin_pv2_4_4_;
  assign pv9_4_4_ = n_n3687 & n_n3650;
  assign pv5_5_5_ = n_n3266 & n_n3408;
  assign pv1_6_6_ = n_n4018 ? n_n3118 : tin_pv1_6_6_;
  assign pv8_6_6_ = n_n3180 & n_n3223;
  assign pv4_7_7_ = n_n4114 ? n_n4166 : tin_pv4_7_7_;
  assign pv7_2_2_ = n_n3497 & n_n4105;
  assign pv3_3_3_ = n_n3274 & n_n4342;
  assign pv6_4_4_ = n_n3093 ? n_n4065 : tin_pv6_4_4_;
  assign pv2_5_5_ = n_n4059 ? n_n3780 : tin_pv2_5_5_;
  assign pv14_7_7_ = n_n3449 & n_n4241;
  assign pv9_5_5_ = n_n3985 & n_n4290;
  assign pv5_6_6_ = n_n3567 & n_n3237;
  assign pv1_7_7_ = n_n3544 ? n_n4199 : tin_pv1_7_7_;
  assign pv15_7_7_ = n_n3079 & n_n3648;
  assign pv8_7_7_ = n_n3525 & n_n3529;
  assign pv4_0_0_ = n_n3826 ? n_n3517 : tin_pv4_0_0_;
  assign pv14_6_6_ = n_n3713 & n_n3262;
  assign pv12_7_7_ = n_n3764 & n_n3720;
  assign pv7_3_3_ = n_n3411 & n_n4303;
  assign pv3_4_4_ = n_n3729 & n_n4162;
  assign pv15_6_6_ = n_n4375 & n_n3020;
  assign pv13_7_7_ = n_n3372 & n_n3394;
  assign pv6_5_5_ = n_n3348 ? n_n4189 : tin_pv6_5_5_;
  assign pv2_6_6_ = n_n3120 ? n_n3385 : tin_pv2_6_6_;
  assign pv14_5_5_ = n_n3008 & n_n3663;
  assign pv12_6_6_ = n_n3782 & n_n3896;
  assign pv10_7_7_ = n_n3521 ? n_n3225 : tin_pv10_7_7_;
  assign pv9_6_6_ = n_n4243 & n_n3239;
  assign pv5_7_7_ = n_n3111 & n_n4005;
  assign pv1_0_0_ = n_n3551 ? n_n4192 : tin_pv1_0_0_;
  assign pv15_5_5_ = n_n3277 & n_n3674;
  assign pv13_6_6_ = n_n3155 & n_n3797;
  assign pv11_7_7_ = n_n3360 ? n_n3376 : tin_pv11_7_7_;
  assign pv8_0_0_ = n_n3014 & n_n4320;
  assign pv4_1_1_ = n_n4089 ? n_n3722 : tin_pv4_1_1_;
  assign pv14_4_4_ = n_n3326 & n_n3089;
  assign pv12_5_5_ = n_n3619 & n_n3337;
  assign pv10_6_6_ = n_n3570 ? n_n3342 : tin_pv10_6_6_;
  assign pv7_4_4_ = n_n3073 & n_n3053;
  assign pv3_5_5_ = n_n3436 & n_n3142;
  assign pv15_4_4_ = n_n3305 & n_n3667;
  assign pv13_5_5_ = n_n4139 & n_n3777;
  assign pv11_6_6_ = n_n3504 ? n_n4279 : tin_pv11_6_6_;
  assign pv6_6_6_ = n_n3836 ? n_n3429 : tin_pv6_6_6_;
  assign pv2_7_7_ = n_n4131 ? n_n3126 : tin_pv2_7_7_;
  assign pv14_3_3_ = n_n3396 & n_n3316;
  assign pv12_4_4_ = n_n3231 & n_n3175;
  assign pv10_5_5_ = n_n3381 ? n_n4247 : tin_pv10_5_5_;
  assign pv9_7_7_ = n_n3319 & n_n3040;
  assign pv5_0_0_ = n_n3195 & n_n3572;
  assign pv1_1_1_ = n_n3215 ? n_n3183 : tin_pv1_1_1_;
  assign pv15_3_3_ = n_n4172 & n_n3051;
  assign pv13_4_4_ = n_n3075 & n_n3758;
  assign pv11_5_5_ = n_n3081 ? n_n3207 : tin_pv11_5_5_;
  assign pv8_1_1_ = n_n3938 & n_n3883;
  assign pv4_2_2_ = n_n4347 ? n_n4372 : tin_pv4_2_2_;
  assign n349 = n2312 | (n_n3724 & ~n1922 & n2315);
  assign n354 = (pv11_1_1_ & n1835) | n2311;
  assign n359 = n2309 | n2307 | n2308;
  assign n364 = n2306 | (n_n3035 & n_n4157 & n1839);
  assign n369 = n2305 | n2303 | n2304;
  assign n374 = ~preset & n1837;
  assign n379 = ~preset & (n_n3144 | (~pdn & n1870));
  assign n384 = ~preset & (n_n3782 | (~pdn & n1870));
  assign n389 = ~preset & (n_n3067 | (~pdn & n1870));
  assign n394 = (pv10_3_3_ & n1838_1) | n2302;
  assign n399 = (n_n4360 & n1839) | n2301;
  assign n404 = ~preset & (n_n3180 | (~pdn & n1870));
  assign n409 = ~preset & (n_n3274 | (~pdn & n1870));
  assign n414 = n_n3475 ? (n1841 | (n1840 & n1990)) : (n1840 & ~n1990);
  assign n419 = (n_n3458 & n1839) | n2300;
  assign n424 = ~preset & (n_n3381 | (~pdn & n1870));
  assign n429 = n2299 | (n_n3688 & n_n3624 & n1839);
  assign n434 = ~preset & n1842;
  assign n439 = n2298 | (n_n3901 & n1839 & n1890);
  assign n444 = n2297 | (n1839 & (~n_n3916 ^ n1930));
  assign n449 = (n1844 & n1845) | n2282;
  assign n454 = (pv6_0_0_ & n1846) | n2281;
  assign n459 = ~preset & (n_n3029 | (~pdn & n1870));
  assign n464 = ~preset & (n_n3619 | (~pdn & n1870));
  assign n469 = ~preset & (n_n3264 | (~pdn & n1870));
  assign n474 = n2280 | (n1839 & (n_n4288 | n2319));
  assign n479 = n1847 & ~preset & ~ngfdn_3;
  assign n484 = ~preset & (n_n4114 | (~pdn & n1870));
  assign n489 = ~preset & (n_n3146 | (~pdn & n1870));
  assign n494 = (pv1_5_5_ & n1848_1) | n2279;
  assign n499 = ~preset & (n_n3152 | (~pdn & n1870));
  assign n504 = preset | (n_n3833 & n1850) | (~n1849 & ~n1850);
  assign n509 = ~preset & (n_n4282 | (~pdn & n1870));
  assign n514 = ~preset & (n_n3305 | (~pdn & n1870));
  assign n519 = n2278 | (n1851 & (~n1905 ^ n1978_1));
  assign n524 = (pv4_5_5_ & n1852) | n2277;
  assign n529 = ~preset & (~n1983_1 | ~n1984) & n2331;
  assign n534 = ~preset & (n_n3204 | (~pdn & n1870));
  assign n539 = ~preset & (n_n3024 | (~pdn & n1870));
  assign n544 = ~preset & (n_n4139 | (~pdn & n1870));
  assign n549 = ~ngfdn_3 & ~preset & ndn3_15;
  assign n554 = n2274 | (n1839 & (n_n3458 | n2332));
  assign n559 = n2262 | (n2038 & (~n1909 ^ n1974));
  assign n564 = (n_n3743 & n1839) | n2261;
  assign n569 = (pv1_2_2_ & n1848_1) | n2260;
  assign n574 = ~preset & (n_n3456 | (~pdn & n1870));
  assign n579 = ~preset & (n_n3521 | (~pdn & n1870));
  assign n584 = ~preset & (n_n3081 | (~pdn & n1870));
  assign n589 = n2257 | (n1853_1 & (n2258_1 | n2336));
  assign n594 = n2256 | (n_n3475 & n1839 & n1890);
  assign n599 = (pv11_2_2_ & n1835) | n2255;
  assign n604 = n_n4045 & n2337 & (n1890 | ~n2335);
  assign n609 = (n1844 & n1851) | n2254;
  assign n614 = n2253_1 | (n1845 & (~n1909 ^ n1974));
  assign n619 = ~preset & (n_n3195 | (~pdn & n1870));
  assign n624 = (n_n3242 & n1839) | n2252;
  assign n629 = (n_n3916 & n1839) | n2251;
  assign n634 = (pv10_4_4_ & n1838_1) | n2250;
  assign n639 = ~preset & ~ngfdn_3 & (ndn3_4 | ndn3_5);
  assign n644 = (n_n3946 & n1839) | n2249;
  assign n649 = ~preset & (n_n3489 | (~pdn & n1870));
  assign n654 = n2248_1 | (n_n3242 & n_n3170 & n1839);
  assign n659 = (pv2_3_3_ & n1854) | n2247;
  assign n664 = n2246 | preset | n1855;
  assign n669 = (n_n4159 & n1839) | n2245;
  assign n674 = (pv4_1_1_ & n1852) | n2244;
  assign n679 = n2243_1 | (n1845 & (~n1905 ^ n1978_1));
  assign n684 = n2242 | (n_n3936 & n_n3099 & n1839);
  assign n689 = (pv6_5_5_ & n1846) | n2241;
  assign n694 = ~preset & (n_n3372 | (~pdn & n1870));
  assign n699 = (n_n4074 & n1839) | n2240;
  assign n704 = n2239 | (n2038 & (n1972 ^ n1973_1));
  assign n709 = n2238_1 | (n1839 & (n_n4233 | n2338));
  assign n714 = n2237 | (n_n3035 & n_n4157 & n1839);
  assign n719 = ~preset & (n_n3411 | (~pdn & n1870));
  assign n724 = n2236 | (n_n4074 & n_n3578 & n1839);
  assign n729 = ~preset & (n_n3396 | (~pdn & n1870));
  assign n734 = ~preset & (n_n3432 | (~pdn & n1870));
  assign n739 = ~preset & (n_n3606 | (~pdn & n1870));
  assign n744 = (n_n4224 & n1839) | n2235;
  assign n749 = (pv11_6_6_ & n1835) | n2234;
  assign n754 = n2233_1 | n2231 | n2232;
  assign n759 = ~preset & (n_n3120 | (~pdn & n1870));
  assign n764 = (n_n4222 & n1839) | n2230;
  assign n769 = (n_n3976 & n1839) | n2229;
  assign n774 = ~preset & (n1987 ? n_n3851 : n1953_1);
  assign n779 = n2228_1 | (n1839 & (n_n3495 | n2341));
  assign n784 = n2212 | n2213_1;
  assign n789 = n2211 | (n_n3556 & n_n4122 & n1839);
  assign n794 = n2210 | (n_n3483 & ~n1922 & n2315);
  assign n799 = ~preset & (n_n4089 | (~pdn & n1870));
  assign n804 = (n_n4392 & n1839) | n2209;
  assign n809 = (n_n4330 & n1839) | n2208_1;
  assign n814 = (pv11_5_5_ & n1835) | n2207;
  assign n819 = n2206 | (n1839 & (~n_n3841 ^ n1901));
  assign n824 = ~preset & (n_n3321 | (~pdn & n1870));
  assign n829 = ~preset & (n_n3443 | (~pdn & n1870));
  assign n834 = ~preset & (n_n3215 | (~pdn & n1870));
  assign n839 = ~preset & ~ngfdn_3 & (ndn3_10 | nen3_10);
  assign n844 = n2205 | (n1839 & (n_n4351 | n2346));
  assign n849 = n1859 & ~preset & ~pdn;
  assign n854 = ~preset & (n_n3590 | (~pdn & n1870));
  assign n859 = ~preset & (n_n4110 | (~pdn & n1870));
  assign n864 = ~n1858_1 & (nlc3_3 | (n1956 & n2347));
  assign n869 = n2204 | (n_n4211 & n_n3657 & n1839);
  assign n874 = ~preset & (n_n4129 | (~pdn & n1870));
  assign n879 = (n_n4071 & n1839) | n2203_1;
  assign n884 = (n1839 & n1860) | n2202;
  assign n889 = (pv4_2_2_ & n1852) | n2201;
  assign n894 = n1870 & ~preset & ~pdn;
  assign n898 = ~preset & (n_n3567 | (~pdn & n1870));
  assign n903 = (pv6_6_6_ & n1846) | n2200;
  assign n908 = ~preset & (n_n3075 | (~pdn & n1870));
  assign n913 = n2199 | (~preset & ~pdn & n1870);
  assign n918 = n2198_1 | (n1839 & (n_n4351 | n2346));
  assign n923 = ~preset & ~ngfdn_3 & (ndn3_5 | ndn3_6);
  assign n928 = ~preset & (n_n3617 | (~pdn & n1870));
  assign n933 = ~preset & (n_n4162 | (~pdn & n1870));
  assign n938 = n2197 | (n_n4012 & ~n1922 & n2315);
  assign n943 = ~preset & (n_n4120 | (~pdn & n1870));
  assign n948 = ~preset & (n_n3065 | (~pdn & n1870));
  assign n953 = ~preset & (n_n4005 | (~pdn & n1870));
  assign n958 = ~preset & (n_n3266 | (~pdn & n1870));
  assign n963 = (pv6_7_7_ & n1846) | n2196;
  assign n968 = ~preset & (n_n3600 | (~pdn & n1870));
  assign n973 = ~preset & (n_n3415 | (~pdn & n1870));
  assign n978 = (n_n4095 & n1839) | n2195;
  assign n983 = ~preset & (n_n3872 | (~pdn & n1870));
  assign n988 = ~preset & (n_n3648 | (~pdn & n1870));
  assign n993 = n2194 | (n_n4211 & n_n3657 & n1839);
  assign n998 = ~preset & (n_n3350 | (~pdn & n1870));
  assign n1003 = ~preset & ~ngfdn_3 & (ndn3_6 | ndn3_7);
  assign n1008 = ~preset & (n_n3116 | (~pdn & n1870));
  assign n1013 = n2193_1 | (n_n3766 & ~n1922 & n2315);
  assign n1018 = (n_n4351 & n1839) | n2192;
  assign n1023 = ~preset & (n_n4131 | (~pdn & n1870));
  assign n1028 = n2191 | (n_n3085 & n_n3250 & n1839);
  assign n1033 = (n_n3976 & n1839) | n2190;
  assign n1038 = (n_n4222 & n1839) | n2189;
  assign n1043 = (pv1_4_4_ & n1848_1) | n2188_1;
  assign n1048 = (pv1_6_6_ & n1848_1) | n2187;
  assign n1053 = (n_n3608 & n1839) | n2186;
  assign n1058 = n2185 | n2183_1 | n2184;
  assign n1063 = ~preset & (n_n4213 | (~pdn & n1870));
  assign n1068 = n2182 | (n_n3688 & n_n3624 & n1839);
  assign n1073 = ~preset & ~ngfdn_3 & (ndn3_7 | ndn3_8);
  assign n1078 = ~preset & (n_n3252 | (~pdn & n1870));
  assign n1083 = n_n4366 ? (n1841 | (n1840 & n1991)) : (n1840 & ~n1991);
  assign n1088 = (pv2_1_1_ & n1854) | n2181;
  assign n1093 = n2180 | n2178_1 | n2179;
  assign n1098 = ~preset & (n_n3348 | (~pdn & n1870));
  assign n1103 = ~preset & (n_n3544 | (~pdn & n1870));
  assign n1108 = ~preset & (n_n3101 | (~pdn & n1870));
  assign n1113 = n2177 | (n_n4334 & ~n1922 & n2315);
  assign n1118 = n2176 | (n_n3556 & n_n4122 & n1839);
  assign n1123 = (n_n3495 & n1839) | n2175;
  assign n1128 = (pv4_6_6_ & n1852) | n2174;
  assign n1133 = ~preset & (n_n3650 | (~pdn & n1870));
  assign n1138 = ~preset & (n_n3307 | (~pdn & n1870));
  assign n1143 = (pv1_3_3_ & n1848_1) | n2173_1;
  assign n1148 = n_n4334 ? (n1872 | n2171) : n1862;
  assign n1153 = n2169 | (n1853_1 & (n2170 | n2350));
  assign n1158 = ~preset & (n_n4164 | (~pdn & n1870));
  assign n1163 = (n_n4145 & n1839) | n2168_1;
  assign n1168 = ~preset & (n_n3749 | (~pdn & n1870));
  assign n1173 = n2166 | n2167;
  assign n1178 = ~preset & (n_n4347 | (~pdn & n1870));
  assign n1183 = ~preset & (n_n3826 | (~pdn & n1870));
  assign n1188 = ~preset & (n_n3360 | (~pdn & n1870));
  assign n1193 = n2165 | (n1851 & (~n1909 ^ n1974));
  assign n1198 = ~preset & (n_n3093 | (~pdn & n1870));
  assign n1203 = ~preset & (n_n3157 | (~pdn & n1870));
  assign n1208 = (n_n4349 & n1839) | n2164;
  assign n1213 = ~preset & (n_n3161 | (~pdn & n1870));
  assign n1218 = (n_n4233 & n1839) | n2163_1;
  assign n1223 = (n_n3892 & n1839) | n2162;
  assign n1228 = n2161 | (n_n4125 & n1839 & n1890);
  assign n1233 = n2160 | (n_n3242 & n_n3170 & n1839);
  assign n1238 = (pv4_7_7_ & n1852) | n2159;
  assign n1243 = (n1851 & n1863_1) | n2158_1;
  assign n1248 = n2157 | (n_n3936 & n_n3099 & n1839);
  assign n1253 = ~preset & (n_n3130 | (~pdn & n1870));
  assign n1258 = ~n1864 & ~preset & nsr4_2;
  assign n1263 = n2156 | (~preset & n_n4047 & ~n1886);
  assign n1268 = (pv2_2_2_ & n1854) | n2155;
  assign n1273 = ~preset & (n_n3239 | (~pdn & n1870));
  assign n1278 = n2153_1 | n2154;
  assign n1283 = ~preset & (n_n3890 | (~pdn & n1870));
  assign n1288 = n2152 | (n1839 & (n_n3608 | n2324));
  assign n1293 = (n_n3085 & n1839) | n2151;
  assign n1298 = (n_n4288 & n1839) | n2150;
  assign n1303 = ~preset & (n_n3326 | (~pdn & n1870));
  assign n1308 = n2147 | (n1853_1 & (n2149 | n2352));
  assign n1313 = pdn | preset | (nsr4_2 & n1864);
  assign n1318 = n2145 | (n1853_1 & (n2146 | n2353));
  assign n1323 = ~preset & (n_n4375 | (~pdn & n1870));
  assign n1328 = n1865 & ~preset & ~n1855;
  assign n1333 = ~preset & (n_n4290 | (~pdn & n1870));
  assign n1338 = (n1845 & n1863_1) | n2144;
  assign n1343 = n2142 | n2143_1;
  assign n1348 = ~preset & (n_n3774 | (~pdn & n1870));
  assign n1353 = ~preset & (n_n3014 | (~pdn & n1870));
  assign n1358 = ~preset & (n_n4241 | (~pdn & n1870));
  assign n1363 = (n_n4201 & n1839) | n2141;
  assign n1368 = n2140 | (n1839 & (~n_n4145 ^ n1895));
  assign n1373 = (pv6_2_2_ & n1846) | n2139;
  assign n1378 = (pv6_4_4_ & n1846) | n2138_1;
  assign n1383 = ~preset & (n_n3551 | (~pdn & n1870));
  assign n1388 = ~preset & (n_n3379 | (~pdn & n1870));
  assign n1393 = (n_n4275 & n1868_1) | n2133_1;
  assign n1398 = ~preset & (n_n3570 | (~pdn & n1870));
  assign n1403 = (pv2_5_5_ & n1854) | n2132;
  assign n1408 = n2131 | n2358;
  assign n1413 = (pv2_7_7_ & n1854) | n2130;
  assign n1418 = ~preset & (n_n4037 | (~pdn & n1870));
  assign n1423 = n2129 | (n1839 & (~n_n3898 ^ n1896));
  assign n1428 = n2127 | n2128_1;
  assign n1433 = (pv6_1_1_ & n1846) | n2126;
  assign n1438 = ~preset & (n_n3339 | (~pdn & n1870));
  assign n1443 = (pv10_5_5_ & n1838_1) | n2125;
  assign n1448 = n2123_1 | (n_n4334 & ~n_n3483 & n1862);
  assign n1453 = ~preset & n2357 & (n_n4099 ^ n1967);
  assign n1458 = ~preset & (n_n4185 | (~pdn & n1870));
  assign n1463 = n2122 | (n_n3934 & n1839 & n1890);
  assign n1468 = ~preset & (n_n3643 | (~pdn & n1870));
  assign n1473 = (n_n4229 & n1839) | n2121;
  assign n1478 = (n_n4145 & n1839) | n2120;
  assign n1483 = n2119 | (n1839 & (n_n4095 | n2345));
  assign n1488 = ~preset & (n_n3828 | (~pdn & n1870));
  assign n1493 = n2118_1 | (n_n3085 & n_n3250 & n1839);
  assign n1498 = (n_n3968 & n1839) | n2117;
  assign n1503 = pdn | preset | (~ngfdn_3 & ~n1870);
  assign n1508 = (n_n3922 & n1839) | n2116;
  assign n1513 = n2115 | (n_n4366 & n1839 & n1890);
  assign n1518 = (n1839 & n1871) | n2114;
  assign n1523 = n2112 | n2113_1;
  assign n1528 = ~preset & (n_n4059 | (~pdn & n1870));
  assign n1533 = (n_n3898 & n1839) | n2111;
  assign n1538 = ~preset & ~ngfdn_3 & (nen3_10 | ndn3_9);
  assign n1543 = ~preset & (n_n3461 | (~pdn & n1870));
  assign n1548 = (n_n4012 & n1872) | n2110;
  assign n1553 = ~preset & (n_n3051 | (~pdn & n1870));
  assign n1558 = n2109 | (n_n4047 & n1839 & n1890);
  assign n1563 = (n_n3898 & n1839) | n2108_1;
  assign n1568 = n2359 & (n2107 | (n1878_1 & n2317));
  assign n1573 = (pv10_2_2_ & n1838_1) | n2106;
  assign n1578 = n2104 | n2105;
  assign n1583 = (pv1_7_7_ & n1848_1) | n2103_1;
  assign n1588 = ~preset & (n_n3504 | (~pdn & n1870));
  assign n1593 = n2362 | (n_n4045 & (n2102 | n2361));
  assign n1598 = ~n2100 & (~n1853_1 | (~n2101 & ~n2363));
  assign n1603 = n2099 | (n_n4324 & n1839 & n1890);
  assign n1608 = (n_n4383 & n1839) | n2098_1;
  assign n1613 = n2097 | (n1839 & (~n_n4229 ^ n1902));
  assign n1618 = ~preset & (n_n3040 | (~pdn & n1870));
  assign n1623 = ~preset & (n_n3874 | (~pdn & n1870));
  assign n1628 = ~preset & (n_n3999 | (~pdn & n1870));
  assign n1633 = (n_n4122 & n1839) | n2096;
  assign n1638 = ndn1_34 & ~preset & ~pdn;
  assign n1643 = (pv10_1_1_ & n1838_1) | n2095;
  assign n1648 = (n2038 & n1844) | n2094;
  assign n1653 = (n_n4258 & n1839) | n2093_1;
  assign n1658 = ~preset & (n_n3095 | (~pdn & n1870));
  assign n1663 = ~preset & (n_n3663 | (~pdn & n1870));
  assign n1668 = n_n3724 ? n1874 : (n_n3814 & n1836);
  assign n1673 = ~preset & (n_n3038 | (~pdn & n1870));
  assign n1678 = (n_n4337 & n1839) | n2092;
  assign n1683 = (pv11_0_0_ & n1835) | n2091;
  assign n1688 = (pv11_4_4_ & n1835) | n2090;
  assign n1693 = n2089 | (n_n3556 & n_n4122 & n1839);
  assign n1698 = n2088_1 | (n_n4074 & n_n3578 & n1839);
  assign n1703 = ~preset & (n_n3211 | (~pdn & n1870));
  assign n1708 = ~preset & (n_n3367 | (~pdn & n1870));
  assign n1713 = ~preset & (n_n3434 | (~pdn & n1870));
  assign n1718 = n2087 | (n1839 & (n_n4233 | n2338));
  assign n1723 = n2086 | (n_n3688 & n_n3624 & n1839);
  assign n1728 = (n_n3876 & n1839) | n2085;
  assign n1733 = ~preset & (n_n3053 | (~pdn & n1870));
  assign n1738 = ~preset & (n_n3938 | (~pdn & n1870));
  assign n1743 = n2084 | (~preset & n_n3769 & ~n1886);
  assign n1748 = n2083_1 | (n_n3936 & n_n3099 & n1839);
  assign n1753 = n1858_1 | (nsr3_17 & (~nen3_10 | ~n1855));
  assign n1758 = ~preset & (n_n3903 | (~pdn & n1870));
  assign n1763 = n2364 & (n_n3658 | (n1890 & n2322));
  assign n1768 = ~preset & ~ngfdn_3 & (nrq3_11 | ~nsr3_14);
  assign n1773 = n2082 | n2080 | n2081;
  assign n1778 = (pv6_3_3_ & n1846) | n2079;
  assign n1783 = (n_n4316 & n1839) | n2078_1;
  assign n1788 = ~preset & (n_n3175 | (~pdn & n1870));
  assign n1793 = (n_n3657 & n1839) | n2077;
  assign n1798 = n2076 | (n1839 & (n_n3495 | n2341));
  assign n1803 = n2075 | (n1839 & (n_n4095 | n2345));
  assign n1808 = ~preset & (n_n4077 | (~pdn & n1870));
  assign n1813 = ~preset & (n_n3142 | (~pdn & n1870));
  assign n1818 = n2074 | (~preset & n_n3901 & ~n1886);
  assign n1823 = n2072 | (~n_n3934 & n_n3976 & n1840);
  assign n1828 = n2071 | (n_n4227 & ~n1922 & n2315);
  assign n1833 = (n_n4160 & n1839) | n2070;
  assign n1838 = (n_n4182 & n1839) | n2069;
  assign n1843 = (pv4_0_0_ & n1852) | n2068_1;
  assign n1848 = (pv4_4_4_ & n1852) | n2067;
  assign n1853 = ~preset & (n_n3836 | (~pdn & n1870));
  assign n1858 = ~preset & (n_n3470 | (~pdn & n1870));
  assign n1863 = (n_n4157 & n1839) | n2066;
  assign n1868 = (n_n3099 & n1839) | n2065;
  assign n1873 = (pv10_6_6_ & n1838_1) | n2064;
  assign n1878 = (n2038 & n1863_1) | n2063_1;
  assign n1883 = ~preset & ~ngfdn_3 & (ndn3_8 | ndn3_9);
  assign n1888 = (pv1_1_1_ & n1848_1) | n2062;
  assign n1893 = ~preset & (n_n3190 | (~pdn & n1870));
  assign n1898 = n2060 | (n1853_1 & (n2061 | n2365));
  assign n1903 = ~preset & (n_n3042 | (~pdn & n1870));
  assign n1908 = n2059 | preset | pdn;
  assign n1913 = n2058_1 | preset | n2057;
  assign n1918 = ~preset & (n_n3188 | (~pdn & n1870));
  assign n1923 = n2056 | (n_n3769 & n1839 & n1890);
  assign n1928 = (pv11_3_3_ & n1835) | n2055;
  assign n1933 = (pv11_7_7_ & n1835) | n2054;
  assign n1938 = (n_n3916 & n1839) | n2053_1;
  assign n1943 = n2052 | (n1839 & (n_n3608 | n2324));
  assign n1948 = n2051 | (n1839 & (n_n4392 | n2339));
  assign n1953 = ~preset & (n_n3150 | (~pdn & n1870));
  assign n1958 = (n_n3688 & n1839) | n2050;
  assign n1963 = (pv10_7_7_ & n1838_1) | n2049;
  assign n1968 = (n_n4362 & n1839) | n2048_1;
  assign n1973 = n2047 | (n_n3242 & n_n3170 & n1839);
  assign n1978 = n2046 | (n_n4275 & ~n1922 & n2315);
  assign n1983 = n2045 | (n1836 & n2366);
  assign n1988 = (pv2_4_4_ & n1854) | n2044;
  assign n1993 = (pv2_6_6_ & n1854) | n2043_1;
  assign n1998 = n2042 | (n_n3814 & ~n1922 & n2315);
  assign n2003 = n2041 | (n1839 & (~n_n4159 ^ ~n_n3976));
  assign n2008 = (n_n4270 & n1839) | n2040;
  assign n2013 = n2039 | (n1845 & (n1972 ^ n1973_1));
  assign n2018 = (n_n3841 & n1839) | n2038_1;
  assign n2023 = n2036 | n2037;
  assign n2028 = ~preset & (n_n3863 | (~pdn & n1870));
  assign n2033 = ~preset & (n_n3720 | (~pdn & n1870));
  assign n2038 = ~ngfdn_3 & ~preset & nrq3_11;
  assign n2043 = (pv10_0_0_ & n1838_1) | n2035;
  assign n2048 = n2034 | (n1839 & (n_n3458 | n2332));
  assign n2053 = (n_n4299 & n1839) | n2033_1;
  assign n2058 = ~preset & (n_n3529 | (~pdn & n1870));
  assign n2063 = (n_n3756 & n1839) | n2032;
  assign n2068 = n_n4324 ? (n1841 | (n1840 & n1994)) : (n1840 & ~n1994);
  assign n2073 = n2031 | (n_n3035 & n_n4157 & n1839);
  assign n2078 = n2030 | (n_n4227 & (n1874 | n2136));
  assign n2083 = ~preset & (n_n4153 | (~pdn & n1870));
  assign n2088 = n2029 | n2368;
  assign n2093 = ~preset & (n_n3233 | (~pdn & n1870));
  assign n2098 = ~preset & n1881;
  assign n2103 = (n_n4251 & n1839) | n2028_1;
  assign n2108 = (pv4_3_3_ & n1852) | n2027;
  assign n2113 = n2025 | n2026;
  assign n2118 = ~preset & (n_n3441 | (~pdn & n1870));
  assign n2123 = ~preset & ~n1855 & (n_n4026 | n2024);
  assign n2128 = (n_n4229 & n1839) | n2023_1;
  assign n2133 = (n_n3841 & n1839) | n2022;
  assign n2138 = n2021 | (n1839 & (n_n4288 | n2319));
  assign n2143 = n2020 | (n_n3085 & n_n3250 & n1839);
  assign n2148 = (pv1_0_0_ & n1848_1) | n2019;
  assign n2153 = (pv2_0_0_ & n1854) | n2018_1;
  assign n2158 = n2016 | (n1853_1 & (n2017 | n2369));
  assign n2163 = n2014 | (n1853_1 & (n2015 | n2370));
  assign n2168 = (n_n3533 & n1839) | n2013_1;
  assign n2173 = n1882 & ~preset & n_n4057;
  assign n2178 = ~preset & (n_n3674 | (~pdn & n1870));
  assign n2183 = n2011 | (n_n3959 & n1884) | n2010;
  assign n2188 = n2009 | (n1851 & (n1972 ^ n1973_1));
  assign n2193 = n2008_1 | n2006 | n2007;
  assign n2198 = ~preset & (n_n4018 | (~pdn & n1870));
  assign n2203 = ~preset & (n_n4354 | (~pdn & n1870));
  assign n2208 = ~preset & (n_n3797 | (~pdn & n1870));
  assign n2213 = (n_n4316 & n1839) | n2005;
  assign n2218 = n2004 | (n1839 & (n_n4392 | n2339));
  assign n2223 = n2003_1 | (n2038 & (~n1905 ^ n1978_1));
  assign n2228 = n2002 | (n_n4211 & n_n3657 & n1839);
  assign n2233 = n2001 | (n_n4074 & n_n3578 & n1839);
  assign n2238 = ~preset & (n_n3087 | (~pdn & n1870));
  assign n2243 = ~preset & (n_n4105 | (~pdn & n1870));
  assign n2248 = ~preset & (n_n3262 | (~pdn & n1870));
  assign n2253 = (n1886 & n2371) | (~preset & n_n4125 & ~n1886);
  assign n2258 = n2000 | (~n_n3814 & n1836);
  assign n2263 = ~n2374 | (~n1997 & (~n1878_1 | ~n2372));
  assign n2268 = n1858_1 | (nsr3_3 & (~n1956 | n1996));
  assign n1835 = ~ndn3_9 & ~preset & ndn3_8;
  assign n1836 = n_n3709 & n_n3707 & ~preset & ~n_n3198;
  assign n1837 = (~n_n3658 & (n1892 ? n2322 : n_n3604)) | (n_n3604 & (n_n3658 | ~n2322));
  assign n1838_1 = ~ndn3_8 & ~preset & ndn3_7;
  assign n1839 = ~n1889 & ~nsr1_2 & ~preset & ~pdn;
  assign n1840 = n_n4056 & ~n_n3557 & ~preset & n_n4057;
  assign n1841 = ~preset & ~n1886;
  assign n1842 = n_n4108 | (pdn & ~ndn1_34) | (~pdn & n1870);
  assign n1843_1 = ~n_n3916 ^ n1930;
  assign n1844 = n1979 ? ((n1906 & ~n1971) | (n1905 & (n1906 | ~n1971))) : ((~n1906 & n1971) | (~n1905 & (~n1906 | n1971)));
  assign n1845 = nen3_10 & ~preset & ~ndn3_10;
  assign n1846 = ~ndn3_7 & ~preset & ndn3_6;
  assign n1847 = ~nsr3_3 | ndn3_4 | (pready_0_0_ & n1956);
  assign n1848_1 = n2328 & (~nsr3_3 | (pready_0_0_ & n1956));
  assign n1849 = (n1857 & n1977) | (~n_n4360 & ((n1857 & n1960) | n1977));
  assign n1850 = n1897 | ~n2316 | n_n4067 | (~n_n4067 & n1922);
  assign n1851 = ngfdn_3 & ~preset & ~ndn3_15;
  assign n1852 = ~ndn3_6 & ~preset & ndn3_5;
  assign n1853_1 = ~preset & (n1886 | n1900);
  assign n1854 = ~ndn3_5 & ~preset & ndn3_4;
  assign n1855 = ~n_n4093 | (n1903_1 & (n1897 | n2310));
  assign n1856 = ((~n_n3916 ^ n_n4040) & (~n1913_1 ^ ~n1930)) | ((~n_n3916 ^ ~n_n4040) & (n1913_1 ^ ~n1930));
  assign n1857 = ~n_n3841 ^ n1901;
  assign n1858_1 = preset | pdn;
  assign n1859 = nlc1_2 | (~preset_0_0_ & nsr1_2 & (~nlc1_2 | n_n4151));
  assign n1860 = n_n4316 ? (~n1938_1 ^ n1959) : (n1938_1 ^ n1959);
  assign n1861 = ((~n_n3988 ^ n_n3898) & (~n1896 ^ ~n1914)) | ((~n_n3988 ^ ~n_n3898) & (n1896 ^ ~n1914));
  assign n1862 = n2349 & n_n4012 & n1836 & n1867;
  assign n1863_1 = n1912 ? ((n1910 & n1911) | (n1909 & (n1910 | n1911))) : ((~n1910 & ~n1911) | (~n1909 & (~n1910 | ~n1911)));
  assign n1864 = 1'b1;
  assign n1865 = n_n4067 | (~n1897 & ~n1922 & n2316);
  assign n1866 = ~n_n4145 ^ n1895;
  assign n1867 = n_n3724 & n_n4227 & n_n3814;
  assign n1868_1 = n1874 | n2134 | n2135 | n2136;
  assign n1869 = ~n_n3898 ^ n1896;
  assign n1870 = ~nsr1_2 | (preset_0_0_ & ~nlc1_2) | (nlc1_2 & ~n_n4151);
  assign n1871 = ((~n_n4160 ^ ~n_n4222) & (~n_n4159 | (n_n4159 & n_n3976))) | (n_n4159 & ~n_n3976 & (~n_n4160 ^ n_n4222));
  assign n1872 = n2172 | (n2318 & (~n1878_1 | ~n2317));
  assign n1873_1 = ~n_n4229 ^ n1902;
  assign n1874 = n2137 | (n2318 & (~n1878_1 | ~n2317));
  assign n1875 = ((~n_n4229 ^ n_n3818) & (~n1902 ^ ~n1944)) | ((~n_n4229 ^ ~n_n3818) & (n1902 ^ ~n1944));
  assign n1876 = ~n_n4159 ^ ~n_n3976;
  assign n1877 = nrq3_11 & ~ngfdn_3;
  assign n1878_1 = n2316 & ~n1897 & ~n2310;
  assign n1879 = n_n3831 & ((n_n3851 & (n_n4026 | n1953_1)) | (~n_n4026 & n1953_1));
  assign n1880 = ~n2331 | ~n_n3709 | (n1983_1 & n1984);
  assign n1881 = n_n4263 | (~nlc3_3 & n1956 & n2347);
  assign n1882 = n1899 | (n_n4056 & (n1950 | ~n2357));
  assign n1883_1 = n_n3959 | (n_n4159 & n_n3976) | (~n_n4159 & ~n_n3976);
  assign n1884 = n2012 | (n2318 & (~n1878_1 | ~n2317));
  assign n1885 = ((~n_n4145 ^ n_n4080) & (~n1895 ^ ~n1907)) | ((~n_n4145 ^ ~n_n4080) & (n1895 ^ ~n1907));
  assign n1886 = n_n4056 ? n2323 : (n1890 & n2322);
  assign n1887 = (n_n3934 & n_n3976 & (n_n4222 ^ ~n_n4125)) | ((~n_n3934 | ~n_n3976) & (n_n4222 ^ n_n4125));
  assign n1888_1 = n_n4159 | n_n4160 | n_n4383;
  assign n1889 = nlc1_2 ? ~n_n4151 : preset_0_0_;
  assign n1890 = n_n3658 ? n_n3604 : (n2320 | n2321);
  assign n1891 = n_n3955 | ~n_n3954 | n_n4029 | n_n3845;
  assign n1892 = n2320 | n2321;
  assign n1893_1 = (~n1856 & n1955) | (n1843_1 & (n1955 | (~n1856 & n1942)));
  assign n1894 = (n1869 & n1893_1) | (~n1861 & (n1893_1 | (n1869 & n1968_1)));
  assign n1895 = n1931 ? ((n_n3898 & (n1932 | n1933_1)) | (n1932 & n1933_1)) : ((~n1932 & ~n1933_1) | (~n_n3898 & (~n1932 | ~n1933_1)));
  assign n1896 = n1932 ? ((n_n3916 & (n1962 | n1975)) | (n1962 & n1975)) : ((~n1962 & ~n1975) | (~n_n3916 & (~n1962 | ~n1975)));
  assign n1897 = n_n4067 ? ~n_n3833 : n1849;
  assign n1898_1 = n_n4056 & n_n4057 & ~n_n3557;
  assign n1899 = n2322 & ~n_n4056 & n1890;
  assign n1900 = ~n_n3493 & (~n_n4045 | (~n1890 & n2335));
  assign n1901 = n1947 ? ((n1931 & n1934) | (n_n4145 & (n1931 | n1934))) : ((~n1931 & ~n1934) | (~n_n4145 & (~n1931 | ~n1934)));
  assign n1902 = n1927 ? ((n_n4316 & (n1938_1 | n1959)) | (n1938_1 & n1959)) : ((~n1938_1 & ~n1959) | (~n_n4316 & (~n1938_1 | ~n1959)));
  assign n1903_1 = nen3_10 & nsr3_17;
  assign n1904 = ~ndn3_15 & ngfdn_3;
  assign n1905 = n2296 | n2294 | n2295;
  assign n1906 = n2325 | (nrq3_11 & ~ngfdn_3 & n1871);
  assign n1907 = (n_n3988 & n1914) | ((n_n3988 | n1914) & (n_n3898 ^ n1896));
  assign n1908_1 = (n_n4080 & n1907) | ((n_n4080 | n1907) & (~n_n4145 ^ ~n1895));
  assign n1909 = (n1957 & n1958_1) | ((n1957 | n1958_1) & (n2272 | n2273));
  assign n1910 = n2334 | (n1877 & (~n_n3916 ^ n1930));
  assign n1911 = n2265 | n2263_1 | n2264;
  assign n1912 = (~n1918_1 & ~n2221 & ~n2222 & ~n2223_1) | (n1918_1 & (n2221 | n2222 | n2223_1));
  assign n1913_1 = (n_n3818 & n1944) | ((n_n3818 | n1944) & (~n_n4229 ^ ~n1902));
  assign n1914 = (n_n4040 & n1913_1) | ((n_n4040 | n1913_1) & (n_n3916 ^ n1930));
  assign n1915 = n2287 | n2285 | n2286;
  assign n1916 = n2327 | n1915 | n2284;
  assign n1917 = ~n_n3865 ^ n1891;
  assign n1918_1 = n2343 | (n1877 & (~n_n3898 ^ n1896));
  assign n1919 = n_n3709 & ~n_n3198 & n_n3707;
  assign n1920 = n2342 | (n1877 & (~n_n3841 ^ n1901));
  assign n1921 = n2226 | n2224 | n2225;
  assign n1922 = n_n4026 ? ~n_n3851 : ~n1953_1;
  assign n1923_1 = (n_n4047 & n1929) | (n_n3916 & (n_n4047 | n1929));
  assign n1924 = (n_n3898 & n1923_1) | (n_n4366 & (n_n3898 | n1923_1));
  assign n1925 = (n1843_1 & n1964) | (~n_n3876 & (n1964 | (n1843_1 & n1981)));
  assign n1926 = (n1869 & n1925) | (~n_n4362 & (n1925 | (n1869 & n1965)));
  assign n1927 = (~n_n4182 & (n_n4160 | n_n4383 | n_n4159)) | (~n_n4160 & ~n_n4383 & ~n_n4159 & n_n4182);
  assign n1928_1 = (~n1940 & ~n2214 & ~n2215 & ~n2216) | (n1940 & (n2214 | n2215 | n2216));
  assign n1929 = (n_n3769 & n1976) | (n_n4229 & (n_n3769 | n1976));
  assign n1930 = n1962 ? ((n1927 & n1982) | (n_n4229 & (n1927 | n1982))) : ((~n1927 & ~n1982) | (~n_n4229 & (~n1927 | ~n1982)));
  assign n1931 = (~n_n4251 & (n_n4224 | n1888_1 | ~n2314)) | (~n_n4224 & n_n4251 & ~n1888_1 & n2314);
  assign n1932 = (~n_n4224 & (n_n4330 | n_n4182 | n1888_1)) | (n_n4224 & ~n_n4330 & ~n_n4182 & ~n1888_1);
  assign n1933_1 = (n_n3916 & n1975) | ((n_n3916 | n1975) & (n_n4330 ^ n1961));
  assign n1934 = (n1932 & n1933_1) | (n_n3898 & (n1932 | n1933_1));
  assign n1935 = (n_n4222 & ((n_n3934 & n_n3976) | n_n4125)) | (n_n3934 & n_n3976 & n_n4125);
  assign n1936 = (n_n3574 & (n_n3959 ? ~n1871 : (n1871 & n1876))) | (~n1871 & (~n_n3959 | ~n1876)) | (~n_n3574 & n1871 & ~n1876);
  assign n1937 = n1983_1 & (~n1857 | (n1857 & (~n_n3726 ^ ~n1908_1)));
  assign n1938_1 = (~n_n4160 & n_n4383 & ~n_n4159) | (~n_n4383 & (n_n4160 | n_n4159));
  assign n1939 = n1918_1 | n2221 | n2222 | n2223_1;
  assign n1940 = n2344 | (n1877 & (~n_n4145 ^ n1895));
  assign n1941 = (n_n3995 & (n1860 ? (n1936 & ~n1943_1) : (~n1936 & n1943_1))) | (~n1860 & n1936) | (~n_n3995 & (n1860 ? (n1936 & n1943_1) : (~n1936 & ~n1943_1)));
  assign n1942 = (n1875 & n1941) | (~n1873_1 & (n1941 | (n1875 & n1954)));
  assign n1943_1 = (~n1871 & n1883_1) | (n_n3574 & (~n1871 | n1883_1));
  assign n1944 = (~n1860 & n1943_1) | (n_n3995 & (~n1860 | n1943_1));
  assign n1945 = (~n_n4381 & ~n_n4052 & ~n_n3865 & ~n1891) | (n_n4381 & (n_n4052 | n_n3865 | n1891));
  assign n1946 = n_n4224 | n_n4251 | n1888_1 | ~n2314;
  assign n1947 = ~n_n4270 ^ ~n1946;
  assign n1948_1 = (~n_n3955 & n_n3954 & ~n_n4029 & ~n_n3845) | (n_n4029 & (n_n3955 | ~n_n3954 | n_n3845));
  assign n1949 = (~n_n3955 & n_n3954 & ~n_n3845) | (n_n3845 & (n_n3955 | ~n_n3954));
  assign n1950 = ~n_n4099 ^ n1967;
  assign n1951 = n_n4052 ^ (n_n3865 | n1891);
  assign n1952 = ~n1957 ^ (n2268_1 | n2333);
  assign n1953_1 = (~n1857 & n1960) | (n_n4360 & (n1960 | (~n1857 & n1977)));
  assign n1954 = (n_n3995 & (n1860 ? (n1936 & n1943_1) : (~n1936 & ~n1943_1))) | (n1860 & ~n1936) | (~n_n3995 & (n1860 ? (n1936 & ~n1943_1) : (~n1936 & n1943_1)));
  assign n1955 = (~n1875 & n1954) | (n1873_1 & (n1954 | (~n1875 & n1941)));
  assign n1956 = nsr1_2 & ((nlc1_2 & n_n4151) | (~preset_0_0_ & (~nlc1_2 | n_n4151)));
  assign n1957 = n2271 | n2269 | n2270;
  assign n1958_1 = n2333 | (n1877 & (~n_n4229 ^ n1902));
  assign n1959 = (n_n4159 & ((n_n4222 & n_n3976) | (~n_n4160 & (n_n4222 | n_n3976)))) | (n_n4160 & n_n4222 & ~n_n4159);
  assign n1960 = (~n1866 & n1966) | (n_n4299 & (n1966 | (~n1866 & n1926)));
  assign n1961 = n_n4160 | n_n4383 | n_n4159 | n_n4182;
  assign n1962 = ~n_n4330 ^ ~n1961;
  assign n1963_1 = (n1860 & n1985) | (~n_n3946 & (n1985 | (n1860 & ~n1985)));
  assign n1964 = (n1873_1 & n1963_1) | (~n_n4258 & (n1963_1 | (n1873_1 & n1980)));
  assign n1965 = (~n1843_1 & n1981) | (n_n3876 & (n1981 | (~n1843_1 & n1964)));
  assign n1966 = (~n1869 & n1965) | (n_n4362 & (n1965 | (~n1869 & n1925)));
  assign n1967 = n_n4381 | n_n4052 | n_n3865 | n1891;
  assign n1968_1 = (n1856 & n1942) | (~n1843_1 & (n1942 | (n1856 & n1955)));
  assign n1969 = (~n1869 & n1968_1) | (n1861 & (n1968_1 | (~n1869 & n1893_1)));
  assign n1970 = n2216 | n2214 | n2215;
  assign n1971 = ~n1973_1 | (~n2289 & ~n2290 & ~n2291);
  assign n1972 = n2291 | n2289 | n2290;
  assign n1973_1 = n2326 | (n_n3934 & n1890 & n1904);
  assign n1974 = (~n1910 & ~n2263_1 & ~n2264 & ~n2265) | (n1910 & (n2263_1 | n2264 | n2265));
  assign n1975 = (n1927 & n1982) | (n_n4229 & (n1927 | n1982));
  assign n1976 = (n_n3901 & n1935) | (n_n4316 & (n_n3901 | n1935));
  assign n1977 = (n1866 & n1926) | (~n_n4299 & (n1926 | (n1866 & n1966)));
  assign n1978_1 = (n1972 & n1973_1 & (n2293 | n2325)) | (~n2293 & (~n1972 | ~n1973_1) & ~n2325);
  assign n1979 = ~n1915 ^ (n2284 | n2327);
  assign n1980 = (~n1860 & ~n1985) | (n_n3946 & (~n1985 | (~n1860 & n1985)));
  assign n1981 = (~n1873_1 & n1980) | (n_n4258 & (n1980 | (~n1873_1 & n1963_1)));
  assign n1982 = (n1938_1 & n1959) | (n_n4316 & (n1938_1 | n1959));
  assign n1983_1 = (n1885 & n1969) | (~n1866 & ((n1885 & n1894) | n1969));
  assign n1984 = (~n_n3841 & n1901) | (n_n3841 & ~n1901) | ((~n_n3841 ^ n1901) & (n_n3726 ^ n1908_1));
  assign n1985 = (n1871 & n2313) | (~n_n3743 & (n1871 | n2313));
  assign n1986 = (~n1970 & ~n2218_1 & ~n2219) | (~n1940 & (~n1970 | (~n2218_1 & ~n2219)));
  assign n1987 = n1897 | n2310 | ~n2316 | n2340;
  assign n1988_1 = ndn3_4 | (nsr3_3 & (~pready_0_0_ | ~n1956));
  assign n1989 = n1890 & ~n_n3493 & ~n_n4045;
  assign n1990 = n_n4145 ? ((n_n4366 & (n_n3898 | n1923_1)) | (n_n3898 & n1923_1)) : ((~n_n3898 & ~n1923_1) | (~n_n4366 & (~n_n3898 | ~n1923_1)));
  assign n1991 = n_n3898 ? ((n_n4047 & n1929) | (n_n3916 & (n_n4047 | n1929))) : ((~n_n4047 & ~n1929) | (~n_n3916 & (~n_n4047 | ~n1929)));
  assign n1992 = n_n4047 ? ((n_n3769 & n1976) | (n_n4229 & (n_n3769 | n1976))) : ((~n_n3769 & ~n1976) | (~n_n4229 & (~n_n3769 | ~n1976)));
  assign n1993_1 = n_n3769 ? ((n_n4316 & (n_n3901 | n1935)) | (n_n3901 & n1935)) : ((~n_n3901 & ~n1935) | (~n_n4316 & (~n_n3901 | ~n1935)));
  assign n1994 = n_n3841 ? ((n_n4145 & n1924) | (n_n3475 & (n_n4145 | n1924))) : ((~n_n4145 & ~n1924) | (~n_n3475 & (~n_n4145 | ~n1924)));
  assign n1995 = ~n_n3707 | (~n_n4026 & ~n1953_1) | (~n_n3851 & n_n4026);
  assign n1996 = nsr4_2 & ((n_n4108 & ~n_n3354) | (~tin_pready_0_0_ & (~n_n4108 | ~n_n3354)));
  assign n1997 = ~preset & (~n_n3831 | n1998_1 | n1999);
  assign n1998_1 = n2373 & n2316 & ~n1897 & ~n2310;
  assign n1999 = n2316 & ~n2310 & ~n1897 & n1995;
  assign n2000 = n_n3814 & (~n1878_1 | ~n2317) & n2318;
  assign n2001 = ~preset & n_n3806 & (pdn | ~n1870);
  assign n2002 = ~preset & n_n3537 & (pdn | ~n1870);
  assign n2003_1 = ~preset & n_n3099 & (~nrq3_11 | ngfdn_3);
  assign n2004 = ~preset & n_n3646 & (pdn | ~n1870);
  assign n2005 = ~preset & n_n3739 & (pdn | ~n1870);
  assign n2006 = n2317 & n1878_1 & ~preset & n_n4299;
  assign n2007 = n_n4080 & (~n1878_1 | ~n2317) & n2318;
  assign n2008_1 = n1836 & (n_n4080 ? (~n1866 ^ ~n1907) : (n1866 ^ ~n1907));
  assign n2009 = ~preset & n_n3608 & (ndn3_15 | ~ngfdn_3);
  assign n2010 = n2317 & n1878_1 & ~preset & n_n3756;
  assign n2011 = ~n_n3959 & n1836 & (~n_n4159 ^ ~n_n3976);
  assign n2012 = n1836 & (~n_n4159 ^ n_n3976);
  assign n2013_1 = ~preset & n_n3486 & (pdn | ~n1870);
  assign n2014 = ~n1900 & ~n1886 & ~preset & n_n3865;
  assign n2015 = n_n3922 & (n1899 | n2259);
  assign n2016 = ~n1900 & ~n1886 & ~preset & n_n3845;
  assign n2017 = n_n3968 & (n1899 | n2259);
  assign n2018_1 = ~preset & n_n3931 & (~ndn3_4 | ndn3_5);
  assign n2019 = n1988_1 & ~preset & n_n3878;
  assign n2020 = ~preset & n_n4180 & (pdn | ~n1870);
  assign n2021 = ~preset & n_n3277 & (pdn | ~n1870);
  assign n2022 = ~preset & n_n4102 & (pdn | ~n1870);
  assign n2023_1 = ~preset & n_n4342 & (pdn | ~n1870);
  assign n2024 = n2316 & ~n2310 & n1879 & ~n1897;
  assign n2025 = ~preset & n_n3841 & (ndn3_10 | ~nen3_10);
  assign n2026 = n1845 & (n1920 ? (~n1921 ^ ~n1986) : (n1921 ^ ~n1986));
  assign n2027 = ~preset & n_n4182 & (~ndn3_5 | ndn3_6);
  assign n2028_1 = ~preset & n_n3413 & (pdn | ~n1870);
  assign n2029 = n_n3831 & (n1897 | n2310 | ~n2316);
  assign n2030 = n1836 & n_n3814 & n_n3724 & ~n_n4227;
  assign n2031 = ~preset & n_n3337 & (pdn | ~n1870);
  assign n2032 = ~preset & n_n4209 & (pdn | ~n1870);
  assign n2033_1 = ~preset & n_n3342 & (pdn | ~n1870);
  assign n2034 = ~preset & n_n3667 & (pdn | ~n1870);
  assign n2035 = ~preset & n_n3756 & (~ndn3_7 | ndn3_8);
  assign n2036 = ~preset & n_n4095 & (ndn3_15 | ~ngfdn_3);
  assign n2037 = n1851 & (n1928_1 ^ (~n2218_1 & ~n2219));
  assign n2038_1 = ~preset & n_n3394 & (pdn | ~n1870);
  assign n2039 = ~preset & n_n3976 & (ndn3_10 | ~nen3_10);
  assign n2040 = ~preset & n_n4166 & (pdn | ~n1870);
  assign n2041 = ~preset & n_n3572 & (pdn | ~n1870);
  assign n2042 = ~preset & n_n3514 & (pdn | ~n1870);
  assign n2043_1 = ~preset & n_n4062 & (~ndn3_4 | ndn3_5);
  assign n2044 = ~preset & n_n4021 & (~ndn3_4 | ndn3_5);
  assign n2045 = n_n3766 & (n1874 | n2135 | n2136);
  assign n2046 = ~preset & n_n3966 & (pdn | ~n1870);
  assign n2047 = ~preset & n_n4199 & (pdn | ~n1870);
  assign n2048_1 = ~preset & n_n4247 & (pdn | ~n1870);
  assign n2049 = ~preset & n_n4360 & (~ndn3_7 | ndn3_8);
  assign n2050 = ~preset & n_n4320 & (pdn | ~n1870);
  assign n2051 = ~preset & n_n3108 & (pdn | ~n1870);
  assign n2052 = ~preset & n_n3910 & (pdn | ~n1870);
  assign n2053_1 = ~preset & n_n3758 & (pdn | ~n1870);
  assign n2054 = ~preset & n_n3170 & (~ndn3_8 | ndn3_9);
  assign n2055 = ~preset & n_n3250 & (~ndn3_8 | ndn3_9);
  assign n2056 = ~preset & n_n4303 & (pdn | ~n1870);
  assign n2057 = nsr1_2 & ~preset_0_0_ & ~nlc1_2;
  assign n2058_1 = n_n4151 & (nlc1_2 | ~nsr1_2 | (preset_0_0_ & ~nlc1_2));
  assign n2059 = nsr3_14 & (nsr3_17 | (n_n4045 & n1890));
  assign n2060 = ~n1900 & ~n1886 & ~preset & n_n4029;
  assign n2061 = n_n3533 & (n1899 | n2259);
  assign n2062 = n1988_1 & ~preset & n_n3208;
  assign n2063_1 = ~preset & n_n4157 & (~nrq3_11 | ngfdn_3);
  assign n2064 = ~preset & n_n4299 & (~ndn3_7 | ndn3_8);
  assign n2065 = ~preset & n_n3883 & (pdn | ~n1870);
  assign n2066 = ~preset & n_n3331 & (pdn | ~n1870);
  assign n2067 = ~preset & n_n4330 & (~ndn3_5 | ndn3_6);
  assign n2068_1 = ~preset & n_n4159 & (~ndn3_5 | ndn3_6);
  assign n2069 = ~preset & n_n4309 & (pdn | ~n1870);
  assign n2070 = ~preset & n_n3722 & (pdn | ~n1870);
  assign n2071 = ~preset & n_n3823 & (pdn | ~n1870);
  assign n2072 = n_n3934 & (n2073_1 | (~preset & ~n1886));
  assign n2073_1 = ~n_n3976 & n1840;
  assign n2074 = n1840 & (n_n4316 ? (~n_n3901 ^ n1935) : (n_n3901 ^ n1935));
  assign n2075 = ~preset & n_n3385 & (pdn | ~n1870);
  assign n2076 = ~preset & n_n3202 & (pdn | ~n1870);
  assign n2077 = ~preset & n_n3055 & (pdn | ~n1870);
  assign n2078_1 = ~preset & n_n3463 & (pdn | ~n1870);
  assign n2079 = ~preset & n_n3533 & (~ndn3_6 | ndn3_7);
  assign n2080 = n2317 & n1878_1 & ~preset & n_n4258;
  assign n2081 = n_n3818 & (~n1878_1 | ~n2317) & n2318;
  assign n2082 = n1836 & (n_n3818 ? (~n1873_1 ^ ~n1944) : (n1873_1 ^ ~n1944));
  assign n2083_1 = ~preset & n_n4390 & (pdn | ~n1870);
  assign n2084 = n1840 & (~n_n4229 ^ n1993_1);
  assign n2085 = ~preset & n_n4136 & (pdn | ~n1870);
  assign n2086 = ~preset & n_n4192 & (pdn | ~n1870);
  assign n2087 = ~preset & n_n3126 & (pdn | ~n1870);
  assign n2088_1 = ~preset & n_n3089 & (pdn | ~n1870);
  assign n2089 = ~preset & n_n3713 & (pdn | ~n1870);
  assign n2090 = ~preset & n_n3578 & (~ndn3_8 | ndn3_9);
  assign n2091 = ~preset & n_n3624 & (~ndn3_8 | ndn3_9);
  assign n2092 = ~preset & n_n3370 & (pdn | ~n1870);
  assign n2093_1 = ~preset & n_n3213 & (pdn | ~n1870);
  assign n2094 = ~preset & n_n3657 & (~nrq3_11 | ngfdn_3);
  assign n2095 = ~preset & n_n3743 & (~ndn3_7 | ndn3_8);
  assign n2096 = ~preset & n_n3223 & (pdn | ~n1870);
  assign n2097 = ~preset & n_n4236 & (pdn | ~n1870);
  assign n2098_1 = ~preset & n_n4372 & (pdn | ~n1870);
  assign n2099 = ~preset & n_n3136 & (pdn | ~n1870);
  assign n2100 = ~n1900 & ~n1886 & ~preset & ~n_n3954;
  assign n2101 = n_n4349 & (n1899 | n2259);
  assign n2102 = n2360 & (~n_n4056 | n1950 | ~n2357);
  assign n2103_1 = n1988_1 & ~preset & n_n3259;
  assign n2104 = ~preset & n_n3085 & (~nrq3_11 | ngfdn_3);
  assign n2105 = n2038 & (n1952 ^ (~n2272 & ~n2273));
  assign n2106 = ~preset & n_n3946 & (~ndn3_7 | ndn3_8);
  assign n2107 = n_n3709 & ((n1983_1 & n1984) | ~n2331);
  assign n2108_1 = ~preset & n_n3777 & (pdn | ~n1870);
  assign n2109 = ~preset & n_n3073 & (pdn | ~n1870);
  assign n2110 = n2349 & n1867 & ~n_n4012 & n1836;
  assign n2111 = ~preset & n_n3436 & (pdn | ~n1870);
  assign n2112 = ~preset & n_n4351 & (ndn3_15 | ~ngfdn_3);
  assign n2113_1 = n1851 & (n1952 ^ (~n2272 & ~n2273));
  assign n2114 = ~preset & n_n3287 & (pdn | ~n1870);
  assign n2115 = ~preset & n_n3679 & (pdn | ~n1870);
  assign n2116 = ~preset & n_n4065 & (pdn | ~n1870);
  assign n2117 = ~preset & n_n3138 & (pdn | ~n1870);
  assign n2118_1 = ~preset & n_n3631 & (pdn | ~n1870);
  assign n2119 = ~preset & n_n3020 & (pdn | ~n1870);
  assign n2120 = ~preset & n_n3057 & (pdn | ~n1870);
  assign n2121 = ~preset & n_n3404 & (pdn | ~n1870);
  assign n2122 = ~preset & n_n3069 & (pdn | ~n1870);
  assign n2123_1 = n_n3483 & (n1872 | n2124 | n2171);
  assign n2124 = ~n_n4334 & n1836;
  assign n2125 = ~preset & n_n4362 & (~ndn3_7 | ndn3_8);
  assign n2126 = ~preset & n_n4201 & (~ndn3_6 | ndn3_7);
  assign n2127 = ~preset & n_n4229 & (ndn3_10 | ~nen3_10);
  assign n2128_1 = n1845 & (n1952 ^ (~n2272 & ~n2273));
  assign n2129 = ~preset & n_n3408 & (pdn | ~n1870);
  assign n2130 = ~preset & n_n3451 & (~ndn3_4 | ndn3_5);
  assign n2131 = n_n4057 & (~n_n4056 | n1950 | ~n2357);
  assign n2132 = ~preset & n_n3854 & (~ndn3_4 | ndn3_5);
  assign n2133_1 = n2354 & (n1919 | (n1878_1 & n2317));
  assign n2134 = ~n_n3766 & n1836;
  assign n2135 = ~n_n4227 & n1836;
  assign n2136 = ~n_n3724 & n1836;
  assign n2137 = ~n_n3814 & n1836;
  assign n2138_1 = ~preset & n_n3922 & (~ndn3_6 | ndn3_7);
  assign n2139 = ~preset & n_n3968 & (~ndn3_6 | ndn3_7);
  assign n2140 = ~preset & n_n3237 & (pdn | ~n1870);
  assign n2141 = ~preset & n_n3952 & (pdn | ~n1870);
  assign n2142 = ~preset & n_n4122 & (~nrq3_11 | ngfdn_3);
  assign n2143_1 = n2038 & (n1928_1 ^ (~n2218_1 & ~n2219));
  assign n2144 = ~preset & n_n3898 & (ndn3_10 | ~nen3_10);
  assign n2145 = ~n1900 & ~n1886 & ~preset & n_n4099;
  assign n2146 = n_n4337 & (n1899 | n2259);
  assign n2147 = ~n1900 & ~n1886 & ~preset & n_n4052;
  assign n2148_1 = n1898_1 & (~n_n4052 ^ (n_n3865 | n1891));
  assign n2149 = n_n4071 & (n1899 | n2259);
  assign n2150 = ~preset & n_n3985 & (pdn | ~n1870);
  assign n2151 = ~preset & n_n3091 & (pdn | ~n1870);
  assign n2152 = ~preset & n_n4003 & (pdn | ~n1870);
  assign n2153_1 = ~preset & n_n4145 & (ndn3_10 | ~nen3_10);
  assign n2154 = n1845 & (n1928_1 ^ (~n2218_1 & ~n2219));
  assign n2155 = ~preset & n_n3978 & (~ndn3_4 | ndn3_5);
  assign n2156 = n1840 & (~n_n3916 ^ n1992);
  assign n2157 = ~preset & n_n3183 & (pdn | ~n1870);
  assign n2158_1 = ~preset & n_n4288 & (ndn3_15 | ~ngfdn_3);
  assign n2159 = ~preset & n_n4270 & (~ndn3_5 | ndn3_6);
  assign n2160 = ~preset & n_n3449 & (pdn | ~n1870);
  assign n2161 = ~preset & n_n3971 & (pdn | ~n1870);
  assign n2162 = ~preset & n_n3429 & (pdn | ~n1870);
  assign n2163_1 = ~preset & n_n3319 & (pdn | ~n1870);
  assign n2164 = ~preset & n_n3506 & (pdn | ~n1870);
  assign n2165 = ~preset & n_n3458 & (ndn3_15 | ~ngfdn_3);
  assign n2166 = ~preset & n_n4233 & (ndn3_15 | ~ngfdn_3);
  assign n2167 = n1851 & (n1920 ? (~n1921 ^ ~n1986) : (n1921 ^ ~n1986));
  assign n2168_1 = ~preset & n_n3155 & (pdn | ~n1870);
  assign n2169 = ~n1900 & ~n1886 & ~preset & n_n3955;
  assign n2170 = n_n4201 & (n1899 | n2259);
  assign n2171 = ~n_n4012 & n1836;
  assign n2172 = n1836 & (~n_n4275 | ~n_n3766 | ~n1867);
  assign n2173_1 = n1988_1 & ~preset & n_n4294;
  assign n2174 = ~preset & n_n4251 & (~ndn3_5 | ndn3_6);
  assign n2175 = ~preset & n_n3736 & (pdn | ~n1870);
  assign n2176 = ~preset & n_n3896 & (pdn | ~n1870);
  assign n2177 = ~preset & n_n4279 & (pdn | ~n1870);
  assign n2178_1 = n2317 & n1878_1 & ~preset & n_n4362;
  assign n2179 = n_n3988 & (~n1878_1 | ~n2317) & n2318;
  assign n2180 = n1836 & (n_n3988 ? (~n1869 ^ ~n1914) : (n1869 ^ ~n1914));
  assign n2181 = ~preset & n_n3328 & (~ndn3_4 | ndn3_5);
  assign n2182 = ~preset & n_n3761 & (pdn | ~n1870);
  assign n2183_1 = n2317 & n1878_1 & ~preset & n_n3946;
  assign n2184 = n_n3995 & (~n1878_1 | ~n2317) & n2318;
  assign n2185 = n1836 & (n_n3995 ? (~n1860 ^ ~n1943_1) : (n1860 ^ ~n1943_1));
  assign n2186 = ~preset & n_n3128 & (pdn | ~n1870);
  assign n2187 = n1988_1 & ~preset & n_n3919;
  assign n2188_1 = n1988_1 & ~preset & n_n3886;
  assign n2189 = ~preset & n_n3048 & (pdn | ~n1870);
  assign n2190 = ~preset & n_n3061 & (pdn | ~n1870);
  assign n2191 = ~preset & n_n3316 & (pdn | ~n1870);
  assign n2192 = ~preset & n_n3906 & (pdn | ~n1870);
  assign n2193_1 = ~preset & n_n3583 & (pdn | ~n1870);
  assign n2194 = ~preset & n_n3358 & (pdn | ~n1870);
  assign n2195 = ~preset & n_n4243 & (pdn | ~n1870);
  assign n2196 = ~preset & n_n4337 & (~ndn3_6 | ndn3_7);
  assign n2197 = ~preset & n_n3207 & (pdn | ~n1870);
  assign n2198_1 = ~preset & n_n3465 & (pdn | ~n1870);
  assign n2199 = n2348 & ((~pdn & ~n1870) | (ndn1_34 & (pdn | ~n1870)));
  assign n2200 = ~preset & n_n3892 & (~ndn3_6 | ndn3_7);
  assign n2201 = ~preset & n_n4383 & (~ndn3_5 | ndn3_6);
  assign n2202 = ~preset & n_n4286 & (pdn | ~n1870);
  assign n2203_1 = ~preset & n_n4189 & (pdn | ~n1870);
  assign n2204 = ~preset & n_n3576 & (pdn | ~n1870);
  assign n2205 = ~preset & n_n4172 & (pdn | ~n1870);
  assign n2206 = ~preset & n_n3111 & (pdn | ~n1870);
  assign n2207 = ~preset & n_n3035 & (~ndn3_8 | ndn3_9);
  assign n2208_1 = ~preset & n_n3627 & (pdn | ~n1870);
  assign n2209 = ~preset & n_n3044 & (pdn | ~n1870);
  assign n2210 = ~preset & n_n3376 & (pdn | ~n1870);
  assign n2211 = ~preset & n_n3118 & (pdn | ~n1870);
  assign n2212 = ~preset & n_n3242 & (~nrq3_11 | ngfdn_3);
  assign n2213_1 = n2038 & (n1920 ? (~n1921 ^ ~n1986) : (n1921 ^ ~n1986));
  assign n2214 = ngfdn_3 & n_n4122 & ~ndn3_15 & n_n3556;
  assign n2215 = nen3_10 & ~ndn3_10 & n_n3919;
  assign n2216 = n_n4145 & nrq3_11 & ~ngfdn_3;
  assign n2217 = n_n4062 & ~ndn3_10 & nen3_10;
  assign n2218_1 = n1939 & ((n1910 & n1911) | (n1909 & (n1910 | n1911)));
  assign n2219 = n1918_1 & (n2221 | n2222 | n2223_1);
  assign n2220 = nen3_10 & ~ndn3_10 & n_n3854;
  assign n2221 = ngfdn_3 & n_n4157 & ~ndn3_15 & n_n3035;
  assign n2222 = nen3_10 & n_n3511 & ~ndn3_10;
  assign n2223_1 = n_n3898 & nrq3_11 & ~ngfdn_3;
  assign n2224 = ngfdn_3 & n_n3170 & ~ndn3_15 & n_n3242;
  assign n2225 = n_n3259 & ~ndn3_10 & nen3_10;
  assign n2226 = n_n3841 & nrq3_11 & ~ngfdn_3;
  assign n2227 = nen3_10 & ~ndn3_10 & n_n3451;
  assign n2228_1 = ~preset & n_n3113 & (pdn | ~n1870);
  assign n2229 = ~preset & n_n3173 & (pdn | ~n1870);
  assign n2230 = ~preset & n_n3221 & (pdn | ~n1870);
  assign n2231 = n2317 & n1878_1 & ~preset & n_n3876;
  assign n2232 = n_n4040 & (~n1878_1 | ~n2317) & n2318;
  assign n2233_1 = n1836 & (n_n4040 ? (~n1843_1 ^ ~n1913_1) : (n1843_1 ^ ~n1913_1));
  assign n2234 = ~preset & n_n3556 & (~ndn3_8 | ndn3_9);
  assign n2235 = ~preset & n_n3733 & (pdn | ~n1870);
  assign n2236 = ~preset & n_n3231 & (pdn | ~n1870);
  assign n2237 = ~preset & n_n3313 & (pdn | ~n1870);
  assign n2238_1 = ~preset & n_n3079 & (pdn | ~n1870);
  assign n2239 = ~preset & n_n3688 & (~nrq3_11 | ngfdn_3);
  assign n2240 = ~preset & n_n3344 & (pdn | ~n1870);
  assign n2241 = ~preset & n_n4071 & (~ndn3_6 | ndn3_7);
  assign n2242 = ~preset & n_n3012 & (pdn | ~n1870);
  assign n2243_1 = ~preset & n_n4222 & (ndn3_10 | ~nen3_10);
  assign n2244 = ~preset & n_n4160 & (~ndn3_5 | ndn3_6);
  assign n2245 = ~preset & n_n3517 & (pdn | ~n1870);
  assign n2246 = n_n3707 & (~n_n3709 | n1937 | ~n2331);
  assign n2247 = ~preset & n_n3281 & (~ndn3_4 | ndn3_5);
  assign n2248_1 = ~preset & n_n3764 & (pdn | ~n1870);
  assign n2249 = ~preset & n_n3549 & (pdn | ~n1870);
  assign n2250 = ~preset & n_n3876 & (~ndn3_7 | ndn3_8);
  assign n2251 = ~preset & n_n3729 & (pdn | ~n1870);
  assign n2252 = ~preset & n_n3525 & (pdn | ~n1870);
  assign n2253_1 = ~preset & n_n3916 & (ndn3_10 | ~nen3_10);
  assign n2254 = ~preset & n_n3495 & (ndn3_15 | ~ngfdn_3);
  assign n2255 = ~preset & n_n4211 & (~ndn3_8 | ndn3_9);
  assign n2256 = ~preset & n_n3670 & (pdn | ~n1870);
  assign n2257 = ~n1900 & ~n1886 & ~preset & n_n4381;
  assign n2258_1 = n_n3892 & (n1899 | n2259);
  assign n2259 = ~n_n3493 & ~n1890 & (~n_n4045 | n2335);
  assign n2260 = n1988_1 & ~preset & n_n3858;
  assign n2261 = ~preset & n_n3270 & (pdn | ~n1870);
  assign n2262 = ~preset & n_n4074 & (~nrq3_11 | ngfdn_3);
  assign n2263_1 = ngfdn_3 & n_n3578 & ~ndn3_15 & n_n4074;
  assign n2264 = nen3_10 & ~ndn3_10 & n_n3886;
  assign n2265 = n_n3916 & nrq3_11 & ~ngfdn_3;
  assign n2266 = n_n4021 & ~ndn3_10 & nen3_10;
  assign n2267 = nen3_10 & n_n3281 & ~ndn3_10;
  assign n2268_1 = nrq3_11 & ~ngfdn_3 & (n_n4229 ^ ~n1902);
  assign n2269 = ngfdn_3 & n_n3250 & ~ndn3_15 & n_n3085;
  assign n2270 = nen3_10 & ~ndn3_10 & n_n4294;
  assign n2271 = n_n4229 & nrq3_11 & ~ngfdn_3;
  assign n2272 = n1916 & ((n1906 & ~n1971) | (n1905 & (n1906 | ~n1971)));
  assign n2273 = n1915 & (n2284 | n2327);
  assign n2274 = ~preset & n_n3133 & (pdn | ~n1870);
  assign n2275 = ~n1894 & (~n1969 | n2329);
  assign n2276 = (~n_n4145 ^ ~n1895) & (~n_n4080 ^ n1907);
  assign n2277 = ~preset & n_n4224 & (~ndn3_5 | ndn3_6);
  assign n2278 = ~preset & n_n4392 & (ndn3_15 | ~ngfdn_3);
  assign n2279 = n1988_1 & ~preset & n_n3511;
  assign n2280 = ~preset & n_n3780 & (pdn | ~n1870);
  assign n2281 = ~preset & n_n4349 & (~ndn3_6 | ndn3_7);
  assign n2282 = ~preset & n_n4316 & (ndn3_10 | ~nen3_10);
  assign n2283 = nen3_10 & ~ndn3_10 & n_n3978;
  assign n2284 = n1877 & (n_n4316 ? (n1938_1 ^ ~n1959) : (~n1938_1 ^ ~n1959));
  assign n2285 = ngfdn_3 & n_n3657 & ~ndn3_15 & n_n4211;
  assign n2286 = nen3_10 & n_n3858 & ~ndn3_10;
  assign n2287 = n_n4316 & nrq3_11 & ~ngfdn_3;
  assign n2288 = nrq3_11 & ~ngfdn_3 & (n_n4159 ^ n_n3976);
  assign n2289 = ngfdn_3 & n_n3624 & ~ndn3_15 & n_n3688;
  assign n2290 = n_n3878 & ~ndn3_10 & nen3_10;
  assign n2291 = nrq3_11 & n_n3976 & ~ngfdn_3;
  assign n2292 = nen3_10 & ~ndn3_10 & n_n3328;
  assign n2293 = n1871 & nrq3_11 & ~ngfdn_3;
  assign n2294 = n_n3099 & ngfdn_3 & n_n3936 & ~ndn3_15;
  assign n2295 = n_n3208 & ~ndn3_10 & nen3_10;
  assign n2296 = n_n4222 & nrq3_11 & ~ngfdn_3;
  assign n2297 = ~preset & n_n3793 & (pdn | ~n1870);
  assign n2298 = ~preset & n_n3497 & (pdn | ~n1870);
  assign n2299 = ~preset & n_n3098 & (pdn | ~n1870);
  assign n2300 = ~preset & n_n3687 & (pdn | ~n1870);
  assign n2301 = ~preset & n_n3225 & (pdn | ~n1870);
  assign n2302 = ~preset & n_n4258 & (~ndn3_7 | ndn3_8);
  assign n2303 = n2317 & n1878_1 & ~preset & n_n4360;
  assign n2304 = n_n3726 & (~n1878_1 | ~n2317) & n2318;
  assign n2305 = n1836 & (n_n3726 ? (~n1857 ^ ~n1908_1) : (n1857 ^ ~n1908_1));
  assign n2306 = ~preset & n_n3008 & (pdn | ~n1870);
  assign n2307 = n2317 & n1878_1 & ~preset & n_n3743;
  assign n2308 = n_n3574 & (~n1878_1 | ~n2317) & n2318;
  assign n2309 = n1836 & (n_n3574 ? (~n1871 ^ ~n1883_1) : (n1871 ^ ~n1883_1));
  assign n2310 = ~n_n4067 & (n_n4026 ? ~n_n3851 : ~n1953_1);
  assign n2311 = ~preset & n_n3936 & (~ndn3_8 | ndn3_9);
  assign n2312 = ~preset & n_n4142 & (pdn | ~n1870);
  assign n2313 = ~n_n3756 & (~n_n4159 ^ ~n_n3976);
  assign n2314 = ~n_n4182 & ~n_n4330;
  assign n2315 = n1839 & ((~n_n4067 & ~n1849) | (n_n3833 & (n_n4067 | ~n1849)));
  assign n2316 = nen3_10 & nsr3_17 & n_n4093;
  assign n2317 = n1879 & ~n_n3709;
  assign n2318 = ~preset & (n_n3198 | ~n_n3707 | ~n_n3709);
  assign n2319 = n_n4157 & n_n3035;
  assign n2320 = n_n4349 | n_n4071 | n_n3892 | n_n4337;
  assign n2321 = n_n3968 | n_n3922 | n_n4201 | n_n3533;
  assign n2322 = nsr3_14 & n_n4045 & ~nsr3_17;
  assign n2323 = ~n_n3557 & n_n4057;
  assign n2324 = n_n3624 & n_n3688;
  assign n2325 = n2292 | (n_n4125 & n1890 & n1904);
  assign n2326 = n2288 | (~ndn3_10 & nen3_10 & n_n3931);
  assign n2327 = n2283 | (n_n3901 & n1890 & n1904);
  assign n2328 = ~ndn3_4 & ~preset;
  assign n2329 = (n_n4145 & ~n1895) | (~n_n4145 & n1895) | ((~n_n4145 ^ n1895) & (n_n4080 ^ n1907));
  assign n2330 = n1857 | n2276 | (~n1857 & (~n_n3726 ^ ~n1908_1));
  assign n2331 = n1919 & (n2275 | n2330);
  assign n2332 = n_n3578 & n_n4074;
  assign n2333 = n2267 | (n_n3769 & n1890 & n1904);
  assign n2334 = n2266 | (n_n4047 & n1890 & n1904);
  assign n2335 = nsr3_14 & ~nsr3_17;
  assign n2336 = (n1898_1 & n1945) | (n_n4381 & n1989);
  assign n2337 = n_n3493 & ~preset;
  assign n2338 = n_n3170 & n_n3242;
  assign n2339 = n_n3099 & n_n3936;
  assign n2340 = n_n4026 | ~n_n3831 | (~n_n4026 & ~n1953_1);
  assign n2341 = n_n3657 & n_n4211;
  assign n2342 = n2227 | (n_n4324 & n1890 & n1904);
  assign n2343 = n2220 | (n_n4366 & n1890 & n1904);
  assign n2344 = n2217 | (n_n3475 & n1890 & n1904);
  assign n2345 = n_n4122 & n_n3556;
  assign n2346 = n_n3250 & n_n3085;
  assign n2347 = nsr3_3 & ((n_n4108 & ~n_n3354) | (~tin_pready_0_0_ & (~n_n4108 | ~n_n3354)));
  assign n2348 = n_n3354 & ~preset;
  assign n2349 = n_n3766 & n_n4275;
  assign n2350 = n_n3955 ? (n1989 | (~n_n3954 & n1898_1)) : (n_n3954 & n1898_1);
  assign n2351 = nlak4_2 | (nlc3_3 & ~n_n4263);
  assign n2352 = (n_n4052 & n1989) | n2148_1;
  assign n2353 = n_n4099 ? ((n1898_1 & n1967) | n1989) : (n1898_1 & ~n1967);
  assign n2354 = n1867 & n1836 & ~n_n4275 & n_n3766;
  assign n2355 = ~n_n3954 & ~n_n3955;
  assign n2356 = n2355 & ~n1949 & n1898_1 & ~n1948_1;
  assign n2357 = n2356 & n1951 & ~n1917 & ~n1945;
  assign n2358 = ~n_n4045 | preset | (~n1890 & n2335);
  assign n2359 = n_n3707 & ~preset;
  assign n2360 = n1890 & n_n4057;
  assign n2361 = ~nsr3_14 | nsr3_17;
  assign n2362 = ~n_n4045 | preset | (~n1890 & n2335);
  assign n2363 = n_n3954 ? n1898_1 : n1989;
  assign n2364 = ~preset & n_n4045 & (n1890 | ~n2335);
  assign n2365 = (n1898_1 & n1948_1) | (n_n4029 & n1989);
  assign n2366 = n_n3814 & n_n4227 & n_n3724 & ~n_n3766;
  assign n2367 = n1879 & n_n3707;
  assign n2368 = n1855 | preset | (n1880 & n2367);
  assign n2369 = (n1898_1 & n1949) | (n_n3845 & n1989);
  assign n2370 = n_n3865 ? ((n1891 & n1898_1) | n1989) : (~n1891 & n1898_1);
  assign n2371 = n1887 & n1840;
  assign n2372 = n2331 & ~n1937 & ~preset & n_n3709;
  assign n2373 = n1849 & ~n_n4067;
  assign n2374 = ~n2310 & n1903_1 & n_n4093 & ~n1897;
  always @ (posedge clock) begin
    n_n4142 <= n349;
    n_n3936 <= n354;
    n_n3574 <= n359;
    n_n3008 <= n364;
    n_n3726 <= n369;
    n_n3604 <= n374;
    n_n3144 <= n379;
    n_n3782 <= n384;
    n_n3067 <= n389;
    n_n4258 <= n394;
    n_n3225 <= n399;
    n_n3180 <= n404;
    n_n3274 <= n409;
    n_n3475 <= n414;
    n_n3687 <= n419;
    n_n3381 <= n424;
    n_n3098 <= n429;
    n_n4108 <= n434;
    n_n3497 <= n439;
    n_n3793 <= n444;
    n_n4316 <= n449;
    n_n4349 <= n454;
    n_n3029 <= n459;
    n_n3619 <= n464;
    n_n3264 <= n469;
    n_n3780 <= n474;
    ndn3_4 <= n479;
    n_n4114 <= n484;
    n_n3146 <= n489;
    n_n3511 <= n494;
    n_n3152 <= n499;
    n_n3833 <= n504;
    n_n4282 <= n509;
    n_n3305 <= n514;
    n_n4392 <= n519;
    n_n4224 <= n524;
    n_n3198 <= n529;
    n_n3204 <= n534;
    n_n3024 <= n539;
    n_n4139 <= n544;
    ndn3_15 <= n549;
    n_n3133 <= n554;
    n_n4074 <= n559;
    n_n3270 <= n564;
    n_n3858 <= n569;
    n_n3456 <= n574;
    n_n3521 <= n579;
    n_n3081 <= n584;
    n_n4381 <= n589;
    n_n3670 <= n594;
    n_n4211 <= n599;
    n_n3493 <= n604;
    n_n3495 <= n609;
    n_n3916 <= n614;
    n_n3195 <= n619;
    n_n3525 <= n624;
    n_n3729 <= n629;
    n_n3876 <= n634;
    ndn3_5 <= n639;
    n_n3549 <= n644;
    n_n3489 <= n649;
    n_n3764 <= n654;
    n_n3281 <= n659;
    n_n3707 <= n664;
    n_n3517 <= n669;
    n_n4160 <= n674;
    n_n4222 <= n679;
    n_n3012 <= n684;
    n_n4071 <= n689;
    n_n3372 <= n694;
    n_n3344 <= n699;
    n_n3688 <= n704;
    n_n3079 <= n709;
    n_n3313 <= n714;
    n_n3411 <= n719;
    n_n3231 <= n724;
    n_n3396 <= n729;
    n_n3432 <= n734;
    n_n3606 <= n739;
    n_n3733 <= n744;
    n_n3556 <= n749;
    n_n4040 <= n754;
    n_n3120 <= n759;
    n_n3221 <= n764;
    n_n3173 <= n769;
    n_n3851 <= n774;
    n_n3113 <= n779;
    n_n3242 <= n784;
    n_n3118 <= n789;
    n_n3376 <= n794;
    n_n4089 <= n799;
    n_n3044 <= n804;
    n_n3627 <= n809;
    n_n3035 <= n814;
    n_n3111 <= n819;
    n_n3321 <= n824;
    n_n3443 <= n829;
    n_n3215 <= n834;
    ndn3_10 <= n839;
    n_n4172 <= n844;
    nlc1_2 <= n849;
    n_n3590 <= n854;
    n_n4110 <= n859;
    nlc3_3 <= n864;
    n_n3576 <= n869;
    n_n4129 <= n874;
    n_n4189 <= n879;
    n_n4286 <= n884;
    n_n4383 <= n889;
    pdn <= n894;
    n_n3567 <= n898;
    n_n3892 <= n903;
    n_n3075 <= n908;
    n_n3354 <= n913;
    n_n3465 <= n918;
    ndn3_6 <= n923;
    n_n3617 <= n928;
    n_n4162 <= n933;
    n_n3207 <= n938;
    n_n4120 <= n943;
    n_n3065 <= n948;
    n_n4005 <= n953;
    n_n3266 <= n958;
    n_n4337 <= n963;
    n_n3600 <= n968;
    n_n3415 <= n973;
    n_n4243 <= n978;
    n_n3872 <= n983;
    n_n3648 <= n988;
    n_n3358 <= n993;
    n_n3350 <= n998;
    ndn3_7 <= n1003;
    n_n3116 <= n1008;
    n_n3583 <= n1013;
    n_n3906 <= n1018;
    n_n4131 <= n1023;
    n_n3316 <= n1028;
    n_n3061 <= n1033;
    n_n3048 <= n1038;
    n_n3886 <= n1043;
    n_n3919 <= n1048;
    n_n3128 <= n1053;
    n_n3995 <= n1058;
    n_n4213 <= n1063;
    n_n3761 <= n1068;
    ndn3_8 <= n1073;
    n_n3252 <= n1078;
    n_n4366 <= n1083;
    n_n3328 <= n1088;
    n_n3988 <= n1093;
    n_n3348 <= n1098;
    n_n3544 <= n1103;
    n_n3101 <= n1108;
    n_n4279 <= n1113;
    n_n3896 <= n1118;
    n_n3736 <= n1123;
    n_n4251 <= n1128;
    n_n3650 <= n1133;
    n_n3307 <= n1138;
    n_n4294 <= n1143;
    n_n4334 <= n1148;
    n_n3955 <= n1153;
    n_n4164 <= n1158;
    n_n3155 <= n1163;
    n_n3749 <= n1168;
    n_n4233 <= n1173;
    n_n4347 <= n1178;
    n_n3826 <= n1183;
    n_n3360 <= n1188;
    n_n3458 <= n1193;
    n_n3093 <= n1198;
    n_n3157 <= n1203;
    n_n3506 <= n1208;
    n_n3161 <= n1213;
    n_n3319 <= n1218;
    n_n3429 <= n1223;
    n_n3971 <= n1228;
    n_n3449 <= n1233;
    n_n4270 <= n1238;
    n_n4288 <= n1243;
    n_n3183 <= n1248;
    n_n3130 <= n1253;
    nlak4_2 <= n1258;
    n_n4047 <= n1263;
    n_n3978 <= n1268;
    n_n3239 <= n1273;
    n_n4145 <= n1278;
    n_n3890 <= n1283;
    n_n4003 <= n1288;
    n_n3091 <= n1293;
    n_n3985 <= n1298;
    n_n3326 <= n1303;
    n_n4052 <= n1308;
    nsr4_2 <= n1313;
    n_n4099 <= n1318;
    n_n4375 <= n1323;
    n_n4067 <= n1328;
    n_n4290 <= n1333;
    n_n3898 <= n1338;
    n_n4122 <= n1343;
    n_n3774 <= n1348;
    n_n3014 <= n1353;
    n_n4241 <= n1358;
    n_n3952 <= n1363;
    n_n3237 <= n1368;
    n_n3968 <= n1373;
    n_n3922 <= n1378;
    n_n3551 <= n1383;
    n_n3379 <= n1388;
    n_n4275 <= n1393;
    n_n3570 <= n1398;
    n_n3854 <= n1403;
    n_n4057 <= n1408;
    n_n3451 <= n1413;
    n_n4037 <= n1418;
    n_n3408 <= n1423;
    n_n4229 <= n1428;
    n_n4201 <= n1433;
    n_n3339 <= n1438;
    n_n4362 <= n1443;
    n_n3483 <= n1448;
    n_n3557 <= n1453;
    n_n4185 <= n1458;
    n_n3069 <= n1463;
    n_n3643 <= n1468;
    n_n3404 <= n1473;
    n_n3057 <= n1478;
    n_n3020 <= n1483;
    n_n3828 <= n1488;
    n_n3631 <= n1493;
    n_n3138 <= n1498;
    nsr1_2 <= n1503;
    n_n4065 <= n1508;
    n_n3679 <= n1513;
    n_n3287 <= n1518;
    n_n4351 <= n1523;
    n_n4059 <= n1528;
    n_n3436 <= n1533;
    nen3_10 <= n1538;
    n_n3461 <= n1543;
    n_n4012 <= n1548;
    n_n3051 <= n1553;
    n_n3073 <= n1558;
    n_n3777 <= n1563;
    n_n3709 <= n1568;
    n_n3946 <= n1573;
    n_n3085 <= n1578;
    n_n3259 <= n1583;
    n_n3504 <= n1588;
    n_n4045 <= n1593;
    n_n3954 <= n1598;
    n_n3136 <= n1603;
    n_n4372 <= n1608;
    n_n4236 <= n1613;
    n_n3040 <= n1618;
    n_n3874 <= n1623;
    n_n3999 <= n1628;
    n_n3223 <= n1633;
    ndn1_34 <= n1638;
    n_n3743 <= n1643;
    n_n3657 <= n1648;
    n_n3213 <= n1653;
    n_n3095 <= n1658;
    n_n3663 <= n1663;
    n_n3724 <= n1668;
    n_n3038 <= n1673;
    n_n3370 <= n1678;
    n_n3624 <= n1683;
    n_n3578 <= n1688;
    n_n3713 <= n1693;
    n_n3089 <= n1698;
    n_n3211 <= n1703;
    n_n3367 <= n1708;
    n_n3434 <= n1713;
    n_n3126 <= n1718;
    n_n4192 <= n1723;
    n_n4136 <= n1728;
    n_n3053 <= n1733;
    n_n3938 <= n1738;
    n_n3769 <= n1743;
    n_n4390 <= n1748;
    nsr3_17 <= n1753;
    n_n3903 <= n1758;
    n_n3658 <= n1763;
    nrq3_11 <= n1768;
    n_n3818 <= n1773;
    n_n3533 <= n1778;
    n_n3463 <= n1783;
    n_n3175 <= n1788;
    n_n3055 <= n1793;
    n_n3202 <= n1798;
    n_n3385 <= n1803;
    n_n4077 <= n1808;
    n_n3142 <= n1813;
    n_n3901 <= n1818;
    n_n3934 <= n1823;
    n_n3823 <= n1828;
    n_n3722 <= n1833;
    n_n4309 <= n1838;
    n_n4159 <= n1843;
    n_n4330 <= n1848;
    n_n3836 <= n1853;
    n_n3470 <= n1858;
    n_n3331 <= n1863;
    n_n3883 <= n1868;
    n_n4299 <= n1873;
    n_n4157 <= n1878;
    ndn3_9 <= n1883;
    n_n3208 <= n1888;
    n_n3190 <= n1893;
    n_n4029 <= n1898;
    n_n3042 <= n1903;
    nsr3_14 <= n1908;
    n_n4151 <= n1913;
    n_n3188 <= n1918;
    n_n4303 <= n1923;
    n_n3250 <= n1928;
    n_n3170 <= n1933;
    n_n3758 <= n1938;
    n_n3910 <= n1943;
    n_n3108 <= n1948;
    n_n3150 <= n1953;
    n_n4320 <= n1958;
    n_n4360 <= n1963;
    n_n4247 <= n1968;
    n_n4199 <= n1973;
    n_n3966 <= n1978;
    n_n3766 <= n1983;
    n_n4021 <= n1988;
    n_n4062 <= n1993;
    n_n3514 <= n1998;
    n_n3572 <= n2003;
    n_n4166 <= n2008;
    n_n3976 <= n2013;
    n_n3394 <= n2018;
    n_n4095 <= n2023;
    n_n3863 <= n2028;
    n_n3720 <= n2033;
    ngfdn_3 <= n2038;
    n_n3756 <= n2043;
    n_n3667 <= n2048;
    n_n3342 <= n2053;
    n_n3529 <= n2058;
    n_n4209 <= n2063;
    n_n4324 <= n2068;
    n_n3337 <= n2073;
    n_n4227 <= n2078;
    n_n4153 <= n2083;
    n_n3831 <= n2088;
    n_n3233 <= n2093;
    n_n4263 <= n2098;
    n_n3413 <= n2103;
    n_n4182 <= n2108;
    n_n3841 <= n2113;
    n_n3441 <= n2118;
    n_n4026 <= n2123;
    n_n4342 <= n2128;
    n_n4102 <= n2133;
    n_n3277 <= n2138;
    n_n4180 <= n2143;
    n_n3878 <= n2148;
    n_n3931 <= n2153;
    n_n3845 <= n2158;
    n_n3865 <= n2163;
    n_n3486 <= n2168;
    n_n4056 <= n2173;
    n_n3674 <= n2178;
    n_n3959 <= n2183;
    n_n3608 <= n2188;
    n_n4080 <= n2193;
    n_n4018 <= n2198;
    n_n4354 <= n2203;
    n_n3797 <= n2208;
    n_n3739 <= n2213;
    n_n3646 <= n2218;
    n_n3099 <= n2223;
    n_n3537 <= n2228;
    n_n3806 <= n2233;
    n_n3087 <= n2238;
    n_n4105 <= n2243;
    n_n3262 <= n2248;
    n_n4125 <= n2253;
    n_n3814 <= n2258;
    n_n4093 <= n2263;
    nsr3_3 <= n2268;
  end
endmodule


