// Benchmark "top" written by ABC on Tue Mar  5 10:01:57 2019

module dsip ( clk, 
    pcount_3_, pkey_5_, pkey_131_, pkey_144_, pkey_157_, pkey_230_,
    pkey_243_, pcount_2_, pkey_4_, pkey_132_, pkey_158_, pkey_169_,
    pkey_242_, pcount_1_, pkey_146_, pkey_168_, pkey_245_, pcount_0_,
    pkey_6_, pkey_130_, pkey_145_, pkey_244_, pkey_9_, pkey_16_, pkey_27_,
    pkey_38_, pkey_49_, pkey_122_, pkey_148_, pkey_153_, pkey_166_,
    pkey_221_, pkey_252_, pkey_8_, pkey_17_, pkey_26_, pkey_48_, pkey_110_,
    pkey_121_, pkey_147_, pkey_154_, pkey_165_, pkey_220_, pkey_246_,
    pkey_253_, pkey_18_, pkey_29_, pkey_36_, pkey_120_, pkey_155_,
    pkey_164_, pkey_210_, pkey_249_, pkey_254_, pkey_19_, pkey_28_,
    pkey_37_, pkey_46_, pkey_112_, pkey_149_, pkey_156_, pkey_163_,
    pkey_211_, pkey_248_, pkey_56_, pkey_67_, pkey_78_, pkey_89_,
    pkey_113_, pkey_126_, pkey_139_, pkey_162_, pkey_212_, pkey_225_,
    pkey_238_, pkey_57_, pkey_66_, pkey_88_, pkey_114_, pkey_125_,
    pkey_150_, pkey_161_, pkey_213_, pkey_224_, pkey_58_, pkey_69_,
    pkey_76_, pkey_115_, pkey_124_, pkey_137_, pkey_160_, pkey_214_,
    pkey_250_, pkey_59_, pkey_68_, pkey_77_, pkey_86_, pkey_116_,
    pkey_123_, pkey_138_, pkey_152_, pkey_222_, pkey_237_, pkey_251_,
    pkey_1_, pkey_96_, pkey_117_, pkey_140_, pkey_216_, pkey_229_,
    pkey_234_, pkey_0_, pkey_97_, pkey_118_, pkey_129_, pkey_136_,
    pkey_217_, pkey_228_, pkey_235_, pkey_3_, pkey_98_, pkey_128_,
    pkey_133_, pkey_142_, pkey_218_, pkey_227_, pkey_232_, pkey_241_,
    pkey_2_, pkey_99_, pkey_134_, pkey_141_, pkey_219_, pkey_226_,
    pkey_233_, pkey_240_, pkey_70_, pkey_81_, pkey_92_, pkey_180_,
    pkey_193_, pkey_80_, pkey_93_, pkey_107_, pkey_194_, pkey_206_, 
    pkey_50_, pkey_61_, pkey_94_, pkey_182_, pkey_195_, pkey_209_,
    pstart_0_, pkey_51_, pkey_60_, pkey_109_, pkey_181_, pkey_196_,
    pkey_208_, pkey_52_, pkey_74_, pkey_85_, pkey_104_, pkey_171_,
    pkey_197_, pkey_203_, pencrypt_0_, pkey_53_, pkey_62_, pkey_75_,
    pkey_84_, pkey_172_, pkey_198_, pkey_202_, pkey_54_, pkey_65_,
    pkey_72_, pkey_83_, pkey_90_, pkey_106_, pkey_205_, pkey_64_, pkey_73_,
    pkey_82_, pkey_91_, pkey_105_, pkey_170_, pkey_204_, pkey_12_,
    pkey_34_, pkey_45_, pkey_100_, pkey_188_, pkey_13_, pkey_22_, pkey_35_,
    pkey_44_, pkey_176_, pkey_187_, pkey_14_, pkey_25_, pkey_32_, pkey_43_,
    pkey_102_, pkey_173_, pkey_201_, pkey_24_, pkey_33_, pkey_42_,
    pkey_101_, pkey_174_, pkey_189_, pkey_200_, pkey_30_, pkey_41_,
    pkey_179_, pkey_184_, pkey_40_, pkey_190_, pkey_10_, pkey_21_,
    pkey_177_, pkey_186_, pkey_11_, pkey_20_, pkey_178_, pkey_185_,
    pkey_192_,
    pksi_50_, pksi_61_, pksi_72_, pksi_83_, pksi_94_, pksi_102_, pksi_115_,
    pksi_128_, pdata_ready_0_, pksi_51_, pksi_60_, pksi_73_, pksi_82_,
    pksi_95_, pksi_101_, pksi_116_, pksi_127_, pksi_52_, pksi_63_,
    pksi_70_, pksi_81_, pksi_96_, pksi_100_, pksi_113_, pksi_53_, pksi_62_,
    pksi_71_, pksi_80_, pksi_97_, pksi_114_, pksi_129_, pksi_54_, pksi_65_,
    pksi_76_, pksi_87_, pksi_90_, pksi_119_, pksi_124_, pksi_191_,
    pksi_55_, pksi_64_, pksi_77_, pksi_86_, pksi_91_, pksi_123_, pksi_56_,
    pksi_67_, pksi_74_, pksi_85_, pksi_92_, pksi_117_, pksi_126_, pksi_57_,
    pksi_66_, pksi_75_, pksi_84_, pksi_93_, pksi_118_, pksi_125_,
    pksi_190_, pksi_14_, pksi_25_, pksi_36_, pksi_47_, pksi_120_, pksi_15_,
    pksi_24_, pksi_37_, pksi_46_, pksi_109_, pnew_count_3_, pksi_16_,
    pksi_27_, pksi_34_, pksi_45_, pksi_108_, pksi_122_, pksi_17_, pksi_26_,
    pksi_35_, pksi_44_, pksi_107_, pksi_121_, pksi_10_, pksi_21_, pksi_32_,
    pksi_43_, pksi_106_, pksi_111_, pnew_count_0_, pksi_11_, pksi_20_,
    pksi_33_, pksi_42_, pksi_105_, pksi_112_, pksi_12_, pksi_23_, pksi_30_,
    pksi_41_, pksi_104_, pnew_count_2_, pksi_13_, pksi_22_, pksi_31_,
    pksi_40_, pksi_103_, pksi_110_, pnew_count_1_, pksi_3_, pksi_151_,
    pksi_164_, pksi_177_, pksi_2_, pksi_152_, pksi_163_, pksi_178_,
    pksi_189_, pksi_1_, pksi_166_, pksi_179_, pksi_188_, pksi_0_,
    pksi_150_, pksi_165_, pksi_187_, pksi_18_, pksi_29_, pksi_142_,
    pksi_168_, pksi_173_, pksi_186_, pksi_19_, pksi_28_, pksi_130_,
    pksi_141_, pksi_167_, pksi_174_, pksi_185_, pksi_38_, pksi_49_,
    pksi_131_, pksi_140_, pksi_175_, pksi_184_, pksi_39_, pksi_48_,
    pksi_132_, pksi_169_, pksi_176_, pksi_183_, pksi_58_, pksi_69_,
    pksi_133_, pksi_146_, pksi_159_, pksi_182_, pksi_59_, pksi_68_,
    pksi_134_, pksi_145_, pksi_170_, pksi_181_, pksi_9_, pksi_78_,
    pksi_89_, pksi_135_, pksi_144_, pksi_157_, pksi_171_, pksi_180_,
    pksi_8_, pksi_79_, pksi_88_, pksi_136_, pksi_143_, pksi_158_,
    pksi_172_, pksi_7_, pksi_98_, pksi_137_, pksi_155_, pksi_160_, pksi_6_,
    pksi_99_, pksi_138_, pksi_149_, pksi_156_, pksi_5_, pksi_139_,
    pksi_148_, pksi_153_, pksi_162_, pksi_4_, pksi_147_, pksi_154_,
    pksi_161_  );
  input  pcount_3_, pkey_5_, pkey_131_, pkey_144_, pkey_157_, pkey_230_,
    pkey_243_, pcount_2_, pkey_4_, pkey_132_, pkey_158_, pkey_169_,
    pkey_242_, pcount_1_, pkey_146_, pkey_168_, pkey_245_, pcount_0_,
    pkey_6_, pkey_130_, pkey_145_, pkey_244_, pkey_9_, pkey_16_, pkey_27_,
    pkey_38_, pkey_49_, pkey_122_, pkey_148_, pkey_153_, pkey_166_,
    pkey_221_, pkey_252_, pkey_8_, pkey_17_, pkey_26_, pkey_48_, pkey_110_,
    pkey_121_, pkey_147_, pkey_154_, pkey_165_, pkey_220_, pkey_246_,
    pkey_253_, pkey_18_, pkey_29_, pkey_36_, pkey_120_, pkey_155_,
    pkey_164_, pkey_210_, pkey_249_, pkey_254_, pkey_19_, pkey_28_,
    pkey_37_, pkey_46_, pkey_112_, pkey_149_, pkey_156_, pkey_163_,
    pkey_211_, pkey_248_, pkey_56_, pkey_67_, pkey_78_, pkey_89_,
    pkey_113_, pkey_126_, pkey_139_, pkey_162_, pkey_212_, pkey_225_,
    pkey_238_, pkey_57_, pkey_66_, pkey_88_, pkey_114_, pkey_125_,
    pkey_150_, pkey_161_, pkey_213_, pkey_224_, pkey_58_, pkey_69_,
    pkey_76_, pkey_115_, pkey_124_, pkey_137_, pkey_160_, pkey_214_,
    pkey_250_, pkey_59_, pkey_68_, pkey_77_, pkey_86_, pkey_116_,
    pkey_123_, pkey_138_, pkey_152_, pkey_222_, pkey_237_, pkey_251_,
    pkey_1_, pkey_96_, pkey_117_, pkey_140_, pkey_216_, pkey_229_,
    pkey_234_, pkey_0_, pkey_97_, pkey_118_, pkey_129_, pkey_136_,
    pkey_217_, pkey_228_, pkey_235_, pkey_3_, pkey_98_, pkey_128_,
    pkey_133_, pkey_142_, pkey_218_, pkey_227_, pkey_232_, pkey_241_,
    pkey_2_, pkey_99_, pkey_134_, pkey_141_, pkey_219_, pkey_226_,
    pkey_233_, pkey_240_, pkey_70_, pkey_81_, pkey_92_, pkey_180_,
    pkey_193_, pkey_80_, pkey_93_, pkey_107_, pkey_194_, pkey_206_, clk,
    pkey_50_, pkey_61_, pkey_94_, pkey_182_, pkey_195_, pkey_209_,
    pstart_0_, pkey_51_, pkey_60_, pkey_109_, pkey_181_, pkey_196_,
    pkey_208_, pkey_52_, pkey_74_, pkey_85_, pkey_104_, pkey_171_,
    pkey_197_, pkey_203_, pencrypt_0_, pkey_53_, pkey_62_, pkey_75_,
    pkey_84_, pkey_172_, pkey_198_, pkey_202_, pkey_54_, pkey_65_,
    pkey_72_, pkey_83_, pkey_90_, pkey_106_, pkey_205_, pkey_64_, pkey_73_,
    pkey_82_, pkey_91_, pkey_105_, pkey_170_, pkey_204_, pkey_12_,
    pkey_34_, pkey_45_, pkey_100_, pkey_188_, pkey_13_, pkey_22_, pkey_35_,
    pkey_44_, pkey_176_, pkey_187_, pkey_14_, pkey_25_, pkey_32_, pkey_43_,
    pkey_102_, pkey_173_, pkey_201_, pkey_24_, pkey_33_, pkey_42_,
    pkey_101_, pkey_174_, pkey_189_, pkey_200_, pkey_30_, pkey_41_,
    pkey_179_, pkey_184_, pkey_40_, pkey_190_, pkey_10_, pkey_21_,
    pkey_177_, pkey_186_, pkey_11_, pkey_20_, pkey_178_, pkey_185_,
    pkey_192_;
  output pksi_50_, pksi_61_, pksi_72_, pksi_83_, pksi_94_, pksi_102_,
    pksi_115_, pksi_128_, pdata_ready_0_, pksi_51_, pksi_60_, pksi_73_,
    pksi_82_, pksi_95_, pksi_101_, pksi_116_, pksi_127_, pksi_52_,
    pksi_63_, pksi_70_, pksi_81_, pksi_96_, pksi_100_, pksi_113_, pksi_53_,
    pksi_62_, pksi_71_, pksi_80_, pksi_97_, pksi_114_, pksi_129_, pksi_54_,
    pksi_65_, pksi_76_, pksi_87_, pksi_90_, pksi_119_, pksi_124_,
    pksi_191_, pksi_55_, pksi_64_, pksi_77_, pksi_86_, pksi_91_, pksi_123_,
    pksi_56_, pksi_67_, pksi_74_, pksi_85_, pksi_92_, pksi_117_, pksi_126_,
    pksi_57_, pksi_66_, pksi_75_, pksi_84_, pksi_93_, pksi_118_, pksi_125_,
    pksi_190_, pksi_14_, pksi_25_, pksi_36_, pksi_47_, pksi_120_, pksi_15_,
    pksi_24_, pksi_37_, pksi_46_, pksi_109_, pnew_count_3_, pksi_16_,
    pksi_27_, pksi_34_, pksi_45_, pksi_108_, pksi_122_, pksi_17_, pksi_26_,
    pksi_35_, pksi_44_, pksi_107_, pksi_121_, pksi_10_, pksi_21_, pksi_32_,
    pksi_43_, pksi_106_, pksi_111_, pnew_count_0_, pksi_11_, pksi_20_,
    pksi_33_, pksi_42_, pksi_105_, pksi_112_, pksi_12_, pksi_23_, pksi_30_,
    pksi_41_, pksi_104_, pnew_count_2_, pksi_13_, pksi_22_, pksi_31_,
    pksi_40_, pksi_103_, pksi_110_, pnew_count_1_, pksi_3_, pksi_151_,
    pksi_164_, pksi_177_, pksi_2_, pksi_152_, pksi_163_, pksi_178_,
    pksi_189_, pksi_1_, pksi_166_, pksi_179_, pksi_188_, pksi_0_,
    pksi_150_, pksi_165_, pksi_187_, pksi_18_, pksi_29_, pksi_142_,
    pksi_168_, pksi_173_, pksi_186_, pksi_19_, pksi_28_, pksi_130_,
    pksi_141_, pksi_167_, pksi_174_, pksi_185_, pksi_38_, pksi_49_,
    pksi_131_, pksi_140_, pksi_175_, pksi_184_, pksi_39_, pksi_48_,
    pksi_132_, pksi_169_, pksi_176_, pksi_183_, pksi_58_, pksi_69_,
    pksi_133_, pksi_146_, pksi_159_, pksi_182_, pksi_59_, pksi_68_,
    pksi_134_, pksi_145_, pksi_170_, pksi_181_, pksi_9_, pksi_78_,
    pksi_89_, pksi_135_, pksi_144_, pksi_157_, pksi_171_, pksi_180_,
    pksi_8_, pksi_79_, pksi_88_, pksi_136_, pksi_143_, pksi_158_,
    pksi_172_, pksi_7_, pksi_98_, pksi_137_, pksi_155_, pksi_160_, pksi_6_,
    pksi_99_, pksi_138_, pksi_149_, pksi_156_, pksi_5_, pksi_139_,
    pksi_148_, pksi_153_, pksi_162_, pksi_4_, pksi_147_, pksi_154_,
    pksi_161_;
  reg pksi_17_, pksi_185_, n_n2410, pksi_170_, pksi_155_, pksi_147_,
    pksi_109_, n_n2513, pksi_19_, n_n2396, n_n2412, n_n121, pksi_148_,
    n_n2448, pksi_107_, pksi_110_, pksi_9_, pksi_176_, pksi_180_,
    pksi_178_, pksi_135_, pksi_129_, pksi_100_, pksi_117_, pksi_118_,
    pksi_5_, pksi_169_, n_n2408, pksi_184_, pksi_125_, pksi_138_,
    pksi_114_, pksi_99_, pksi_85_, pksi_14_, pksi_4_, pksi_186_, n_n2420,
    pksi_141_, pksi_113_, pksi_115_, pksi_98_, pksi_2_, pksi_23_,
    pksi_177_, pksi_189_, n_n2485, n_n2495, pksi_97_, pksi_102_, pksi_11_,
    pksi_173_, pksi_179_, pksi_171_, pksi_104_, pksi_103_, n_n2384,
    pksi_183_, pksi_172_, n_n2416, pksi_116_, pksi_96_, pksi_119_,
    pksi_84_, pksi_159_, n_n2440, pksi_160_, pksi_128_, pksi_127_,
    pksi_142_, n_n2272, pksi_149_, pksi_162_, pksi_154_, pksi_121_,
    pksi_134_, pksi_126_, pksi_82_, n_n2430, pksi_153_, pksi_165_,
    pksi_137_, n_n2481, pksi_101_, pksi_93_, pksi_161_, pksi_156_, n_n2452,
    n_n2462, pksi_123_, pksi_111_, pksi_92_, pksi_15_, n_n109, pksi_145_,
    pksi_144_, pksi_150_, pksi_124_, pksi_132_, pksi_130_, pksi_105_,
    pksi_112_, n_n10, pksi_6_, pksi_188_, pksi_152_, pksi_163_, pksi_166_,
    pksi_131_, n_n2474, pksi_136_, pksi_108_, n_n2517, n_n2268, pksi_175_,
    pksi_190_, pksi_164_, pksi_158_, pksi_167_, pksi_133_, n_n2476,
    pksi_122_, n_n2507, pksi_75_, pksi_182_, pksi_174_, pksi_157_,
    pksi_151_, pksi_146_, pksi_140_, pksi_120_, n_n168, pksi_106_,
    pksi_57_, pksi_36_, pksi_38_, pksi_28_, n_n2374, pksi_53_, pksi_27_,
    pksi_26_, pksi_47_, pksi_1_, pksi_63_, pksi_34_, pksi_24_, pksi_30_,
    pksi_18_, pksi_79_, pksi_54_, n_n2337, pksi_46_, pksi_39_, pksi_8_,
    n_n2277, pksi_91_, pksi_51_, pksi_70_, pksi_0_, pksi_73_, pksi_89_,
    pksi_60_, pksi_48_, pksi_22_, n_n2280, pksi_77_, pksi_64_, pksi_56_,
    pksi_80_, pksi_81_, n_n2301, pksi_66_, pksi_72_, pksi_78_, pksi_69_,
    n_n2320, pksi_40_, pksi_32_, pksi_94_, pksi_87_, pksi_61_, pksi_59_,
    n_n2333, pksi_42_, pksi_86_, pksi_76_, n_n2305, pksi_50_, pksi_33_,
    pksi_12_, pksi_74_, pksi_95_, pksi_58_, pksi_62_, pksi_29_, pksi_3_,
    pksi_83_, pksi_68_, pksi_71_, pksi_37_, pksi_41_, n_n2365, n_n2369,
    n_n2288, pksi_55_, pksi_52_, pksi_45_, pksi_43_, pksi_16_, pksi_10_,
    n_n2310, pksi_67_, pksi_31_, pksi_25_, pksi_35_, pksi_20_, pksi_21_,
    pksi_49_, pksi_65_, pksi_44_, n_n2342, n_n2352, pksi_7_, pksi_13_;
  wire n1327_1, n1328, n1329, n1330, n1331, n1332_1, n1341, n1342, n1343,
    n1344_1, n1345, n1346, n1347, n1348_1, n1349, n1350, n1351, n1352_1,
    n1353, n1354, n1355, n1356_1, n1357, n1358, n1359, n1360, n1361_1,
    n1362, n1363, n1364, n1365_1, n1366, n1367, n1368, n1369, n1370_1,
    n1371, n1372, n1373, n1374_1, n1375, n1376, n1377, n1378_1, n1379,
    n1380, n1381, n1382_1, n1383, n1384, n1385, n1386_1, n1387, n1388,
    n1389, n1390_1, n1391, n1392, n1393, n1394_1, n1395, n1396, n1397,
    n1398_1, n1399, n1400, n1401, n1402_1, n1403, n1404, n1405, n1406,
    n1407_1, n1408, n1409, n1410, n1411_1, n1412, n1413, n1414, n1415_1,
    n1416, n1417, n1418, n1419_1, n1420, n1421, n1422, n1423_1, n1424,
    n1425, n1426, n1427_1, n1428, n1429, n1430, n1431, n1432_1, n1433,
    n1434, n1435, n1436_1, n1437, n1438, n1439, n1440_1, n1441, n1442,
    n1443, n1444_1, n1445, n1446, n1447, n1448_1, n1449, n1450, n1451,
    n1452_1, n1453, n1454, n1455, n1456_1, n1457, n1458, n1459, n1460_1,
    n1461, n1462, n1463, n1464_1, n1465, n1466, n1467, n1468_1, n1469,
    n1470, n1471, n1472_1, n1473, n1474, n1475, n1476_1, n1477, n1478,
    n1479, n1480_1, n1481, n1482, n1483, n1484, n1485_1, n1486, n1487,
    n1488, n1489_1, n1490, n1491, n1492, n1493_1, n1494, n1495, n1496,
    n1497_1, n1498, n1499, n1500, n1501, n1502_1, n1503, n1504, n1505,
    n1506_1, n1507, n1508, n1509, n1510_1, n1511, n1512, n1513, n1514_1,
    n1515, n1516, n1517, n1518_1, n1519, n1520, n1521, n1522_1, n1523,
    n1524, n1525, n1526_1, n1527, n1528, n1529, n1530_1, n1531, n1532,
    n1533, n1534_1, n1535, n1536, n1537, n1538_1, n1539, n1540, n1541,
    n1542, n1543_1, n1544, n1545, n1546, n1547_1, n1548, n1549, n1550,
    n1551_1, n1552, n1553, n1554, n1555_1, n1556, n1557, n1558, n1559_1,
    n1560, n1561, n1562, n1563_1, n1564, n1565, n1566, n1567, n1568_1,
    n1569, n1570, n1571, n1572_1, n1573, n1574, n1575, n1576_1, n1577,
    n1578, n1579, n1580_1, n1581, n1582, n1583, n1584_1, n1585, n1586,
    n1587, n1588, n1589_1, n1590, n1591, n1592, n1593_1, n1594, n1595,
    n1596, n1597_1, n1598, n1599, n1600, n1601_1, n1602, n1603, n1604,
    n1605_1, n1606, n1607, n1608, n1609_1, n1610, n1611, n1612, n1613_1,
    n1614, n1615, n1616, n1617, n1618_1, n1619, n1620, n1621, n1622_1,
    n1623, n1624, n1625, n1626_1, n1627, n1628, n1629, n1630_1, n1631,
    n1632, n1633, n1634, n1635_1, n1636, n1637, n1638, n1639_1, n1640,
    n1641, n1642, n1643_1, n1644, n1645, n1646, n1647_1, n1648, n1649,
    n1650, n1651_1, n1652, n1653, n1654, n1655_1, n1656, n1657, n1658,
    n1659_1, n1660, n1661, n1662, n1663_1, n1664, n1665, n1666, n1667_1,
    n1668, n1669, n1670, n1671_1, n1672, n1673, n1674, n1675_1, n1676,
    n1677, n1678, n1679_1, n1680, n1681, n1682, n1683_1, n1684, n1685,
    n1686, n1687_1, n1688, n1689, n1690, n1691_1, n1692, n1693, n1694,
    n1695, n1696_1, n1697, n1698, n1699, n1700, n1701_1, n1702, n1703,
    n1704, n1705, n1706_1, n1707, n1708, n1709, n1710_1, n1711, n1712,
    n1713, n1714_1, n1715, n1716, n1717, n1718_1, n1719, n1720, n1721,
    n1722_1, n1723, n1724, n1725, n1726_1, n1727, n1728, n1729, n1730_1,
    n1731, n1732, n1733, n1734, n1735_1, n1736, n1737, n1738, n1739_1,
    n1740, n1741, n1742, n1743_1, n1744, n1745, n1746, n1747_1, n1748,
    n1749, n1750, n1751_1, n1752, n1753, n1754, n1755_1, n1756, n1757,
    n1758, n1759_1, n1760, n1761, n1762, n1763_1, n1764, n1765, n1766,
    n1767_1, n1768, n1769, n1770, n1771_1, n1772, n1773, n1774, n1775,
    n1776_1, n1777, n1778, n1779, n1780, n1781_1, n1782, n1783, n1784,
    n1785_1, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
    n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
    n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
    n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
    n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
    n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
    n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
    n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
    n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
    n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
    n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
    n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
    n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
    n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
    n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
    n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
    n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
    n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
    n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
    n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
    n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
    n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
    n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
    n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
    n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
    n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
    n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
    n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
    n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
    n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
    n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
    n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
    n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
    n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
    n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
    n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
    n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
    n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
    n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
    n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
    n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
    n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
    n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
    n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
    n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
    n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
    n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
    n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
    n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
    n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
    n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
    n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
    n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
    n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
    n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
    n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
    n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
    n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
    n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
    n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
    n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
    n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
    n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
    n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
    n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
    n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
    n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
    n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
    n2465, n2466, n2467, n853, n857, n861, n866, n870, n874, n878, n882,
    n887, n891, n896, n901, n906, n910, n915, n919, n923, n927, n931, n935,
    n939, n943, n947, n951, n955, n959, n963, n967, n972, n976, n980, n984,
    n988, n992, n996, n1000, n1004, n1008, n1013, n1017, n1021, n1025,
    n1029, n1033, n1037, n1041, n1045, n1050, n1055, n1059, n1063, n1067,
    n1071, n1075, n1079, n1083, n1087, n1092, n1096, n1100, n1105, n1109,
    n1113, n1117, n1121, n1125, n1130, n1134, n1138, n1142, n1146, n1151,
    n1155, n1159, n1163, n1167, n1171, n1175, n1179, n1184, n1188, n1192,
    n1196, n1201, n1205, n1209, n1213, n1217, n1222, n1227, n1231, n1235,
    n1239, n1243, n1248, n1252, n1256, n1260, n1264, n1268, n1272, n1276,
    n1280, n1285, n1289, n1293, n1297, n1301, n1305, n1309, n1314, n1318,
    n1322, n1327, n1332, n1336, n1340, n1344, n1348, n1352, n1356, n1361,
    n1365, n1370, n1374, n1378, n1382, n1386, n1390, n1394, n1398, n1402,
    n1407, n1411, n1415, n1419, n1423, n1427, n1432, n1436, n1440, n1444,
    n1448, n1452, n1456, n1460, n1464, n1468, n1472, n1476, n1480, n1485,
    n1489, n1493, n1497, n1502, n1506, n1510, n1514, n1518, n1522, n1526,
    n1530, n1534, n1538, n1543, n1547, n1551, n1555, n1559, n1563, n1568,
    n1572, n1576, n1580, n1584, n1589, n1593, n1597, n1601, n1605, n1609,
    n1613, n1618, n1622, n1626, n1630, n1635, n1639, n1643, n1647, n1651,
    n1655, n1659, n1663, n1667, n1671, n1675, n1679, n1683, n1687, n1691,
    n1696, n1701, n1706, n1710, n1714, n1718, n1722, n1726, n1730, n1735,
    n1739, n1743, n1747, n1751, n1755, n1759, n1763, n1767, n1771, n1776,
    n1781, n1785;
  assign pdata_ready_0_ = (n1327_1 & n2465) | (n1328 & n1329);
  assign pnew_count_3_ = n1343 | n1342 | (pstart_0_ & ~pencrypt_0_);
  assign pnew_count_0_ = pstart_0_ ? ~pencrypt_0_ : ~pcount_0_;
  assign pnew_count_2_ = n2467 | (pcount_2_ & ~n1331);
  assign pnew_count_1_ = (pcount_1_ & (pcount_0_ ? ~pencrypt_0_ : (~pstart_0_ & pencrypt_0_))) | (~pcount_1_ & (pcount_0_ ? (~pstart_0_ & pencrypt_0_) : ~pencrypt_0_)) | (pstart_0_ & ~pencrypt_0_);
  assign n853 = n2014 | n2015 | n2016 | n2018;
  assign n857 = n2011 | n2012 | n2013 | n2020;
  assign n861 = n2008 | n2009 | n2010 | n2022;
  assign n866 = n2005 | n2006 | n2007 | n2024;
  assign n870 = n2002 | n2003 | n2004 | n2026;
  assign n874 = n1999 | n2000 | n2001 | n2028;
  assign n878 = n1996 | n1997 | n1998 | n2030;
  assign n882 = n1993 | n1994 | n1995 | n2032;
  assign n887 = n1990 | n1991 | n1992 | n2034;
  assign n891 = n1987 | n1988 | n1989 | n2036;
  assign n896 = n1984 | n1985 | n1986 | n2038;
  assign n901 = n1981 | n1982 | n1983 | n2040;
  assign n906 = n1978 | n1979 | n1980 | n2042;
  assign n910 = n1975 | n1976 | n1977 | n2044;
  assign n915 = n1972 | n1973 | n1974 | n2046;
  assign n919 = n1969 | n1970 | n1971 | n2048;
  assign n923 = n1966 | n1967 | n1968 | n2050;
  assign n927 = n1963 | n1964 | n1965 | n2052;
  assign n931 = n1960 | n1961 | n1962 | n2054;
  assign n935 = n1957 | n1958 | n1959 | n2056;
  assign n939 = n1954 | n1955 | n1956 | n2058;
  assign n943 = n1951 | n1952 | n1953 | n2060;
  assign n947 = n1948 | n1949 | n1950 | n2062;
  assign n951 = n1945 | n1946 | n1947 | n2064;
  assign n955 = n1942 | n1943 | n1944 | n2066;
  assign n959 = n1939 | n1940 | n1941 | n2068;
  assign n963 = n1936 | n1937 | n1938 | n2070;
  assign n967 = n1933 | n1934 | n1935 | n2072;
  assign n972 = n1930 | n1931 | n1932 | n2074;
  assign n976 = n1927 | n1928 | n1929 | n2076;
  assign n980 = n1924 | n1925 | n1926 | n2078;
  assign n984 = n1921 | n1922 | n1923 | n2080;
  assign n988 = n1918 | n1919 | n1920 | n2082;
  assign n992 = n1915 | n1916 | n1917 | n2084;
  assign n996 = n1912 | n1913 | n1914 | n2086;
  assign n1000 = n1909 | n1910 | n1911 | n2088;
  assign n1004 = n1906 | n1907 | n1908 | n2090;
  assign n1008 = n1903 | n1904 | n1905 | n2092;
  assign n1013 = n1900 | n1901 | n1902 | n2094;
  assign n1017 = n1897 | n1898 | n1899 | n2096;
  assign n1021 = n1894 | n1895 | n1896 | n2098;
  assign n1025 = n1891 | n1892 | n1893 | n2100;
  assign n1029 = n1888 | n1889 | n1890 | n2102;
  assign n1033 = n1885 | n1886 | n1887 | n2104;
  assign n1037 = n1882 | n1883 | n1884 | n2106;
  assign n1041 = n1879 | n1880 | n1881 | n2108;
  assign n1045 = n1876 | n1877 | n1878 | n2110;
  assign n1050 = n1873 | n1874 | n1875 | n2112;
  assign n1055 = n1870 | n1871 | n1872 | n2114;
  assign n1059 = n1867 | n1868 | n1869 | n2116;
  assign n1063 = n1864 | n1865 | n1866 | n2118;
  assign n1067 = n1861 | n1862 | n1863 | n2120;
  assign n1071 = n1858 | n1859 | n1860 | n2122;
  assign n1075 = n1855 | n1856 | n1857 | n2124;
  assign n1079 = n1852 | n1853 | n1854 | n2126;
  assign n1083 = n1849 | n1850 | n1851 | n2128;
  assign n1087 = n1846 | n1847 | n1848 | n2130;
  assign n1092 = n1843 | n1844 | n1845 | n2132;
  assign n1096 = n1840 | n1841 | n1842 | n2134;
  assign n1100 = n1837 | n1838 | n1839 | n2136;
  assign n1105 = n1834 | n1835 | n1836 | n2138;
  assign n1109 = n1831 | n1832 | n1833 | n2140;
  assign n1113 = n1828 | n1829 | n1830 | n2142;
  assign n1117 = n1825 | n1826 | n1827 | n2144;
  assign n1121 = n1822 | n1823 | n1824 | n2146;
  assign n1125 = n1819 | n1820 | n1821 | n2148;
  assign n1130 = n1816 | n1817 | n1818 | n2150;
  assign n1134 = n1813 | n1814 | n1815 | n2152;
  assign n1138 = n1810 | n1811 | n1812 | n2154;
  assign n1142 = n1807 | n1808 | n1809 | n2156;
  assign n1146 = n1804 | n1805 | n1806 | n2158;
  assign n1151 = n1801 | n1802 | n1803 | n2160;
  assign n1155 = n1798 | n1799 | n1800 | n2162;
  assign n1159 = n1795 | n1796 | n1797 | n2164;
  assign n1163 = n1792 | n1793 | n1794 | n2166;
  assign n1167 = n1789 | n1790 | n1791 | n2168;
  assign n1171 = n1786 | n1787 | n1788 | n2170;
  assign n1175 = n1783 | n1784 | n1785_1 | n2172;
  assign n1179 = n1780 | n1781_1 | n1782 | n2174;
  assign n1184 = n1777 | n1778 | n1779 | n2176;
  assign n1188 = n1774 | n1775 | n1776_1 | n2178;
  assign n1192 = n1771_1 | n1772 | n1773 | n2180;
  assign n1196 = n1768 | n1769 | n1770 | n2182;
  assign n1201 = n1765 | n1766 | n1767_1 | n2184;
  assign n1205 = n1762 | n1763_1 | n1764 | n2186;
  assign n1209 = n1759_1 | n1760 | n1761 | n2188;
  assign n1213 = n1756 | n1757 | n1758 | n2190;
  assign n1217 = n1753 | n1754 | n1755_1 | n2192;
  assign n1222 = n1750 | n1751_1 | n1752 | n2194;
  assign n1227 = n1747_1 | n1748 | n1749 | n2196;
  assign n1231 = n1744 | n1745 | n1746 | n2198;
  assign n1235 = n1741 | n1742 | n1743_1 | n2200;
  assign n1239 = n1738 | n1739_1 | n1740 | n2202;
  assign n1243 = n1735_1 | n1736 | n1737 | n2204;
  assign n1248 = n1732 | n1733 | n1734 | n2206;
  assign n1252 = n1729 | n1730_1 | n1731 | n2208;
  assign n1256 = n1726_1 | n1727 | n1728 | n2210;
  assign n1260 = n1723 | n1724 | n1725 | n2212;
  assign n1264 = n1720 | n1721 | n1722_1 | n2214;
  assign n1268 = n1717 | n1718_1 | n1719 | n2216;
  assign n1272 = n1714_1 | n1715 | n1716 | n2218;
  assign n1276 = n1711 | n1712 | n1713 | n2220;
  assign n1280 = n1708 | n1709 | n1710_1 | n2222;
  assign n1285 = n1705 | n1706_1 | n1707 | n2224;
  assign n1289 = n1702 | n1703 | n1704 | n2226;
  assign n1293 = n1699 | n1700 | n1701_1 | n2228;
  assign n1297 = n1696_1 | n1697 | n1698 | n2230;
  assign n1301 = n1693 | n1694 | n1695 | n2232;
  assign n1305 = n1690 | n1691_1 | n1692 | n2234;
  assign n1309 = n1687_1 | n1688 | n1689 | n2236;
  assign n1314 = n1684 | n1685 | n1686 | n2238;
  assign n1318 = n1681 | n1682 | n1683_1 | n2240;
  assign n1322 = n1678 | n1679_1 | n1680 | n2242;
  assign n1327 = n1675_1 | n1676 | n1677 | n2244;
  assign n1332 = n1672 | n1673 | n1674 | n2246;
  assign n1336 = n1669 | n1670 | n1671_1 | n2248;
  assign n1340 = n1666 | n1667_1 | n1668 | n2250;
  assign n1344 = n1663_1 | n1664 | n1665 | n2252;
  assign n1348 = n1660 | n1661 | n1662 | n2254;
  assign n1352 = n1657 | n1658 | n1659_1 | n2256;
  assign n1356 = n1654 | n1655_1 | n1656 | n2258;
  assign n1361 = n1651_1 | n1652 | n1653 | n2260;
  assign n1365 = n1648 | n1649 | n1650 | n2262;
  assign n1370 = n1645 | n1646 | n1647_1 | n2264;
  assign n1374 = n1642 | n1643_1 | n1644 | n2266;
  assign n1378 = n1639_1 | n1640 | n1641 | n2268;
  assign n1382 = n1636 | n1637 | n1638 | n2270;
  assign n1386 = n1633 | n1634 | n1635_1 | n2272;
  assign n1390 = n1630_1 | n1631 | n1632 | n2274;
  assign n1394 = n1627 | n1628 | n1629 | n2276;
  assign n1398 = n1624 | n1625 | n1626_1 | n2278;
  assign n1402 = n1621 | n1622_1 | n1623 | n2280;
  assign n1407 = n1618_1 | n1619 | n1620 | n2282;
  assign n1411 = n1615 | n1616 | n1617 | n2284;
  assign n1415 = n1612 | n1613_1 | n1614 | n2286;
  assign n1419 = n1609_1 | n1610 | n1611 | n2288;
  assign n1423 = n1606 | n1607 | n1608 | n2290;
  assign n1427 = n1603 | n1604 | n1605_1 | n2292;
  assign n1432 = n1600 | n1601_1 | n1602 | n2294;
  assign n1436 = n1597_1 | n1598 | n1599 | n2296;
  assign n1440 = n1594 | n1595 | n1596 | n2298;
  assign n1444 = n1591 | n1592 | n1593_1 | n2300;
  assign n1448 = n1588 | n1589_1 | n1590 | n2302;
  assign n1452 = n1585 | n1586 | n1587 | n2304;
  assign n1456 = n1582 | n1583 | n1584_1 | n2306;
  assign n1460 = n1579 | n1580_1 | n1581 | n2308;
  assign n1464 = n1576_1 | n1577 | n1578 | n2310;
  assign n1468 = n1573 | n1574 | n1575 | n2312;
  assign n1472 = n1570 | n1571 | n1572_1 | n2314;
  assign n1476 = n1567 | n1568_1 | n1569 | n2316;
  assign n1480 = n1564 | n1565 | n1566 | n2318;
  assign n1485 = n1561 | n1562 | n1563_1 | n2320;
  assign n1489 = n1558 | n1559_1 | n1560 | n2322;
  assign n1493 = n1555_1 | n1556 | n1557 | n2324;
  assign n1497 = n1552 | n1553 | n1554 | n2326;
  assign n1502 = n1549 | n1550 | n1551_1 | n2328;
  assign n1506 = n1546 | n1547_1 | n1548 | n2330;
  assign n1510 = n1543_1 | n1544 | n1545 | n2332;
  assign n1514 = n1540 | n1541 | n1542 | n2334;
  assign n1518 = n1537 | n1538_1 | n1539 | n2336;
  assign n1522 = n1534_1 | n1535 | n1536 | n2338;
  assign n1526 = n1531 | n1532 | n1533 | n2340;
  assign n1530 = n1528 | n1529 | n1530_1 | n2342;
  assign n1534 = n1525 | n1526_1 | n1527 | n2344;
  assign n1538 = n1522_1 | n1523 | n1524 | n2346;
  assign n1543 = n1519 | n1520 | n1521 | n2348;
  assign n1547 = n1516 | n1517 | n1518_1 | n2350;
  assign n1551 = n1513 | n1514_1 | n1515 | n2352;
  assign n1555 = n1510_1 | n1511 | n1512 | n2354;
  assign n1559 = n1507 | n1508 | n1509 | n2356;
  assign n1563 = n1504 | n1505 | n1506_1 | n2358;
  assign n1568 = n1501 | n1502_1 | n1503 | n2360;
  assign n1572 = n1498 | n1499 | n1500 | n2362;
  assign n1576 = n1495 | n1496 | n1497_1 | n2364;
  assign n1580 = n1492 | n1493_1 | n1494 | n2366;
  assign n1584 = n1489_1 | n1490 | n1491 | n2368;
  assign n1589 = n1486 | n1487 | n1488 | n2370;
  assign n1593 = n1483 | n1484 | n1485_1 | n2372;
  assign n1597 = n1480_1 | n1481 | n1482 | n2374;
  assign n1601 = n1477 | n1478 | n1479 | n2376;
  assign n1605 = n1474 | n1475 | n1476_1 | n2378;
  assign n1609 = n1471 | n1472_1 | n1473 | n2380;
  assign n1613 = n1468_1 | n1469 | n1470 | n2382;
  assign n1618 = n1465 | n1466 | n1467 | n2384;
  assign n1622 = n1462 | n1463 | n1464_1 | n2386;
  assign n1626 = n1459 | n1460_1 | n1461 | n2388;
  assign n1630 = n1456_1 | n1457 | n1458 | n2390;
  assign n1635 = n1453 | n1454 | n1455 | n2392;
  assign n1639 = n1450 | n1451 | n1452_1 | n2394;
  assign n1643 = n1447 | n1448_1 | n1449 | n2396;
  assign n1647 = n1444_1 | n1445 | n1446 | n2398;
  assign n1651 = n1441 | n1442 | n1443 | n2400;
  assign n1655 = n1438 | n1439 | n1440_1 | n2402;
  assign n1659 = n1435 | n1436_1 | n1437 | n2404;
  assign n1663 = n1432_1 | n1433 | n1434 | n2406;
  assign n1667 = n1429 | n1430 | n1431 | n2408;
  assign n1671 = n1426 | n1427_1 | n1428 | n2410;
  assign n1675 = n1423_1 | n1424 | n1425 | n2412;
  assign n1679 = n1420 | n1421 | n1422 | n2414;
  assign n1683 = n1417 | n1418 | n1419_1 | n2416;
  assign n1687 = n1414 | n1415_1 | n1416 | n2418;
  assign n1691 = n1411_1 | n1412 | n1413 | n2420;
  assign n1696 = n1408 | n1409 | n1410 | n2422;
  assign n1701 = n1405 | n1406 | n1407_1 | n2424;
  assign n1706 = n1402_1 | n1403 | n1404 | n2426;
  assign n1710 = n1399 | n1400 | n1401 | n2428;
  assign n1714 = n1396 | n1397 | n1398_1 | n2430;
  assign n1718 = n1393 | n1394_1 | n1395 | n2432;
  assign n1722 = n1390_1 | n1391 | n1392 | n2434;
  assign n1726 = n1387 | n1388 | n1389 | n2436;
  assign n1730 = n1384 | n1385 | n1386_1 | n2438;
  assign n1735 = n1381 | n1382_1 | n1383 | n2440;
  assign n1739 = n1378_1 | n1379 | n1380 | n2442;
  assign n1743 = n1375 | n1376 | n1377 | n2444;
  assign n1747 = n1372 | n1373 | n1374_1 | n2446;
  assign n1751 = n1369 | n1370_1 | n1371 | n2448;
  assign n1755 = n1366 | n1367 | n1368 | n2450;
  assign n1759 = n1363 | n1364 | n1365_1 | n2452;
  assign n1763 = n1360 | n1361_1 | n1362 | n2454;
  assign n1767 = n1357 | n1358 | n1359 | n2456;
  assign n1771 = n1354 | n1355 | n1356_1 | n2458;
  assign n1776 = n1351 | n1352_1 | n1353 | n2460;
  assign n1781 = n1348_1 | n1349 | n1350 | n2462;
  assign n1785 = n1345 | n1346 | n1347 | n2464;
  assign n1327_1 = (~pcount_3_ & (pcount_2_ ? (pcount_1_ & pcount_0_) : (~pcount_1_ & ~pcount_0_))) | (pcount_1_ & ~pcount_0_ & pcount_3_ & pcount_2_);
  assign n1328 = (~pcount_2_ & ~pcount_1_ & (~pcount_3_ | ~pcount_0_)) | (pcount_1_ & pcount_0_ & pcount_3_ & pcount_2_);
  assign n1329 = pencrypt_0_ & ~pstart_0_ & pcount_1_ & pcount_0_;
  assign n1330 = ~pstart_0_ | pencrypt_0_;
  assign n1331 = (pencrypt_0_ & (pstart_0_ | (pcount_1_ & pcount_0_))) | (~pcount_1_ & ~pcount_0_ & ~pencrypt_0_);
  assign n1332_1 = ~pstart_0_ & pencrypt_0_;
  assign pksi_90_ = n_n10;
  assign pksi_191_ = n_n121;
  assign pksi_187_ = n_n121;
  assign pksi_168_ = n_n109;
  assign pksi_181_ = n_n109;
  assign pksi_88_ = n_n10;
  assign pksi_143_ = n_n168;
  assign pksi_139_ = n_n168;
  assign n1341 = ~pencrypt_0_ & ~pcount_0_ & ~pcount_2_ & ~pcount_1_;
  assign n1342 = ~pcount_3_ & (n1344_1 | (pcount_2_ & n1329));
  assign n1343 = pcount_3_ & (~n1331 | n2466);
  assign n1344_1 = ~pencrypt_0_ & ~pcount_0_ & ~pcount_2_ & ~pcount_1_;
  assign n1345 = n1328 & n_n2374 & ~pstart_0_ & ~pencrypt_0_;
  assign n1346 = ~n1328 & pksi_1_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1347 = ~n1327_1 & pksi_10_ & ~pstart_0_ & pencrypt_0_;
  assign n1348_1 = ~n1328 & pksi_16_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1349 = n1328 & pksi_20_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1350 = ~n1327_1 & pksi_47_ & ~pstart_0_ & pencrypt_0_;
  assign n1351 = ~n1328 & pksi_43_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1352_1 = n1328 & pksi_41_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1353 = ~n1327_1 & pksi_26_ & ~pstart_0_ & pencrypt_0_;
  assign n1354 = ~n1328 & pksi_42_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1355 = n1328 & pksi_25_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1356_1 = ~n1327_1 & pksi_45_ & ~pstart_0_ & pencrypt_0_;
  assign n1357 = ~n1328 & n_n2333 & ~pstart_0_ & ~pencrypt_0_;
  assign n1358 = n1328 & pksi_40_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1359 = ~n1327_1 & pksi_52_ & ~pstart_0_ & pencrypt_0_;
  assign n1360 = ~n1328 & pksi_57_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1361_1 = n1328 & pksi_67_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1362 = ~n1327_1 & pksi_59_ & ~pstart_0_ & pencrypt_0_;
  assign n1363 = ~n1328 & pksi_56_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1364 = n1328 & pksi_66_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1365_1 = ~n1327_1 & pksi_61_ & ~pstart_0_ & pencrypt_0_;
  assign n1366 = ~n1328 & n_n2374 & ~pstart_0_ & ~pencrypt_0_;
  assign n1367 = n1327_1 & pksi_10_ & ~pstart_0_ & pencrypt_0_;
  assign n1368 = n1328 & pksi_13_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1369 = ~n1328 & n_n2365 & ~pstart_0_ & ~pencrypt_0_;
  assign n1370_1 = n1328 & pksi_16_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1371 = ~n1327_1 & pksi_28_ & ~pstart_0_ & pencrypt_0_;
  assign n1372 = n1328 & n_n2352 & ~pstart_0_ & ~pencrypt_0_;
  assign n1373 = ~n1328 & pksi_41_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1374_1 = ~n1327_1 & pksi_38_ & ~pstart_0_ & pencrypt_0_;
  assign n1375 = ~n1328 & pksi_32_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1376 = n1328 & pksi_42_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1377 = ~n1327_1 & pksi_37_ & ~pstart_0_ & pencrypt_0_;
  assign n1378_1 = ~n1328 & pksi_40_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1379 = n1328 & pksi_44_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1380 = ~n1327_1 & pksi_71_ & ~pstart_0_ & pencrypt_0_;
  assign n1381 = ~n1328 & pksi_53_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1382_1 = n1327_1 & pksi_65_ & ~pstart_0_ & pencrypt_0_;
  assign n1383 = n1328 & pksi_57_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1384 = ~n1328 & pksi_66_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1385 = n1328 & pksi_49_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1386_1 = ~n1327_1 & pksi_69_ & ~pstart_0_ & pencrypt_0_;
  assign n1387 = ~n1328 & pksi_13_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1388 = n1328 & pksi_21_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1389 = ~n1327_1 & pksi_12_ & ~pstart_0_ & pencrypt_0_;
  assign n1390_1 = n1328 & n_n2365 & ~pstart_0_ & ~pencrypt_0_;
  assign n1391 = ~n1328 & pksi_3_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1392 = ~n1327_1 & pksi_7_ & ~pstart_0_ & pencrypt_0_;
  assign n1393 = ~n1328 & pksi_29_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1394_1 = n1327_1 & pksi_41_ & ~pstart_0_ & pencrypt_0_;
  assign n1395 = n1328 & pksi_33_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1396 = ~n1328 & n_n2342 & ~pstart_0_ & ~pencrypt_0_;
  assign n1397 = n1327_1 & pksi_34_ & ~pstart_0_ & pencrypt_0_;
  assign n1398_1 = n1328 & pksi_37_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1399 = ~n1328 & pksi_44_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1400 = n1328 & pksi_31_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1401 = ~n1327_1 & pksi_54_ & ~pstart_0_ & pencrypt_0_;
  assign n1402_1 = ~n1328 & pksi_64_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1403 = n1328 & pksi_68_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1404 = ~n1327_1 & pksi_95_ & ~pstart_0_ & pencrypt_0_;
  assign n1405 = ~n1328 & pksi_91_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1406 = n1328 & pksi_89_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1407_1 = ~n1327_1 & pksi_74_ & ~pstart_0_ & pencrypt_0_;
  assign n1408 = ~n1328 & pksi_21_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1409 = n1328 & pksi_10_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1410 = ~n1327_1 & pksi_3_ & ~pstart_0_ & pencrypt_0_;
  assign n1411_1 = ~n1328 & pksi_12_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1412 = n1328 & pksi_3_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1413 = ~n1327_1 & pksi_20_ & ~pstart_0_ & pencrypt_0_;
  assign n1414 = ~n1328 & pksi_33_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1415_1 = n1328 & pksi_43_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1416 = ~n1327_1 & pksi_35_ & ~pstart_0_ & pencrypt_0_;
  assign n1417 = n1328 & n_n2342 & ~pstart_0_ & ~pencrypt_0_;
  assign n1418 = ~n1328 & pksi_25_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1419_1 = ~n1327_1 & pksi_34_ & ~pstart_0_ & pencrypt_0_;
  assign n1420 = ~n1328 & pksi_31_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1421 = n1328 & pksi_52_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1422 = ~n1327_1 & pksi_63_ & ~pstart_0_ & pencrypt_0_;
  assign n1423_1 = ~n1328 & n_n2301 & ~pstart_0_ & ~pencrypt_0_;
  assign n1424 = n1328 & pksi_64_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1425 = ~n1327_1 & pksi_76_ & ~pstart_0_ & pencrypt_0_;
  assign n1426 = ~n1328 & pksi_89_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1427_1 = n1328 & n_n2288 & ~pstart_0_ & ~pencrypt_0_;
  assign n1428 = ~n1327_1 & pksi_86_ & ~pstart_0_ & pencrypt_0_;
  assign n1429 = ~n1328 & n_n2369 & ~pstart_0_ & ~pencrypt_0_;
  assign n1430 = n1328 & pksi_12_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1431 = ~n1327_1 & pksi_16_ & ~pstart_0_ & pencrypt_0_;
  assign n1432_1 = ~n1328 & pksi_30_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1433 = n1328 & pksi_39_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1434 = ~n1327_1 & pksi_43_ & ~pstart_0_ & pencrypt_0_;
  assign n1435 = ~n1328 & pksi_59_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1436_1 = n1328 & pksi_50_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1437 = ~n1327_1 & pksi_48_ & ~pstart_0_ & pencrypt_0_;
  assign n1438 = ~n1328 & pksi_61_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1439 = n1328 & pksi_69_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1440_1 = ~n1327_1 & pksi_60_ & ~pstart_0_ & pencrypt_0_;
  assign n1441 = ~n1328 & pksi_55_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1442 = n1328 & pksi_76_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1443 = ~n1327_1 & pksi_87_ & ~pstart_0_ & pencrypt_0_;
  assign n1444_1 = ~n1328 & n_n2288 & ~pstart_0_ & ~pencrypt_0_;
  assign n1445 = n1328 & pksi_83_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1446 = ~n1327_1 & pksi_94_ & ~pstart_0_ & pencrypt_0_;
  assign n1447 = n1328 & n_n2369 & ~pstart_0_ & ~pencrypt_0_;
  assign n1448_1 = ~n1328 & pksi_10_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1449 = n1327_1 & pksi_3_ & ~pstart_0_ & pencrypt_0_;
  assign n1450 = ~n1328 & pksi_39_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1451 = n1328 & pksi_29_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1452_1 = ~n1327_1 & pksi_41_ & ~pstart_0_ & pencrypt_0_;
  assign n1453 = ~n1328 & n_n2320 & ~pstart_0_ & ~pencrypt_0_;
  assign n1454 = n1328 & pksi_59_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1455 = ~n1327_1 & pksi_70_ & ~pstart_0_ & pencrypt_0_;
  assign n1456_1 = ~n1328 & pksi_69_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1457 = n1328 & pksi_58_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1458 = ~n1327_1 & pksi_51_ & ~pstart_0_ & pencrypt_0_;
  assign n1459 = ~n1328 & pksi_68_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1460_1 = n1328 & pksi_55_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1461 = ~n1327_1 & pksi_78_ & ~pstart_0_ & pencrypt_0_;
  assign n1462 = ~n1328 & pksi_83_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1463 = n1328 & pksi_74_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1464_1 = ~n1327_1 & pksi_72_ & ~pstart_0_ & pencrypt_0_;
  assign n1465 = ~n1328 & pksi_24_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1466 = n1327_1 & pksi_25_ & ~pstart_0_ & pencrypt_0_;
  assign n1467 = n1328 & pksi_32_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1468_1 = ~n1328 & pksi_36_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1469 = n1328 & pksi_27_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1470 = ~n1327_1 & pksi_44_ & ~pstart_0_ & pencrypt_0_;
  assign n1471 = n1328 & n_n2320 & ~pstart_0_ & ~pencrypt_0_;
  assign n1472_1 = ~n1328 & pksi_65_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1473 = ~n1327_1 & pksi_62_ & ~pstart_0_ & pencrypt_0_;
  assign n1474 = ~n1328 & pksi_49_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1475 = n1328 & n_n2310 & ~pstart_0_ & ~pencrypt_0_;
  assign n1476_1 = ~n1327_1 & pksi_58_ & ~pstart_0_ & pencrypt_0_;
  assign n1477 = ~n1328 & pksi_95_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1478 = n1328 & pksi_78_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1479 = ~n1327_1 & pksi_81_ & ~pstart_0_ & pencrypt_0_;
  assign n1480_1 = ~n1328 & pksi_74_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1481 = n1328 & pksi_86_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1482 = ~n1327_1 & pksi_80_ & ~pstart_0_ & pencrypt_0_;
  assign n1483 = ~n1328 & pksi_46_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1484 = n1328 & pksi_24_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1485_1 = ~n1327_1 & pksi_25_ & ~pstart_0_ & pencrypt_0_;
  assign n1486 = n1328 & n_n2333 & ~pstart_0_ & ~pencrypt_0_;
  assign n1487 = ~n1328 & pksi_27_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1488 = ~n1327_1 & pksi_31_ & ~pstart_0_ & pencrypt_0_;
  assign n1489_1 = ~n1328 & pksi_67_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1490 = n1328 & pksi_65_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1491 = ~n1327_1 & pksi_50_ & ~pstart_0_ & pencrypt_0_;
  assign n1492 = ~n1328 & n_n2310 & ~pstart_0_ & ~pencrypt_0_;
  assign n1493_1 = ~n1327_1 & n_n2305 & ~pstart_0_ & pencrypt_0_;
  assign n1494 = n1328 & pksi_61_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1495 = ~n1328 & pksi_76_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1496 = n1328 & pksi_95_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1497_1 = ~n1327_1 & pksi_77_ & ~pstart_0_ & pencrypt_0_;
  assign n1498 = ~n1328 & pksi_86_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1499 = ~n1327_1 & n_n2280 & ~pstart_0_ & pencrypt_0_;
  assign n1500 = n1328 & pksi_94_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1501 = ~n1328 & pksi_48_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1502_1 = n1328 & pksi_56_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1503 = ~n1327_1 & n_n2310 & ~pstart_0_ & pencrypt_0_;
  assign n1504 = ~n1328 & pksi_60_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1505 = n1328 & pksi_51_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1506_1 = ~n1327_1 & pksi_68_ & ~pstart_0_ & pencrypt_0_;
  assign n1507 = ~n1328 & pksi_87_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1508 = n1328 & pksi_77_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1509 = ~n1327_1 & pksi_89_ & ~pstart_0_ & pencrypt_0_;
  assign n1510_1 = ~n1328 & pksi_94_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1511 = n1328 & pksi_72_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1512 = ~n1327_1 & pksi_73_ & ~pstart_0_ & pencrypt_0_;
  assign n1513 = ~n1328 & pksi_70_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1514_1 = n1328 & pksi_48_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1515 = ~n1327_1 & pksi_49_ & ~pstart_0_ & pencrypt_0_;
  assign n1516 = ~n1328 & pksi_51_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1517 = n1328 & n_n2301 & ~pstart_0_ & ~pencrypt_0_;
  assign n1518_1 = ~n1327_1 & pksi_55_ & ~pstart_0_ & pencrypt_0_;
  assign n1519 = ~n1328 & pksi_78_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1520 = n1328 & pksi_87_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1521 = ~n1327_1 & pksi_91_ & ~pstart_0_ & pencrypt_0_;
  assign n1522_1 = ~n1328 & pksi_72_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1523 = n1327_1 & pksi_73_ & ~pstart_0_ & pencrypt_0_;
  assign n1524 = n1328 & pksi_80_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1525 = ~n1328 & pksi_2_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1526_1 = n1328 & pksi_14_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1527 = ~n1327_1 & pksi_8_ & ~pstart_0_ & pencrypt_0_;
  assign n1528 = ~n1328 & pksi_62_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1529 = n1328 & pksi_70_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1530_1 = ~n1327_1 & pksi_66_ & ~pstart_0_ & pencrypt_0_;
  assign n1531 = ~n1328 & pksi_58_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1532 = n1328 & n_n2305 & ~pstart_0_ & ~pencrypt_0_;
  assign n1533 = ~n1327_1 & n_n2301 & ~pstart_0_ & pencrypt_0_;
  assign n1534_1 = ~n1328 & pksi_81_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1535 = n1328 & pksi_91_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1536 = ~n1327_1 & pksi_83_ & ~pstart_0_ & pencrypt_0_;
  assign n1537 = ~n1328 & pksi_80_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1538_1 = n1328 & n_n2280 & ~pstart_0_ & ~pencrypt_0_;
  assign n1539 = ~n1327_1 & pksi_85_ & ~pstart_0_ & pencrypt_0_;
  assign n1540 = ~n1328 & pksi_14_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1541 = n1328 & pksi_22_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1542 = ~n1327_1 & pksi_18_ & ~pstart_0_ & pencrypt_0_;
  assign n1543_1 = ~n1328 & pksi_50_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1544 = n1328 & pksi_62_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1545 = ~n1327_1 & pksi_56_ & ~pstart_0_ & pencrypt_0_;
  assign n1546 = ~n1328 & n_n2305 & ~pstart_0_ & ~pencrypt_0_;
  assign n1547_1 = n1328 & pksi_60_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1548 = ~n1327_1 & pksi_64_ & ~pstart_0_ & pencrypt_0_;
  assign n1549 = ~n1328 & pksi_77_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1550 = n1328 & pksi_81_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1551_1 = ~n1327_1 & n_n2288 & ~pstart_0_ & pencrypt_0_;
  assign n1552 = ~n1328 & n_n2280 & ~pstart_0_ & ~pencrypt_0_;
  assign n1553 = n1328 & pksi_73_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1554 = ~n1327_1 & pksi_93_ & ~pstart_0_ & pencrypt_0_;
  assign n1555_1 = ~n1328 & pksi_22_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1556 = n1328 & pksi_0_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1557 = ~n1327_1 & pksi_1_ & ~pstart_0_ & pencrypt_0_;
  assign n1558 = ~n1328 & pksi_47_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1559_1 = n1328 & pksi_30_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1560 = ~n1327_1 & pksi_33_ & ~pstart_0_ & pencrypt_0_;
  assign n1561 = ~n1328 & pksi_26_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1562 = n1328 & pksi_38_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1563_1 = ~n1327_1 & pksi_32_ & ~pstart_0_ & pencrypt_0_;
  assign n1564 = ~n1328 & pksi_45_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1565 = n1328 & pksi_34_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1566 = ~n1327_1 & pksi_27_ & ~pstart_0_ & pencrypt_0_;
  assign n1567 = ~n1328 & pksi_52_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1568_1 = n1328 & pksi_71_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1569 = ~n1327_1 & pksi_53_ & ~pstart_0_ & pencrypt_0_;
  assign n1570 = ~n1328 & n_n10 & ~pstart_0_ & ~pencrypt_0_;
  assign n1571 = n1328 & pksi_92_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1572_1 = ~n1327_1 & pksi_23_ & ~pstart_0_ & pencrypt_0_;
  assign n1573 = ~n1328 & pksi_0_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1574 = n1327_1 & pksi_1_ & ~pstart_0_ & pencrypt_0_;
  assign n1575 = n1328 & pksi_8_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1576_1 = ~n1328 & pksi_28_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1577 = n1328 & pksi_47_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1578 = ~n1327_1 & pksi_29_ & ~pstart_0_ & pencrypt_0_;
  assign n1579 = ~n1328 & pksi_38_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1580_1 = n1328 & pksi_46_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1581 = ~n1327_1 & pksi_42_ & ~pstart_0_ & pencrypt_0_;
  assign n1582 = ~n1328 & pksi_37_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1583 = n1328 & pksi_45_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1584_1 = ~n1327_1 & pksi_36_ & ~pstart_0_ & pencrypt_0_;
  assign n1585 = ~n1328 & pksi_71_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1586 = n1328 & pksi_54_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1587 = ~n1327_1 & pksi_57_ & ~pstart_0_ & pencrypt_0_;
  assign n1588 = ~n1328 & pksi_8_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1589_1 = n1328 & pksi_18_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1590 = ~n1327_1 & pksi_13_ & ~pstart_0_ & pencrypt_0_;
  assign n1591 = ~n1328 & pksi_7_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1592 = n1328 & pksi_28_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1593_1 = ~n1327_1 & pksi_39_ & ~pstart_0_ & pencrypt_0_;
  assign n1594 = ~n1328 & n_n2352 & ~pstart_0_ & ~pencrypt_0_;
  assign n1595 = n1328 & pksi_35_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1596 = ~n1327_1 & pksi_46_ & ~pstart_0_ & pencrypt_0_;
  assign n1597_1 = ~n1328 & n_n2337 & ~pstart_0_ & ~pencrypt_0_;
  assign n1598 = n1328 & pksi_36_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1599 = ~n1327_1 & pksi_40_ & ~pstart_0_ & pencrypt_0_;
  assign n1600 = ~n1328 & pksi_54_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1601_1 = n1328 & pksi_63_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1602 = ~n1327_1 & pksi_67_ & ~pstart_0_ & pencrypt_0_;
  assign n1603 = ~n1328 & pksi_18_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1604 = n1328 & pksi_1_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1605_1 = ~n1327_1 & pksi_21_ & ~pstart_0_ & pencrypt_0_;
  assign n1606 = ~n1328 & pksi_20_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1607 = n1328 & pksi_7_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1608 = ~n1327_1 & pksi_30_ & ~pstart_0_ & pencrypt_0_;
  assign n1609_1 = ~n1328 & pksi_35_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1610 = n1328 & pksi_26_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1611 = ~n1327_1 & pksi_24_ & ~pstart_0_ & pencrypt_0_;
  assign n1612 = n1328 & n_n2337 & ~pstart_0_ & ~pencrypt_0_;
  assign n1613_1 = ~n1328 & pksi_34_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1614 = n1327_1 & pksi_27_ & ~pstart_0_ & pencrypt_0_;
  assign n1615 = ~n1328 & pksi_63_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1616 = n1328 & pksi_53_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1617 = ~n1327_1 & pksi_65_ & ~pstart_0_ & pencrypt_0_;
  assign n1618_1 = ~n1328 & pksi_98_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1619 = n1327_1 & pksi_112_ & ~pstart_0_ & pencrypt_0_;
  assign n1620 = n1328 & pksi_119_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1621 = ~n1328 & pksi_126_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1622_1 = n1328 & pksi_122_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1623 = ~n1327_1 & pksi_136_ & ~pstart_0_ & pencrypt_0_;
  assign n1624 = ~n1328 & pksi_134_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1625 = n1327_1 & n_n2476 & ~pstart_0_ & pencrypt_0_;
  assign n1626_1 = n1328 & pksi_127_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1627 = ~n1328 & pksi_131_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1628 = n1328 & pksi_133_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1629 = ~n1327_1 & pksi_121_ & ~pstart_0_ & pencrypt_0_;
  assign n1630_1 = ~n1328 & pksi_166_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1631 = n1328 & pksi_150_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1632 = ~n1327_1 & pksi_154_ & ~pstart_0_ & pencrypt_0_;
  assign n1633 = ~n1328 & n_n2448 & ~pstart_0_ & ~pencrypt_0_;
  assign n1634 = n1328 & pksi_158_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1635_1 = ~n1327_1 & pksi_163_ & ~pstart_0_ & pencrypt_0_;
  assign n1636 = ~n1328 & pksi_148_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1637 = n1328 & pksi_155_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1638 = ~n1327_1 & pksi_152_ & ~pstart_0_ & pencrypt_0_;
  assign n1639_1 = ~n1328 & pksi_159_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1640 = n1328 & pksi_190_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1641 = ~n1327_1 & n_n121 & ~pstart_0_ & pencrypt_0_;
  assign n1642 = ~n1328 & pksi_171_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1643_1 = n1328 & n_n2416 & ~pstart_0_ & ~pencrypt_0_;
  assign n1644 = ~n1327_1 & n_n2412 & ~pstart_0_ & pencrypt_0_;
  assign n1645 = ~n1328 & n_n2272 & ~pstart_0_ & ~pencrypt_0_;
  assign n1646 = n1328 & pksi_84_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1647_1 = ~n1327_1 & n_n10 & ~pstart_0_ & pencrypt_0_;
  assign n1648 = ~n1328 & pksi_96_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1649 = n1328 & pksi_115_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1650 = ~n1327_1 & pksi_105_ & ~pstart_0_ & pencrypt_0_;
  assign n1651_1 = ~n1328 & pksi_142_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1652 = n1328 & pksi_126_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1653 = ~n1327_1 & pksi_130_ & ~pstart_0_ & pencrypt_0_;
  assign n1654 = ~n1328 & pksi_127_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1655_1 = n1328 & pksi_120_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1656 = ~n1327_1 & pksi_132_ & ~pstart_0_ & pencrypt_0_;
  assign n1657 = ~n1328 & pksi_124_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1658 = n1328 & pksi_131_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1659_1 = ~n1327_1 & pksi_128_ & ~pstart_0_ & pencrypt_0_;
  assign n1660 = ~n1328 & pksi_150_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1661 = n1328 & pksi_146_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1662 = ~n1327_1 & pksi_160_ & ~pstart_0_ & pencrypt_0_;
  assign n1663_1 = ~n1328 & pksi_147_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1664 = n1328 & n_n2448 & ~pstart_0_ & ~pencrypt_0_;
  assign n1665 = ~n1327_1 & pksi_144_ & ~pstart_0_ & pencrypt_0_;
  assign n1666 = ~n1328 & pksi_155_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1667_1 = n1328 & pksi_157_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1668 = ~n1327_1 & pksi_145_ & ~pstart_0_ & pencrypt_0_;
  assign n1669 = ~n1328 & pksi_149_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1670 = n1328 & pksi_159_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1671_1 = ~n1327_1 & pksi_170_ & ~pstart_0_ & pencrypt_0_;
  assign n1672 = ~n1328 & n_n2416 & ~pstart_0_ & ~pencrypt_0_;
  assign n1673 = n1328 & pksi_182_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1674 = ~n1327_1 & n_n2410 & ~pstart_0_ & pencrypt_0_;
  assign n1675_1 = ~n1328 & pksi_84_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1676 = n1328 & pksi_75_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1677 = ~n1327_1 & pksi_92_ & ~pstart_0_ & pencrypt_0_;
  assign n1678 = ~n1328 & pksi_106_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1679_1 = n1328 & pksi_112_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1680 = ~n1327_1 & pksi_99_ & ~pstart_0_ & pencrypt_0_;
  assign n1681 = ~n1328 & pksi_115_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1682 = n1328 & n_n2507 & ~pstart_0_ & ~pencrypt_0_;
  assign n1683_1 = ~n1327_1 & pksi_114_ & ~pstart_0_ & pencrypt_0_;
  assign n1684 = ~n1328 & n_n168 & ~pstart_0_ & ~pencrypt_0_;
  assign n1685 = n1328 & pksi_130_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1686 = ~n1327_1 & pksi_141_ & ~pstart_0_ & pencrypt_0_;
  assign n1687_1 = ~n1328 & pksi_120_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1688 = n1328 & n_n2476 & ~pstart_0_ & ~pencrypt_0_;
  assign n1689 = ~n1327_1 & pksi_129_ & ~pstart_0_ & pencrypt_0_;
  assign n1690 = ~n1328 & pksi_138_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1691_1 = n1328 & pksi_124_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1692 = ~n1327_1 & pksi_140_ & ~pstart_0_ & pencrypt_0_;
  assign n1693 = ~n1328 & pksi_125_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1694 = n1328 & pksi_135_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1695 = ~n1327_1 & pksi_146_ & ~pstart_0_ & pencrypt_0_;
  assign n1696_1 = ~n1328 & pksi_151_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1697 = n1328 & pksi_144_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1698 = ~n1327_1 & pksi_156_ & ~pstart_0_ & pencrypt_0_;
  assign n1699 = ~n1328 & pksi_157_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1700 = n1328 & pksi_164_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1701_1 = ~n1327_1 & pksi_161_ & ~pstart_0_ & pencrypt_0_;
  assign n1702 = ~n1328 & pksi_179_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1703 = n1328 & n_n109 & ~pstart_0_ & ~pencrypt_0_;
  assign n1704 = ~n1327_1 & pksi_169_ & ~pstart_0_ & pencrypt_0_;
  assign n1705 = ~n1328 & pksi_4_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1706_1 = n1328 & pksi_23_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1707 = ~n1327_1 & pksi_5_ & ~pstart_0_ & pencrypt_0_;
  assign n1708 = n1328 & n_n2268 & ~pstart_0_ & ~pencrypt_0_;
  assign n1709 = ~n1328 & pksi_75_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1710_1 = ~n1327_1 & pksi_79_ & ~pstart_0_ & pencrypt_0_;
  assign n1711 = ~n1328 & pksi_119_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1712 = n1328 & pksi_106_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1713 = ~n1327_1 & pksi_117_ & ~pstart_0_ & pencrypt_0_;
  assign n1714_1 = ~n1328 & n_n2507 & ~pstart_0_ & ~pencrypt_0_;
  assign n1715 = n1328 & pksi_108_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1716 = ~n1327_1 & pksi_100_ & ~pstart_0_ & pencrypt_0_;
  assign n1717 = ~n1328 & pksi_122_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1718_1 = ~n1327_1 & n_n2485 & ~pstart_0_ & pencrypt_0_;
  assign n1719 = n1328 & n_n168 & ~pstart_0_ & ~pencrypt_0_;
  assign n1720 = n1328 & n_n2474 & ~pstart_0_ & ~pencrypt_0_;
  assign n1721 = ~n1328 & n_n2476 & ~pstart_0_ & ~pencrypt_0_;
  assign n1722_1 = ~n1327_1 & pksi_138_ & ~pstart_0_ & pencrypt_0_;
  assign n1723 = ~n1328 & pksi_129_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1724 = n1328 & pksi_138_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1725 = ~n1327_1 & pksi_133_ & ~pstart_0_ & pencrypt_0_;
  assign n1726_1 = ~n1328 & pksi_135_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1727 = n1328 & pksi_166_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1728 = ~n1327_1 & pksi_167_ & ~pstart_0_ & pencrypt_0_;
  assign n1729 = ~n1328 & pksi_158_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1730_1 = n1328 & pksi_151_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1731 = ~n1327_1 & pksi_153_ & ~pstart_0_ & pencrypt_0_;
  assign n1732 = ~n1328 & pksi_164_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1733 = n1327_1 & pksi_161_ & ~pstart_0_ & pencrypt_0_;
  assign n1734 = n1328 & pksi_152_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1735_1 = ~n1328 & pksi_172_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1736 = n1328 & pksi_179_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1737 = ~n1327_1 & pksi_176_ & ~pstart_0_ & pencrypt_0_;
  assign n1738 = ~n1328 & pksi_23_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1739_1 = n1328 & pksi_6_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1740 = ~n1327_1 & pksi_9_ & ~pstart_0_ & pencrypt_0_;
  assign n1741 = ~n1328 & n_n2268 & ~pstart_0_ & ~pencrypt_0_;
  assign n1742 = n1328 & n_n10 & ~pstart_0_ & ~pencrypt_0_;
  assign n1743_1 = ~n1327_1 & pksi_4_ & ~pstart_0_ & pencrypt_0_;
  assign n1744 = ~n1328 & n_n2495 & ~pstart_0_ & ~pencrypt_0_;
  assign n1745 = n1328 & pksi_101_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1746 = ~n1327_1 & pksi_126_ & ~pstart_0_ & pencrypt_0_;
  assign n1747_1 = ~n1328 & n_n2485 & ~pstart_0_ & ~pencrypt_0_;
  assign n1748 = n1328 & pksi_141_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1749 = ~n1327_1 & pksi_134_ & ~pstart_0_ & pencrypt_0_;
  assign n1750 = ~n1328 & pksi_121_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1751_1 = n1328 & pksi_137_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1752 = ~n1327_1 & pksi_135_ & ~pstart_0_ & pencrypt_0_;
  assign n1753 = ~n1328 & pksi_154_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1754 = n1328 & pksi_160_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1755_1 = ~n1327_1 & pksi_147_ & ~pstart_0_ & pencrypt_0_;
  assign n1756 = ~n1328 & pksi_163_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1757 = n1328 & pksi_153_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1758 = ~n1327_1 & pksi_162_ & ~pstart_0_ & pencrypt_0_;
  assign n1759_1 = ~n1328 & pksi_152_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1760 = n1328 & pksi_145_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1761 = ~n1327_1 & pksi_149_ & ~pstart_0_ & pencrypt_0_;
  assign n1762 = ~n1328 & n_n2277 & ~pstart_0_ & ~pencrypt_0_;
  assign n1763_1 = ~n1327_1 & n_n2272 & ~pstart_0_ & pencrypt_0_;
  assign n1764 = n1328 & pksi_85_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1765 = ~n1328 & pksi_113_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1766 = n1328 & n_n2495 & ~pstart_0_ & ~pencrypt_0_;
  assign n1767_1 = ~n1327_1 & pksi_142_ & ~pstart_0_ & pencrypt_0_;
  assign n1768 = ~n1328 & pksi_141_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1769 = n1328 & pksi_123_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1770 = ~n1327_1 & pksi_127_ & ~pstart_0_ & pencrypt_0_;
  assign n1771_1 = ~n1328 & pksi_128_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1772 = n1328 & pksi_121_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1773 = ~n1327_1 & pksi_125_ & ~pstart_0_ & pencrypt_0_;
  assign n1774 = n1328 & n_n2452 & ~pstart_0_ & ~pencrypt_0_;
  assign n1775 = ~n1328 & pksi_160_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1776_1 = ~n1327_1 & n_n2448 & ~pstart_0_ & pencrypt_0_;
  assign n1777 = ~n1328 & pksi_144_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1778 = ~n1327_1 & n_n2440 & ~pstart_0_ & pencrypt_0_;
  assign n1779 = n1328 & pksi_163_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1780 = ~n1328 & pksi_145_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1781_1 = n1328 & pksi_161_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1782 = ~n1327_1 & pksi_159_ & ~pstart_0_ & pencrypt_0_;
  assign n1783 = ~n1328 & pksi_85_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1784 = n1328 & pksi_93_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1785_1 = ~n1327_1 & pksi_84_ & ~pstart_0_ & pencrypt_0_;
  assign n1786 = ~n1328 & pksi_111_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1787 = n1328 & pksi_142_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1788 = ~n1327_1 & n_n168 & ~pstart_0_ & pencrypt_0_;
  assign n1789 = ~n1328 & pksi_123_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1790 = n1328 & n_n2481 & ~pstart_0_ & ~pencrypt_0_;
  assign n1791 = ~n1327_1 & pksi_120_ & ~pstart_0_ & pencrypt_0_;
  assign n1792 = ~n1328 & pksi_140_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1793 = n1327_1 & pksi_137_ & ~pstart_0_ & pencrypt_0_;
  assign n1794 = n1328 & pksi_128_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1795 = ~n1328 & pksi_146_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1796 = n1327_1 & pksi_160_ & ~pstart_0_ & pencrypt_0_;
  assign n1797 = n1328 & pksi_167_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1798 = ~n1328 & pksi_156_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1799 = n1328 & n_n2440 & ~pstart_0_ & ~pencrypt_0_;
  assign n1800 = ~n1327_1 & pksi_155_ & ~pstart_0_ & pencrypt_0_;
  assign n1801 = ~n1328 & pksi_161_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1802 = n1328 & n_n2430 & ~pstart_0_ & ~pencrypt_0_;
  assign n1803 = ~n1327_1 & pksi_190_ & ~pstart_0_ & pencrypt_0_;
  assign n1804 = ~n1328 & pksi_93_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1805 = n1328 & pksi_82_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1806 = ~n1327_1 & pksi_75_ & ~pstart_0_ & pencrypt_0_;
  assign n1807 = ~n1328 & pksi_101_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1808 = n1328 & pksi_111_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1809 = ~n1327_1 & pksi_122_ & ~pstart_0_ & pencrypt_0_;
  assign n1810 = ~n1328 & n_n2481 & ~pstart_0_ & ~pencrypt_0_;
  assign n1811 = n1327_1 & pksi_120_ & ~pstart_0_ & pencrypt_0_;
  assign n1812 = n1328 & pksi_134_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1813 = ~n1328 & pksi_133_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1814 = n1328 & pksi_140_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1815 = ~n1327_1 & pksi_137_ & ~pstart_0_ & pencrypt_0_;
  assign n1816 = ~n1328 & pksi_167_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1817 = n1328 & pksi_154_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1818 = ~n1327_1 & pksi_165_ & ~pstart_0_ & pencrypt_0_;
  assign n1819 = ~n1328 & pksi_153_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1820 = n1328 & pksi_156_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1821 = ~n1327_1 & pksi_148_ & ~pstart_0_ & pencrypt_0_;
  assign n1822 = ~n1328 & n_n2430 & ~pstart_0_ & ~pencrypt_0_;
  assign n1823 = n1328 & pksi_149_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1824 = ~n1327_1 & pksi_174_ & ~pstart_0_ & pencrypt_0_;
  assign n1825 = ~n1328 & pksi_82_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1826 = n1327_1 & pksi_75_ & ~pstart_0_ & pencrypt_0_;
  assign n1827 = n1328 & n_n2272 & ~pstart_0_ & ~pencrypt_0_;
  assign n1828 = ~n1328 & pksi_102_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1829 = n1328 & pksi_98_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1830 = ~n1327_1 & pksi_112_ & ~pstart_0_ & pencrypt_0_;
  assign n1831 = ~n1328 & pksi_110_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1832 = n1327_1 & pksi_115_ & ~pstart_0_ & pencrypt_0_;
  assign n1833 = n1328 & pksi_103_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1834 = ~n1328 & pksi_107_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1835 = n1328 & pksi_109_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1836 = ~n1327_1 & pksi_97_ & ~pstart_0_ & pencrypt_0_;
  assign n1837 = ~n1328 & pksi_189_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1838 = n1328 & pksi_171_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1839 = ~n1327_1 & pksi_175_ & ~pstart_0_ & pencrypt_0_;
  assign n1840 = ~n1328 & pksi_177_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1841 = n1328 & pksi_186_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1842 = ~n1327_1 & n_n109 & ~pstart_0_ & pencrypt_0_;
  assign n1843 = ~n1328 & n_n2396 & ~pstart_0_ & ~pencrypt_0_;
  assign n1844 = n1328 & pksi_173_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1845 = ~n1327_1 & pksi_102_ & ~pstart_0_ & pencrypt_0_;
  assign n1846 = ~n1328 & pksi_19_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1847 = n1328 & pksi_17_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1848 = ~n1327_1 & pksi_2_ & ~pstart_0_ & pencrypt_0_;
  assign n1849 = ~n1328 & n_n2513 & ~pstart_0_ & ~pencrypt_0_;
  assign n1850 = n1328 & pksi_110_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1851 = ~n1327_1 & pksi_115_ & ~pstart_0_ & pencrypt_0_;
  assign n1852 = ~n1328 & pksi_109_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1853 = n1328 & pksi_116_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1854 = ~n1327_1 & pksi_113_ & ~pstart_0_ & pencrypt_0_;
  assign n1855 = ~n1328 & n_n2420 & ~pstart_0_ & ~pencrypt_0_;
  assign n1856 = n1328 & pksi_189_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1857 = ~n1327_1 & pksi_182_ & ~pstart_0_ & pencrypt_0_;
  assign n1858 = ~n1328 & pksi_186_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1859 = n1328 & pksi_172_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1860 = ~n1327_1 & pksi_188_ & ~pstart_0_ & pencrypt_0_;
  assign n1861 = ~n1328 & pksi_185_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1862 = n1328 & n_n2396 & ~pstart_0_ & ~pencrypt_0_;
  assign n1863 = ~n1327_1 & pksi_118_ & ~pstart_0_ & pencrypt_0_;
  assign n1864 = ~n1328 & pksi_17_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1865 = n1328 & n_n2384 & ~pstart_0_ & ~pencrypt_0_;
  assign n1866 = ~n1327_1 & pksi_14_ & ~pstart_0_ & pencrypt_0_;
  assign n1867 = ~n1328 & pksi_183_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1868 = n1328 & pksi_118_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1869 = ~n1327_1 & pksi_119_ & ~pstart_0_ & pencrypt_0_;
  assign n1870 = ~n1328 & pksi_116_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1871 = ~n1327_1 & n_n2495 & ~pstart_0_ & pencrypt_0_;
  assign n1872 = n1328 & pksi_104_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1873 = ~n1328 & pksi_97_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1874 = n1328 & pksi_113_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1875 = ~n1327_1 & pksi_111_ & ~pstart_0_ & pencrypt_0_;
  assign n1876 = ~n1328 & pksi_130_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1877 = n1328 & pksi_136_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1878 = ~n1327_1 & pksi_123_ & ~pstart_0_ & pencrypt_0_;
  assign n1879 = ~n1328 & pksi_184_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1880 = ~n1327_1 & n_n2416 & ~pstart_0_ & pencrypt_0_;
  assign n1881 = n1328 & n_n2420 & ~pstart_0_ & ~pencrypt_0_;
  assign n1882 = ~n1328 & n_n2408 & ~pstart_0_ & ~pencrypt_0_;
  assign n1883 = n1328 & pksi_180_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1884 = ~n1327_1 & pksi_172_ & ~pstart_0_ & pencrypt_0_;
  assign n1885 = ~n1328 & pksi_79_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1886 = n1328 & pksi_4_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1887 = ~n1327_1 & pksi_15_ & ~pstart_0_ & pencrypt_0_;
  assign n1888 = ~n1328 & n_n2384 & ~pstart_0_ & ~pencrypt_0_;
  assign n1889 = n1328 & pksi_11_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1890 = ~n1327_1 & pksi_22_ & ~pstart_0_ & pencrypt_0_;
  assign n1891 = ~n1328 & pksi_118_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1892 = n1328 & pksi_102_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1893 = ~n1327_1 & pksi_106_ & ~pstart_0_ & pencrypt_0_;
  assign n1894 = ~n1328 & pksi_103_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1895 = n1328 & pksi_96_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1896 = ~n1327_1 & pksi_108_ & ~pstart_0_ & pencrypt_0_;
  assign n1897 = ~n1328 & pksi_104_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1898 = n1328 & pksi_97_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1899 = ~n1327_1 & pksi_101_ & ~pstart_0_ & pencrypt_0_;
  assign n1900 = ~n1328 & pksi_136_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1901 = n1327_1 & pksi_123_ & ~pstart_0_ & pencrypt_0_;
  assign n1902 = n1328 & n_n2485 & ~pstart_0_ & ~pencrypt_0_;
  assign n1903 = ~n1328 & pksi_178_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1904 = n1328 & pksi_184_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1905 = ~n1327_1 & pksi_171_ & ~pstart_0_ & pencrypt_0_;
  assign n1906 = ~n1328 & pksi_180_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1907 = n1328 & pksi_177_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1908 = ~n1327_1 & pksi_179_ & ~pstart_0_ & pencrypt_0_;
  assign n1909 = ~n1328 & pksi_92_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1910 = n1328 & pksi_79_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1911 = ~n1327_1 & pksi_6_ & ~pstart_0_ & pencrypt_0_;
  assign n1912 = ~n1328 & pksi_11_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1913 = n1328 & pksi_2_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1914 = ~n1327_1 & pksi_0_ & ~pstart_0_ & pencrypt_0_;
  assign n1915 = n1328 & n_n2277 & ~pstart_0_ & ~pencrypt_0_;
  assign n1916 = ~n1328 & pksi_73_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1917 = ~n1327_1 & pksi_82_ & ~pstart_0_ & pencrypt_0_;
  assign n1918 = ~n1328 & n_n2517 & ~pstart_0_ & ~pencrypt_0_;
  assign n1919 = n1328 & pksi_117_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1920 = ~n1327_1 & pksi_110_ & ~pstart_0_ & pencrypt_0_;
  assign n1921 = ~n1328 & pksi_108_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1922 = n1328 & pksi_105_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1923 = ~n1327_1 & pksi_107_ & ~pstart_0_ & pencrypt_0_;
  assign n1924 = ~n1328 & pksi_132_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1925 = n1328 & pksi_129_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1926 = ~n1327_1 & pksi_131_ & ~pstart_0_ & pencrypt_0_;
  assign n1927 = n1328 & n_n2462 & ~pstart_0_ & ~pencrypt_0_;
  assign n1928 = ~n1328 & pksi_137_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1929 = ~n1327_1 & pksi_166_ & ~pstart_0_ & pencrypt_0_;
  assign n1930 = ~n1328 & n_n121 & ~pstart_0_ & ~pencrypt_0_;
  assign n1931 = n1328 & pksi_178_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1932 = ~n1327_1 & pksi_189_ & ~pstart_0_ & pencrypt_0_;
  assign n1933 = ~n1328 & n_n2412 & ~pstart_0_ & ~pencrypt_0_;
  assign n1934 = n1328 & n_n2410 & ~pstart_0_ & ~pencrypt_0_;
  assign n1935 = ~n1327_1 & pksi_177_ & ~pstart_0_ & pencrypt_0_;
  assign n1936 = ~n1328 & pksi_188_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1937 = n1328 & pksi_176_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1938 = ~n1327_1 & n_n2396 & ~pstart_0_ & pencrypt_0_;
  assign n1939 = ~n1328 & pksi_6_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1940 = n1328 & pksi_15_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1941 = ~n1327_1 & pksi_19_ & ~pstart_0_ & pencrypt_0_;
  assign n1942 = ~n1328 & pksi_173_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1943 = n1328 & pksi_183_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1944 = ~n1327_1 & pksi_98_ & ~pstart_0_ & pencrypt_0_;
  assign n1945 = ~n1328 & pksi_112_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1946 = n1328 & n_n2517 & ~pstart_0_ & ~pencrypt_0_;
  assign n1947 = ~n1327_1 & n_n2513 & ~pstart_0_ & pencrypt_0_;
  assign n1948 = ~n1328 & pksi_105_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1949 = n1328 & pksi_114_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1950 = ~n1327_1 & pksi_109_ & ~pstart_0_ & pencrypt_0_;
  assign n1951 = ~n1328 & n_n2474 & ~pstart_0_ & ~pencrypt_0_;
  assign n1952 = n1328 & pksi_132_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1953 = ~n1327_1 & pksi_124_ & ~pstart_0_ & pencrypt_0_;
  assign n1954 = ~n1328 & n_n2462 & ~pstart_0_ & ~pencrypt_0_;
  assign n1955 = n1328 & pksi_125_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1956 = ~n1327_1 & pksi_150_ & ~pstart_0_ & pencrypt_0_;
  assign n1957 = ~n1328 & pksi_170_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1958 = ~n1327_1 & n_n2420 & ~pstart_0_ & pencrypt_0_;
  assign n1959 = n1328 & n_n121 & ~pstart_0_ & ~pencrypt_0_;
  assign n1960 = ~n1328 & n_n2410 & ~pstart_0_ & ~pencrypt_0_;
  assign n1961 = n1328 & n_n2408 & ~pstart_0_ & ~pencrypt_0_;
  assign n1962 = ~n1327_1 & pksi_186_ & ~pstart_0_ & pencrypt_0_;
  assign n1963 = ~n1328 & n_n109 & ~pstart_0_ & ~pencrypt_0_;
  assign n1964 = n1328 & pksi_188_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1965 = ~n1327_1 & pksi_185_ & ~pstart_0_ & pencrypt_0_;
  assign n1966 = ~n1328 & pksi_15_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1967 = n1328 & pksi_5_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1968 = ~n1327_1 & pksi_17_ & ~pstart_0_ & pencrypt_0_;
  assign n1969 = ~n1328 & pksi_99_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1970 = n1328 & n_n2513 & ~pstart_0_ & ~pencrypt_0_;
  assign n1971 = ~n1327_1 & pksi_96_ & ~pstart_0_ & pencrypt_0_;
  assign n1972 = ~n1328 & pksi_114_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1973 = n1328 & pksi_100_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1974 = ~n1327_1 & pksi_116_ & ~pstart_0_ & pencrypt_0_;
  assign n1975 = ~n1328 & pksi_165_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1976 = n1328 & pksi_147_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1977 = ~n1327_1 & pksi_151_ & ~pstart_0_ & pencrypt_0_;
  assign n1978 = ~n1328 & n_n2440 & ~pstart_0_ & ~pencrypt_0_;
  assign n1979 = n1328 & pksi_162_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1980 = ~n1327_1 & pksi_157_ & ~pstart_0_ & pencrypt_0_;
  assign n1981 = ~n1328 & pksi_174_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1982 = n1328 & pksi_170_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1983 = ~n1327_1 & pksi_184_ & ~pstart_0_ & pencrypt_0_;
  assign n1984 = ~n1328 & pksi_182_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1985 = ~n1327_1 & n_n2408 & ~pstart_0_ & pencrypt_0_;
  assign n1986 = n1328 & pksi_175_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1987 = ~n1328 & pksi_169_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1988 = n1328 & pksi_185_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1989 = ~n1327_1 & pksi_183_ & ~pstart_0_ & pencrypt_0_;
  assign n1990 = ~n1328 & pksi_5_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1991 = ~n1327_1 & n_n2384 & ~pstart_0_ & pencrypt_0_;
  assign n1992 = n1328 & pksi_9_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1993 = ~n1328 & pksi_117_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1994 = n1328 & pksi_99_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1995 = ~n1327_1 & pksi_103_ & ~pstart_0_ & pencrypt_0_;
  assign n1996 = ~n1328 & pksi_100_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1997 = n1328 & pksi_107_ & ~pstart_0_ & ~pencrypt_0_;
  assign n1998 = ~n1327_1 & pksi_104_ & ~pstart_0_ & pencrypt_0_;
  assign n1999 = ~n1328 & n_n2452 & ~pstart_0_ & ~pencrypt_0_;
  assign n2000 = n1328 & pksi_165_ & ~pstart_0_ & ~pencrypt_0_;
  assign n2001 = ~n1327_1 & pksi_158_ & ~pstart_0_ & pencrypt_0_;
  assign n2002 = ~n1328 & pksi_162_ & ~pstart_0_ & ~pencrypt_0_;
  assign n2003 = n1328 & pksi_148_ & ~pstart_0_ & ~pencrypt_0_;
  assign n2004 = ~n1327_1 & pksi_164_ & ~pstart_0_ & pencrypt_0_;
  assign n2005 = ~n1328 & pksi_190_ & ~pstart_0_ & ~pencrypt_0_;
  assign n2006 = n1328 & pksi_174_ & ~pstart_0_ & ~pencrypt_0_;
  assign n2007 = ~n1327_1 & pksi_178_ & ~pstart_0_ & pencrypt_0_;
  assign n2008 = ~n1328 & pksi_175_ & ~pstart_0_ & ~pencrypt_0_;
  assign n2009 = n1328 & n_n2412 & ~pstart_0_ & ~pencrypt_0_;
  assign n2010 = ~n1327_1 & pksi_180_ & ~pstart_0_ & pencrypt_0_;
  assign n2011 = ~n1328 & pksi_176_ & ~pstart_0_ & ~pencrypt_0_;
  assign n2012 = n1328 & pksi_169_ & ~pstart_0_ & ~pencrypt_0_;
  assign n2013 = ~n1327_1 & pksi_173_ & ~pstart_0_ & pencrypt_0_;
  assign n2014 = ~n1328 & pksi_9_ & ~pstart_0_ & ~pencrypt_0_;
  assign n2015 = n1328 & pksi_19_ & ~pstart_0_ & ~pencrypt_0_;
  assign n2016 = ~n1327_1 & pksi_11_ & ~pstart_0_ & pencrypt_0_;
  assign n2017 = pstart_0_ & (pencrypt_0_ ? pkey_57_ : pkey_0_);
  assign n2018 = n2017 | (n_n2384 & n1327_1 & n1332_1);
  assign n2019 = pstart_0_ & (pencrypt_0_ ? pkey_211_ : pkey_219_);
  assign n2020 = n2019 | (n_n2396 & n1327_1 & n1332_1);
  assign n2021 = pstart_0_ & (pencrypt_0_ ? pkey_205_ : pkey_213_);
  assign n2022 = n2021 | (n_n2408 & n1327_1 & n1332_1);
  assign n2023 = pstart_0_ & (pencrypt_0_ ? pkey_230_ : pkey_238_);
  assign n2024 = n2023 | (n_n121 & n1327_1 & n1332_1);
  assign n2025 = pstart_0_ & (pencrypt_0_ ? pkey_156_ : pkey_164_);
  assign n2026 = n2025 | (pksi_157_ & n1327_1 & n1332_1);
  assign n2027 = pstart_0_ & (pencrypt_0_ ? pkey_181_ : pkey_189_);
  assign n2028 = n2027 | (n_n2448 & n1327_1 & n1332_1);
  assign n2029 = pstart_0_ & (pencrypt_0_ ? pkey_20_ : pkey_28_);
  assign n2030 = n2029 | (pksi_116_ & n1327_1 & n1332_1);
  assign n2031 = pstart_0_ & (pencrypt_0_ ? pkey_45_ : pkey_53_);
  assign n2032 = n2031 | (pksi_110_ & n1327_1 & n1332_1);
  assign n2033 = pstart_0_ & (pencrypt_0_ ? pkey_0_ : pkey_8_);
  assign n2034 = n2033 | (pksi_17_ & n1327_1 & n1332_1);
  assign n2035 = pstart_0_ & (pencrypt_0_ ? pkey_203_ : pkey_211_);
  assign n2036 = n2035 | (pksi_173_ & n1327_1 & n1332_1);
  assign n2037 = pstart_0_ & (pencrypt_0_ ? pkey_213_ : pkey_221_);
  assign n2038 = n2037 | (n_n2410 & n1327_1 & n1332_1);
  assign n2039 = pstart_0_ & (pencrypt_0_ ? pkey_222_ : pkey_230_);
  assign n2040 = n2039 | (pksi_178_ & n1327_1 & n1332_1);
  assign n2041 = pstart_0_ & (pencrypt_0_ ? pkey_164_ : pkey_172_);
  assign n2042 = n2041 | (pksi_155_ & n1327_1 & n1332_1);
  assign n2043 = pstart_0_ & (pencrypt_0_ ? pkey_173_ : pkey_181_);
  assign n2044 = n2043 | (pksi_158_ & n1327_1 & n1332_1);
  assign n2045 = pstart_0_ & (pencrypt_0_ ? pkey_28_ : pkey_36_);
  assign n2046 = n2045 | (pksi_109_ & n1327_1 & n1332_1);
  assign n2047 = pstart_0_ & (pencrypt_0_ ? pkey_37_ : pkey_45_);
  assign n2048 = n2047 | (pksi_103_ & n1327_1 & n1332_1);
  assign n2049 = pstart_0_ & (pencrypt_0_ ? pkey_8_ : pkey_16_);
  assign n2050 = n2049 | (pksi_19_ & n1327_1 & n1332_1);
  assign n2051 = pstart_0_ & (pencrypt_0_ ? pkey_196_ : pkey_204_);
  assign n2052 = n2051 | (pksi_169_ & n1327_1 & n1332_1);
  assign n2053 = pstart_0_ & (pencrypt_0_ ? pkey_252_ : pkey_197_);
  assign n2054 = n2053 | (pksi_177_ & n1327_1 & n1332_1);
  assign n2055 = pstart_0_ & (pencrypt_0_ ? pkey_214_ : pkey_222_);
  assign n2056 = n2055 | (pksi_184_ & n1327_1 & n1332_1);
  assign n2057 = pstart_0_ & (pencrypt_0_ ? pkey_190_ : pkey_67_);
  assign n2058 = n2057 | (pksi_166_ & n1327_1 & n1332_1);
  assign n2059 = pstart_0_ & (pencrypt_0_ ? pkey_116_ : pkey_124_);
  assign n2060 = n2059 | (pksi_138_ & n1327_1 & n1332_1);
  assign n2061 = pstart_0_ & (pencrypt_0_ ? pkey_36_ : pkey_44_);
  assign n2062 = n2061 | (pksi_107_ & n1327_1 & n1332_1);
  assign n2063 = pstart_0_ & (pencrypt_0_ ? pkey_61_ : pkey_6_);
  assign n2064 = n2063 | (pksi_99_ & n1327_1 & n1332_1);
  assign n2065 = pstart_0_ & (pencrypt_0_ ? pkey_54_ : pkey_62_);
  assign n2066 = n2065 | (pksi_102_ & n1327_1 & n1332_1);
  assign n2067 = pstart_0_ & (pencrypt_0_ ? pkey_16_ : pkey_24_);
  assign n2068 = n2067 | (pksi_9_ & n1327_1 & n1332_1);
  assign n2069 = pstart_0_ & (pencrypt_0_ ? pkey_219_ : pkey_196_);
  assign n2070 = n2069 | (pksi_185_ & n1327_1 & n1332_1);
  assign n2071 = pstart_0_ & (pencrypt_0_ ? pkey_197_ : pkey_205_);
  assign n2072 = n2071 | (pksi_180_ & n1327_1 & n1332_1);
  assign n2073 = pstart_0_ & (pencrypt_0_ ? pkey_206_ : pkey_214_);
  assign n2074 = n2073 | (n_n2420 & n1327_1 & n1332_1);
  assign n2075 = pstart_0_ & (pencrypt_0_ ? pkey_67_ : pkey_75_);
  assign n2076 = n2075 | (pksi_135_ & n1327_1 & n1332_1);
  assign n2077 = pstart_0_ & (pencrypt_0_ ? pkey_44_ : pkey_116_);
  assign n2078 = n2077 | (pksi_124_ & n1327_1 & n1332_1);
  assign n2079 = pstart_0_ & (pencrypt_0_ ? pkey_44_ : pkey_52_);
  assign n2080 = n2079 | (pksi_100_ & n1327_1 & n1332_1);
  assign n2081 = pstart_0_ & (pencrypt_0_ ? pkey_53_ : pkey_61_);
  assign n2082 = n2081 | (n_n2513 & n1327_1 & n1332_1);
  assign n2083 = pstart_0_ & (pencrypt_0_ ? pkey_226_ : pkey_234_);
  assign n2084 = n2083 | (pksi_93_ & n1327_1 & n1332_1);
  assign n2085 = pstart_0_ & (pencrypt_0_ ? pkey_25_ : pkey_33_);
  assign n2086 = n2085 | (pksi_22_ & n1327_1 & n1332_1);
  assign n2087 = pstart_0_ & (pencrypt_0_ ? pkey_48_ : pkey_56_);
  assign n2088 = n2087 | (pksi_23_ & n1327_1 & n1332_1);
  assign n2089 = pstart_0_ & (pencrypt_0_ ? pkey_172_ : pkey_244_);
  assign n2090 = n2089 | (pksi_172_ & n1327_1 & n1332_1);
  assign n2091 = pstart_0_ & (pencrypt_0_ ? pkey_198_ : pkey_206_);
  assign n2092 = n2091 | (pksi_189_ & n1327_1 & n1332_1);
  assign n2093 = pstart_0_ & (pencrypt_0_ ? pkey_125_ : pkey_70_);
  assign n2094 = n2093 | (n_n2481 & ~n1327_1 & n1332_1);
  assign n2095 = pstart_0_ & (pencrypt_0_ ? pkey_19_ : pkey_27_);
  assign n2096 = n2095 | (n_n2495 & n1327_1 & n1332_1);
  assign n2097 = pstart_0_ & (pencrypt_0_ ? pkey_13_ : pkey_21_);
  assign n2098 = n2097 | (n_n2507 & n1327_1 & n1332_1);
  assign n2099 = pstart_0_ & (pencrypt_0_ ? pkey_38_ : pkey_46_);
  assign n2100 = n2099 | (pksi_119_ & n1327_1 & n1332_1);
  assign n2101 = pstart_0_ & (pencrypt_0_ ? pkey_33_ : pkey_41_);
  assign n2102 = n2101 | (pksi_14_ & n1327_1 & n1332_1);
  assign n2103 = pstart_0_ & (pencrypt_0_ ? pkey_40_ : pkey_48_);
  assign n2104 = n2103 | (pksi_6_ & n1327_1 & n1332_1);
  assign n2105 = pstart_0_ & (pencrypt_0_ ? pkey_244_ : pkey_252_);
  assign n2106 = n2105 | (pksi_186_ & n1327_1 & n1332_1);
  assign n2107 = pstart_0_ & (pencrypt_0_ ? pkey_253_ : pkey_198_);
  assign n2108 = n2107 | (pksi_171_ & n1327_1 & n1332_1);
  assign n2109 = pstart_0_ & (pencrypt_0_ ? pkey_70_ : pkey_78_);
  assign n2110 = n2109 | (pksi_141_ & n1327_1 & n1332_1);
  assign n2111 = pstart_0_ & (pencrypt_0_ ? pkey_11_ : pkey_19_);
  assign n2112 = n2111 | (pksi_101_ & n1327_1 & n1332_1);
  assign n2113 = pstart_0_ & (pencrypt_0_ ? pkey_27_ : pkey_4_);
  assign n2114 = n2113 | (pksi_113_ & n1327_1 & n1332_1);
  assign n2115 = pstart_0_ & (pencrypt_0_ ? pkey_46_ : pkey_54_);
  assign n2116 = n2115 | (pksi_98_ & n1327_1 & n1332_1);
  assign n2117 = pstart_0_ & (pencrypt_0_ ? pkey_41_ : pkey_49_);
  assign n2118 = n2117 | (pksi_2_ & n1327_1 & n1332_1);
  assign n2119 = pstart_0_ & (pencrypt_0_ ? pkey_195_ : pkey_203_);
  assign n2120 = n2119 | (pksi_183_ & n1327_1 & n1332_1);
  assign n2121 = pstart_0_ & (pencrypt_0_ ? pkey_220_ : pkey_228_);
  assign n2122 = n2121 | (n_n109 & n1327_1 & n1332_1);
  assign n2123 = pstart_0_ & (pencrypt_0_ ? pkey_245_ : pkey_253_);
  assign n2124 = n2123 | (n_n2416 & n1327_1 & n1332_1);
  assign n2125 = pstart_0_ & (pencrypt_0_ ? pkey_4_ : pkey_12_);
  assign n2126 = n2125 | (pksi_97_ & n1327_1 & n1332_1);
  assign n2127 = pstart_0_ & (pencrypt_0_ ? pkey_29_ : pkey_37_);
  assign n2128 = n2127 | (pksi_96_ & n1327_1 & n1332_1);
  assign n2129 = pstart_0_ & (pencrypt_0_ ? pkey_49_ : pkey_57_);
  assign n2130 = n2129 | (pksi_11_ & n1327_1 & n1332_1);
  assign n2131 = pstart_0_ & (pencrypt_0_ ? pkey_62_ : pkey_195_);
  assign n2132 = n2131 | (pksi_118_ & n1327_1 & n1332_1);
  assign n2133 = pstart_0_ & (pencrypt_0_ ? pkey_228_ : pkey_172_);
  assign n2134 = n2133 | (pksi_179_ & n1327_1 & n1332_1);
  assign n2135 = pstart_0_ & (pencrypt_0_ ? pkey_237_ : pkey_245_);
  assign n2136 = n2135 | (pksi_182_ & n1327_1 & n1332_1);
  assign n2137 = pstart_0_ & (pencrypt_0_ ? pkey_12_ : pkey_20_);
  assign n2138 = n2137 | (pksi_104_ & n1327_1 & n1332_1);
  assign n2139 = pstart_0_ & (pencrypt_0_ ? pkey_21_ : pkey_29_);
  assign n2140 = n2139 | (n_n2507 & ~n1327_1 & n1332_1);
  assign n2141 = pstart_0_ & (pencrypt_0_ ? pkey_30_ : pkey_38_);
  assign n2142 = n2141 | (pksi_106_ & n1327_1 & n1332_1);
  assign n2143 = pstart_0_ & (pencrypt_0_ ? pkey_194_ : pkey_202_);
  assign n2144 = n2143 | (n_n2268 & ~n1327_1 & n1332_1);
  assign n2145 = pstart_0_ & (pencrypt_0_ ? pkey_254_ : pkey_131_);
  assign n2146 = n2145 | (pksi_190_ & n1327_1 & n1332_1);
  assign n2147 = pstart_0_ & (pencrypt_0_ ? pkey_180_ : pkey_188_);
  assign n2148 = n2147 | (pksi_162_ & n1327_1 & n1332_1);
  assign n2149 = pstart_0_ & (pencrypt_0_ ? pkey_142_ : pkey_150_);
  assign n2150 = n2149 | (n_n2452 & n1327_1 & n1332_1);
  assign n2151 = pstart_0_ & (pencrypt_0_ ? pkey_68_ : pkey_76_);
  assign n2152 = n2151 | (pksi_121_ & n1327_1 & n1332_1);
  assign n2153 = pstart_0_ & (pencrypt_0_ ? pkey_93_ : pkey_101_);
  assign n2154 = n2153 | (n_n2476 & ~n1327_1 & n1332_1);
  assign n2155 = pstart_0_ & (pencrypt_0_ ? pkey_118_ : pkey_126_);
  assign n2156 = n2155 | (pksi_126_ & n1327_1 & n1332_1);
  assign n2157 = pstart_0_ & (pencrypt_0_ ? pkey_202_ : pkey_210_);
  assign n2158 = n2157 | (pksi_84_ & n1327_1 & n1332_1);
  assign n2159 = pstart_0_ & (pencrypt_0_ ? pkey_131_ : pkey_139_);
  assign n2160 = n2159 | (pksi_159_ & n1327_1 & n1332_1);
  assign n2161 = pstart_0_ & (pencrypt_0_ ? pkey_172_ : pkey_180_);
  assign n2162 = n2161 | (pksi_148_ & n1327_1 & n1332_1);
  assign n2163 = pstart_0_ & (pencrypt_0_ ? pkey_150_ : pkey_158_);
  assign n2164 = n2163 | (n_n2452 & ~n1327_1 & n1332_1);
  assign n2165 = pstart_0_ & (pencrypt_0_ ? pkey_91_ : pkey_68_);
  assign n2166 = n2165 | (n_n2462 & ~n1327_1 & n1332_1);
  assign n2167 = pstart_0_ & (pencrypt_0_ ? pkey_101_ : pkey_109_);
  assign n2168 = n2167 | (pksi_127_ & n1327_1 & n1332_1);
  assign n2169 = pstart_0_ & (pencrypt_0_ ? pkey_110_ : pkey_118_);
  assign n2170 = n2169 | (pksi_122_ & n1327_1 & n1332_1);
  assign n2171 = pstart_0_ & (pencrypt_0_ ? pkey_210_ : pkey_218_);
  assign n2172 = n2171 | (n_n2272 & n1327_1 & n1332_1);
  assign n2173 = pstart_0_ & (pencrypt_0_ ? pkey_139_ : pkey_147_);
  assign n2174 = n2173 | (pksi_149_ & n1327_1 & n1332_1);
  assign n2175 = pstart_0_ & (pencrypt_0_ ? pkey_133_ : pkey_141_);
  assign n2176 = n2175 | (pksi_156_ & n1327_1 & n1332_1);
  assign n2177 = pstart_0_ & (pencrypt_0_ ? pkey_189_ : pkey_134_);
  assign n2178 = n2177 | (pksi_147_ & n1327_1 & n1332_1);
  assign n2179 = pstart_0_ & (pencrypt_0_ ? pkey_83_ : pkey_91_);
  assign n2180 = n2179 | (n_n2462 & n1327_1 & n1332_1);
  assign n2181 = pstart_0_ & (pencrypt_0_ ? pkey_109_ : pkey_117_);
  assign n2182 = n2181 | (pksi_134_ & n1327_1 & n1332_1);
  assign n2183 = pstart_0_ & (pencrypt_0_ ? pkey_3_ : pkey_11_);
  assign n2184 = n2183 | (pksi_111_ & n1327_1 & n1332_1);
  assign n2185 = pstart_0_ & (pencrypt_0_ ? pkey_218_ : pkey_226_);
  assign n2186 = n2185 | (pksi_82_ & n1327_1 & n1332_1);
  assign n2187 = pstart_0_ & (pencrypt_0_ ? pkey_147_ : pkey_155_);
  assign n2188 = n2187 | (n_n2430 & n1327_1 & n1332_1);
  assign n2189 = pstart_0_ & (pencrypt_0_ ? pkey_188_ : pkey_133_);
  assign n2190 = n2189 | (n_n2440 & n1327_1 & n1332_1);
  assign n2191 = pstart_0_ & (pencrypt_0_ ? pkey_134_ : pkey_142_);
  assign n2192 = n2191 | (pksi_165_ & n1327_1 & n1332_1);
  assign n2193 = pstart_0_ & (pencrypt_0_ ? pkey_75_ : pkey_83_);
  assign n2194 = n2193 | (pksi_125_ & n1327_1 & n1332_1);
  assign n2195 = pstart_0_ & (pencrypt_0_ ? pkey_117_ : pkey_125_);
  assign n2196 = n2195 | (n_n2481 & n1327_1 & n1332_1);
  assign n2197 = pstart_0_ & (pencrypt_0_ ? pkey_126_ : pkey_3_);
  assign n2198 = n2197 | (pksi_142_ & n1327_1 & n1332_1);
  assign n2199 = pstart_0_ & (pencrypt_0_ ? pkey_227_ : pkey_235_);
  assign n2200 = n2199 | (pksi_79_ & n1327_1 & n1332_1);
  assign n2201 = pstart_0_ & (pencrypt_0_ ? pkey_24_ : pkey_32_);
  assign n2202 = n2201 | (pksi_5_ & n1327_1 & n1332_1);
  assign n2203 = pstart_0_ & (pencrypt_0_ ? pkey_212_ : pkey_220_);
  assign n2204 = n2203 | (pksi_188_ & n1327_1 & n1332_1);
  assign n2205 = pstart_0_ & (pencrypt_0_ ? pkey_155_ : pkey_132_);
  assign n2206 = n2205 | (n_n2430 & ~n1327_1 & n1332_1);
  assign n2207 = pstart_0_ & (pencrypt_0_ ? pkey_149_ : pkey_157_);
  assign n2208 = n2207 | (pksi_163_ & n1327_1 & n1332_1);
  assign n2209 = pstart_0_ & (pencrypt_0_ ? pkey_174_ : pkey_182_);
  assign n2210 = n2209 | (pksi_146_ & n1327_1 & n1332_1);
  assign n2211 = pstart_0_ & (pencrypt_0_ ? pkey_100_ : pkey_44_);
  assign n2212 = n2211 | (pksi_131_ & n1327_1 & n1332_1);
  assign n2213 = pstart_0_ & (pencrypt_0_ ? pkey_124_ : pkey_69_);
  assign n2214 = n2213 | (pksi_129_ & n1327_1 & n1332_1);
  assign n2215 = pstart_0_ & (pencrypt_0_ ? pkey_86_ : pkey_94_);
  assign n2216 = n2215 | (pksi_136_ & n1327_1 & n1332_1);
  assign n2217 = pstart_0_ & (pencrypt_0_ ? pkey_52_ : pkey_60_);
  assign n2218 = n2217 | (pksi_114_ & n1327_1 & n1332_1);
  assign n2219 = pstart_0_ & (pencrypt_0_ ? pkey_14_ : pkey_22_);
  assign n2220 = n2219 | (n_n2517 & n1327_1 & n1332_1);
  assign n2221 = pstart_0_ & (pencrypt_0_ ? pkey_235_ : pkey_243_);
  assign n2222 = n2221 | (pksi_92_ & n1327_1 & n1332_1);
  assign n2223 = pstart_0_ & (pencrypt_0_ ? pkey_32_ : pkey_40_);
  assign n2224 = n2223 | (pksi_15_ & n1327_1 & n1332_1);
  assign n2225 = pstart_0_ & (pencrypt_0_ ? pkey_204_ : pkey_212_);
  assign n2226 = n2225 | (pksi_176_ & n1327_1 & n1332_1);
  assign n2227 = pstart_0_ & (pencrypt_0_ ? pkey_132_ : pkey_140_);
  assign n2228 = n2227 | (pksi_145_ & n1327_1 & n1332_1);
  assign n2229 = pstart_0_ & (pencrypt_0_ ? pkey_141_ : pkey_149_);
  assign n2230 = n2229 | (pksi_153_ & n1327_1 & n1332_1);
  assign n2231 = pstart_0_ & (pencrypt_0_ ? pkey_182_ : pkey_190_);
  assign n2232 = n2231 | (pksi_150_ & n1327_1 & n1332_1);
  assign n2233 = pstart_0_ & (pencrypt_0_ ? pkey_92_ : pkey_100_);
  assign n2234 = n2233 | (pksi_133_ & n1327_1 & n1332_1);
  assign n2235 = pstart_0_ & (pencrypt_0_ ? pkey_69_ : pkey_77_);
  assign n2236 = n2235 | (pksi_132_ & n1327_1 & n1332_1);
  assign n2237 = pstart_0_ & (pencrypt_0_ ? pkey_78_ : pkey_86_);
  assign n2238 = n2237 | (n_n2485 & n1327_1 & n1332_1);
  assign n2239 = pstart_0_ & (pencrypt_0_ ? pkey_60_ : pkey_5_);
  assign n2240 = n2239 | (pksi_105_ & n1327_1 & n1332_1);
  assign n2241 = pstart_0_ & (pencrypt_0_ ? pkey_6_ : pkey_14_);
  assign n2242 = n2241 | (pksi_117_ & n1327_1 & n1332_1);
  assign n2243 = pstart_0_ & (pencrypt_0_ ? pkey_243_ : pkey_251_);
  assign n2244 = n2243 | (n_n10 & n1327_1 & n1332_1);
  assign n2245 = pstart_0_ & (pencrypt_0_ ? pkey_221_ : pkey_229_);
  assign n2246 = n2245 | (n_n2412 & n1327_1 & n1332_1);
  assign n2247 = pstart_0_ & (pencrypt_0_ ? pkey_246_ : pkey_254_);
  assign n2248 = n2247 | (pksi_174_ & n1327_1 & n1332_1);
  assign n2249 = pstart_0_ & (pencrypt_0_ ? pkey_140_ : pkey_148_);
  assign n2250 = n2249 | (pksi_152_ & n1327_1 & n1332_1);
  assign n2251 = pstart_0_ & (pencrypt_0_ ? pkey_165_ : pkey_173_);
  assign n2252 = n2251 | (pksi_151_ & n1327_1 & n1332_1);
  assign n2253 = pstart_0_ & (pencrypt_0_ ? pkey_158_ : pkey_166_);
  assign n2254 = n2253 | (pksi_154_ & n1327_1 & n1332_1);
  assign n2255 = pstart_0_ & (pencrypt_0_ ? pkey_84_ : pkey_92_);
  assign n2256 = n2255 | (pksi_140_ & n1327_1 & n1332_1);
  assign n2257 = pstart_0_ & (pencrypt_0_ ? pkey_77_ : pkey_85_);
  assign n2258 = n2257 | (n_n2474 & n1327_1 & n1332_1);
  assign n2259 = pstart_0_ & (pencrypt_0_ ? pkey_102_ : pkey_110_);
  assign n2260 = n2259 | (n_n168 & n1327_1 & n1332_1);
  assign n2261 = pstart_0_ & (pencrypt_0_ ? pkey_5_ : pkey_13_);
  assign n2262 = n2261 | (pksi_108_ & n1327_1 & n1332_1);
  assign n2263 = pstart_0_ & (pencrypt_0_ ? pkey_251_ : pkey_194_);
  assign n2264 = n2263 | (n_n2268 & n1327_1 & n1332_1);
  assign n2265 = pstart_0_ & (pencrypt_0_ ? pkey_229_ : pkey_237_);
  assign n2266 = n2265 | (pksi_175_ & n1327_1 & n1332_1);
  assign n2267 = pstart_0_ & (pencrypt_0_ ? pkey_238_ : pkey_246_);
  assign n2268 = n2267 | (pksi_170_ & n1327_1 & n1332_1);
  assign n2269 = pstart_0_ & (pencrypt_0_ ? pkey_148_ : pkey_156_);
  assign n2270 = n2269 | (pksi_164_ & n1327_1 & n1332_1);
  assign n2271 = pstart_0_ & (pencrypt_0_ ? pkey_157_ : pkey_165_);
  assign n2272 = n2271 | (pksi_144_ & n1327_1 & n1332_1);
  assign n2273 = pstart_0_ & (pencrypt_0_ ? pkey_166_ : pkey_174_);
  assign n2274 = n2273 | (pksi_167_ & n1327_1 & n1332_1);
  assign n2275 = pstart_0_ & (pencrypt_0_ ? pkey_76_ : pkey_84_);
  assign n2276 = n2275 | (pksi_128_ & n1327_1 & n1332_1);
  assign n2277 = pstart_0_ & (pencrypt_0_ ? pkey_85_ : pkey_93_);
  assign n2278 = n2277 | (n_n2474 & ~n1327_1 & n1332_1);
  assign n2279 = pstart_0_ & (pencrypt_0_ ? pkey_94_ : pkey_102_);
  assign n2280 = n2279 | (pksi_130_ & n1327_1 & n1332_1);
  assign n2281 = pstart_0_ & (pencrypt_0_ ? pkey_22_ : pkey_30_);
  assign n2282 = n2281 | (n_n2517 & ~n1327_1 & n1332_1);
  assign n2283 = pstart_0_ & (pencrypt_0_ ? pkey_136_ : pkey_144_);
  assign n2284 = n2283 | (pksi_67_ & n1327_1 & n1332_1);
  assign n2285 = pstart_0_ & (pencrypt_0_ ? pkey_66_ : pkey_74_);
  assign n2286 = n2285 | (n_n2333 & ~n1327_1 & n1332_1);
  assign n2287 = pstart_0_ & (pencrypt_0_ ? pkey_89_ : pkey_97_);
  assign n2288 = n2287 | (pksi_46_ & n1327_1 & n1332_1);
  assign n2289 = pstart_0_ & (pencrypt_0_ ? pkey_112_ : pkey_120_);
  assign n2290 = n2289 | (pksi_47_ & n1327_1 & n1332_1);
  assign n2291 = pstart_0_ & (pencrypt_0_ ? pkey_42_ : pkey_50_);
  assign n2292 = n2291 | (pksi_13_ & n1327_1 & n1332_1);
  assign n2293 = pstart_0_ & (pencrypt_0_ ? pkey_144_ : pkey_152_);
  assign n2294 = n2293 | (pksi_57_ & n1327_1 & n1332_1);
  assign n2295 = pstart_0_ & (pencrypt_0_ ? pkey_123_ : pkey_66_);
  assign n2296 = n2295 | (n_n2333 & n1327_1 & n1332_1);
  assign n2297 = pstart_0_ & (pencrypt_0_ ? pkey_97_ : pkey_105_);
  assign n2298 = n2297 | (pksi_38_ & n1327_1 & n1332_1);
  assign n2299 = pstart_0_ & (pencrypt_0_ ? pkey_104_ : pkey_112_);
  assign n2300 = n2299 | (pksi_30_ & n1327_1 & n1332_1);
  assign n2301 = pstart_0_ & (pencrypt_0_ ? pkey_50_ : pkey_58_);
  assign n2302 = n2301 | (n_n2374 & n1327_1 & n1332_1);
  assign n2303 = pstart_0_ & (pencrypt_0_ ? pkey_152_ : pkey_160_);
  assign n2304 = n2303 | (pksi_53_ & n1327_1 & n1332_1);
  assign n2305 = pstart_0_ & (pencrypt_0_ ? pkey_82_ : pkey_90_);
  assign n2306 = n2305 | (n_n2337 & n1327_1 & n1332_1);
  assign n2307 = pstart_0_ & (pencrypt_0_ ? pkey_73_ : pkey_81_);
  assign n2308 = n2307 | (pksi_32_ & n1327_1 & n1332_1);
  assign n2309 = pstart_0_ & (pencrypt_0_ ? pkey_96_ : pkey_104_);
  assign n2310 = n2309 | (pksi_39_ & n1327_1 & n1332_1);
  assign n2311 = pstart_0_ & (pencrypt_0_ ? pkey_58_ : pkey_1_);
  assign n2312 = n2311 | (n_n2374 & ~n1327_1 & n1332_1);
  assign n2313 = pstart_0_ & (pencrypt_0_ ? pkey_56_ : pkey_227_);
  assign n2314 = n2313 | (pksi_4_ & n1327_1 & n1332_1);
  assign n2315 = pstart_0_ & (pencrypt_0_ ? pkey_160_ : pkey_168_);
  assign n2316 = n2315 | (pksi_63_ & n1327_1 & n1332_1);
  assign n2317 = pstart_0_ & (pencrypt_0_ ? pkey_74_ : pkey_82_);
  assign n2318 = n2317 | (pksi_36_ & n1327_1 & n1332_1);
  assign n2319 = pstart_0_ & (pencrypt_0_ ? pkey_81_ : pkey_89_);
  assign n2320 = n2319 | (pksi_24_ & n1327_1 & n1332_1);
  assign n2321 = pstart_0_ & (pencrypt_0_ ? pkey_88_ : pkey_96_);
  assign n2322 = n2321 | (pksi_29_ & n1327_1 & n1332_1);
  assign n2323 = pstart_0_ & (pencrypt_0_ ? pkey_1_ : pkey_9_);
  assign n2324 = n2323 | (pksi_18_ & n1327_1 & n1332_1);
  assign n2325 = pstart_0_ & (pencrypt_0_ ? pkey_234_ : pkey_242_);
  assign n2326 = n2325 | (pksi_85_ & n1327_1 & n1332_1);
  assign n2327 = pstart_0_ & (pencrypt_0_ ? pkey_192_ : pkey_200_);
  assign n2328 = n2327 | (pksi_89_ & n1327_1 & n1332_1);
  assign n2329 = pstart_0_ & (pencrypt_0_ ? pkey_187_ : pkey_130_);
  assign n2330 = n2329 | (n_n2301 & n1327_1 & n1332_1);
  assign n2331 = pstart_0_ & (pencrypt_0_ ? pkey_145_ : pkey_153_);
  assign n2332 = n2331 | (pksi_48_ & n1327_1 & n1332_1);
  assign n2333 = pstart_0_ & (pencrypt_0_ ? pkey_9_ : pkey_17_);
  assign n2334 = n2333 | (pksi_8_ & n1327_1 & n1332_1);
  assign n2335 = pstart_0_ & (pencrypt_0_ ? pkey_242_ : pkey_250_);
  assign n2336 = n2335 | (n_n2277 & n1327_1 & n1332_1);
  assign n2337 = pstart_0_ & (pencrypt_0_ ? pkey_249_ : pkey_192_);
  assign n2338 = n2337 | (n_n2288 & n1327_1 & n1332_1);
  assign n2339 = pstart_0_ & (pencrypt_0_ ? pkey_130_ : pkey_138_);
  assign n2340 = n2339 | (pksi_51_ & n1327_1 & n1332_1);
  assign n2341 = pstart_0_ & (pencrypt_0_ ? pkey_137_ : pkey_145_);
  assign n2342 = n2341 | (pksi_56_ & n1327_1 & n1332_1);
  assign n2343 = pstart_0_ & (pencrypt_0_ ? pkey_17_ : pkey_25_);
  assign n2344 = n2343 | (pksi_0_ & n1327_1 & n1332_1);
  assign n2345 = pstart_0_ & (pencrypt_0_ ? pkey_250_ : pkey_193_);
  assign n2346 = n2345 | (n_n2277 & ~n1327_1 & n1332_1);
  assign n2347 = pstart_0_ & (pencrypt_0_ ? pkey_208_ : pkey_216_);
  assign n2348 = n2347 | (pksi_81_ & n1327_1 & n1332_1);
  assign n2349 = pstart_0_ & (pencrypt_0_ ? pkey_171_ : pkey_179_);
  assign n2350 = n2349 | (pksi_68_ & n1327_1 & n1332_1);
  assign n2351 = pstart_0_ & (pencrypt_0_ ? pkey_129_ : pkey_137_);
  assign n2352 = n2351 | (pksi_66_ & n1327_1 & n1332_1);
  assign n2353 = pstart_0_ & (pencrypt_0_ ? pkey_193_ : pkey_201_);
  assign n2354 = n2353 | (n_n2280 & n1327_1 & n1332_1);
  assign n2355 = pstart_0_ & (pencrypt_0_ ? pkey_200_ : pkey_208_);
  assign n2356 = n2355 | (pksi_91_ & n1327_1 & n1332_1);
  assign n2357 = pstart_0_ & (pencrypt_0_ ? pkey_179_ : pkey_187_);
  assign n2358 = n2357 | (pksi_64_ & n1327_1 & n1332_1);
  assign n2359 = pstart_0_ & (pencrypt_0_ ? pkey_186_ : pkey_129_);
  assign n2360 = n2359 | (pksi_49_ & n1327_1 & n1332_1);
  assign n2361 = pstart_0_ & (pencrypt_0_ ? pkey_201_ : pkey_209_);
  assign n2362 = n2361 | (pksi_80_ & n1327_1 & n1332_1);
  assign n2363 = pstart_0_ & (pencrypt_0_ ? pkey_224_ : pkey_232_);
  assign n2364 = n2363 | (pksi_87_ & n1327_1 & n1332_1);
  assign n2365 = pstart_0_ & (pencrypt_0_ ? pkey_154_ : pkey_162_);
  assign n2366 = n2365 | (pksi_58_ & n1327_1 & n1332_1);
  assign n2367 = pstart_0_ & (pencrypt_0_ ? pkey_177_ : pkey_185_);
  assign n2368 = n2367 | (pksi_59_ & n1327_1 & n1332_1);
  assign n2369 = pstart_0_ & (pencrypt_0_ ? pkey_107_ : pkey_115_);
  assign n2370 = n2369 | (pksi_44_ & n1327_1 & n1332_1);
  assign n2371 = pstart_0_ & (pencrypt_0_ ? pkey_65_ : pkey_73_);
  assign n2372 = n2371 | (pksi_42_ & n1327_1 & n1332_1);
  assign n2373 = pstart_0_ & (pencrypt_0_ ? pkey_209_ : pkey_217_);
  assign n2374 = n2373 | (pksi_72_ & n1327_1 & n1332_1);
  assign n2375 = pstart_0_ & (pencrypt_0_ ? pkey_216_ : pkey_224_);
  assign n2376 = n2375 | (pksi_77_ & n1327_1 & n1332_1);
  assign n2377 = pstart_0_ & (pencrypt_0_ ? pkey_162_ : pkey_170_);
  assign n2378 = n2377 | (pksi_69_ & n1327_1 & n1332_1);
  assign n2379 = pstart_0_ & (pencrypt_0_ ? pkey_169_ : pkey_177_);
  assign n2380 = n2379 | (pksi_50_ & n1327_1 & n1332_1);
  assign n2381 = pstart_0_ & (pencrypt_0_ ? pkey_115_ : pkey_123_);
  assign n2382 = n2381 | (pksi_40_ & n1327_1 & n1332_1);
  assign n2383 = pstart_0_ & (pencrypt_0_ ? pkey_122_ : pkey_65_);
  assign n2384 = n2383 | (n_n2342 & ~n1327_1 & n1332_1);
  assign n2385 = pstart_0_ & (pencrypt_0_ ? pkey_217_ : pkey_225_);
  assign n2386 = n2385 | (pksi_94_ & n1327_1 & n1332_1);
  assign n2387 = pstart_0_ & (pencrypt_0_ ? pkey_240_ : pkey_248_);
  assign n2388 = n2387 | (pksi_95_ & n1327_1 & n1332_1);
  assign n2389 = pstart_0_ & (pencrypt_0_ ? pkey_138_ : pkey_146_);
  assign n2390 = n2389 | (pksi_60_ & n1327_1 & n1332_1);
  assign n2391 = pstart_0_ & (pencrypt_0_ ? pkey_161_ : pkey_169_);
  assign n2392 = n2391 | (pksi_62_ & n1327_1 & n1332_1);
  assign n2393 = pstart_0_ & (pencrypt_0_ ? pkey_72_ : pkey_80_);
  assign n2394 = n2393 | (pksi_43_ & n1327_1 & n1332_1);
  assign n2395 = pstart_0_ & (pencrypt_0_ ? pkey_2_ : pkey_10_);
  assign n2396 = n2395 | (n_n2365 & ~n1327_1 & n1332_1);
  assign n2397 = pstart_0_ & (pencrypt_0_ ? pkey_225_ : pkey_233_);
  assign n2398 = n2397 | (pksi_86_ & n1327_1 & n1332_1);
  assign n2399 = pstart_0_ & (pencrypt_0_ ? pkey_232_ : pkey_240_);
  assign n2400 = n2399 | (pksi_78_ & n1327_1 & n1332_1);
  assign n2401 = pstart_0_ & (pencrypt_0_ ? pkey_146_ : pkey_154_);
  assign n2402 = n2401 | (n_n2305 & n1327_1 & n1332_1);
  assign n2403 = pstart_0_ & (pencrypt_0_ ? pkey_153_ : pkey_161_);
  assign n2404 = n2403 | (pksi_70_ & n1327_1 & n1332_1);
  assign n2405 = pstart_0_ & (pencrypt_0_ ? pkey_80_ : pkey_88_);
  assign n2406 = n2405 | (pksi_33_ & n1327_1 & n1332_1);
  assign n2407 = pstart_0_ & (pencrypt_0_ ? pkey_59_ : pkey_2_);
  assign n2408 = n2407 | (n_n2365 & n1327_1 & n1332_1);
  assign n2409 = pstart_0_ & (pencrypt_0_ ? pkey_233_ : pkey_241_);
  assign n2410 = n2409 | (pksi_74_ & n1327_1 & n1332_1);
  assign n2411 = pstart_0_ & (pencrypt_0_ ? pkey_163_ : pkey_171_);
  assign n2412 = n2411 | (pksi_55_ & n1327_1 & n1332_1);
  assign n2413 = pstart_0_ & (pencrypt_0_ ? pkey_168_ : pkey_176_);
  assign n2414 = n2413 | (pksi_54_ & n1327_1 & n1332_1);
  assign n2415 = pstart_0_ & (pencrypt_0_ ? pkey_98_ : pkey_106_);
  assign n2416 = n2415 | (pksi_45_ & n1327_1 & n1332_1);
  assign n2417 = pstart_0_ & (pencrypt_0_ ? pkey_121_ : pkey_64_);
  assign n2418 = n2417 | (n_n2352 & n1327_1 & n1332_1);
  assign n2419 = pstart_0_ & (pencrypt_0_ ? pkey_51_ : pkey_59_);
  assign n2420 = n2419 | (pksi_16_ & n1327_1 & n1332_1);
  assign n2421 = pstart_0_ & (pencrypt_0_ ? pkey_10_ : pkey_18_);
  assign n2422 = n2421 | (pksi_12_ & n1327_1 & n1332_1);
  assign n2423 = pstart_0_ & (pencrypt_0_ ? pkey_241_ : pkey_249_);
  assign n2424 = n2423 | (pksi_83_ & n1327_1 & n1332_1);
  assign n2425 = pstart_0_ & (pencrypt_0_ ? pkey_248_ : pkey_163_);
  assign n2426 = n2425 | (pksi_76_ & n1327_1 & n1332_1);
  assign n2427 = pstart_0_ & (pencrypt_0_ ? pkey_176_ : pkey_184_);
  assign n2428 = n2427 | (pksi_71_ & n1327_1 & n1332_1);
  assign n2429 = pstart_0_ & (pencrypt_0_ ? pkey_90_ : pkey_98_);
  assign n2430 = n2429 | (n_n2337 & ~n1327_1 & n1332_1);
  assign n2431 = pstart_0_ & (pencrypt_0_ ? pkey_64_ : pkey_72_);
  assign n2432 = n2431 | (n_n2352 & ~n1327_1 & n1332_1);
  assign n2433 = pstart_0_ & (pencrypt_0_ ? pkey_43_ : pkey_51_);
  assign n2434 = n2433 | (pksi_20_ & n1327_1 & n1332_1);
  assign n2435 = pstart_0_ & (pencrypt_0_ ? pkey_18_ : pkey_26_);
  assign n2436 = n2435 | (n_n2369 & n1327_1 & n1332_1);
  assign n2437 = pstart_0_ & (pencrypt_0_ ? pkey_170_ : pkey_178_);
  assign n2438 = n2437 | (pksi_61_ & n1327_1 & n1332_1);
  assign n2439 = pstart_0_ & (pencrypt_0_ ? pkey_128_ : pkey_136_);
  assign n2440 = n2439 | (n_n2320 & ~n1327_1 & n1332_1);
  assign n2441 = pstart_0_ & (pencrypt_0_ ? pkey_184_ : pkey_99_);
  assign n2442 = n2441 | (pksi_52_ & n1327_1 & n1332_1);
  assign n2443 = pstart_0_ & (pencrypt_0_ ? pkey_114_ : pkey_122_);
  assign n2444 = n2443 | (n_n2342 & n1327_1 & n1332_1);
  assign n2445 = pstart_0_ & (pencrypt_0_ ? pkey_105_ : pkey_113_);
  assign n2446 = n2445 | (pksi_26_ & n1327_1 & n1332_1);
  assign n2447 = pstart_0_ & (pencrypt_0_ ? pkey_35_ : pkey_43_);
  assign n2448 = n2447 | (pksi_7_ & n1327_1 & n1332_1);
  assign n2449 = pstart_0_ & (pencrypt_0_ ? pkey_26_ : pkey_34_);
  assign n2450 = n2449 | (n_n2369 & ~n1327_1 & n1332_1);
  assign n2451 = pstart_0_ & (pencrypt_0_ ? pkey_178_ : pkey_186_);
  assign n2452 = n2451 | (n_n2310 & n1327_1 & n1332_1);
  assign n2453 = pstart_0_ & (pencrypt_0_ ? pkey_185_ : pkey_128_);
  assign n2454 = n2453 | (n_n2320 & n1327_1 & n1332_1);
  assign n2455 = pstart_0_ & (pencrypt_0_ ? pkey_99_ : pkey_107_);
  assign n2456 = n2455 | (pksi_31_ & n1327_1 & n1332_1);
  assign n2457 = pstart_0_ & (pencrypt_0_ ? pkey_106_ : pkey_114_);
  assign n2458 = n2457 | (pksi_37_ & n1327_1 & n1332_1);
  assign n2459 = pstart_0_ & (pencrypt_0_ ? pkey_113_ : pkey_121_);
  assign n2460 = n2459 | (pksi_35_ & n1327_1 & n1332_1);
  assign n2461 = pstart_0_ & (pencrypt_0_ ? pkey_120_ : pkey_35_);
  assign n2462 = n2461 | (pksi_28_ & n1327_1 & n1332_1);
  assign n2463 = pstart_0_ & (pencrypt_0_ ? pkey_34_ : pkey_42_);
  assign n2464 = n2463 | (pksi_21_ & n1327_1 & n1332_1);
  assign n2465 = ~pencrypt_0_ & ~pstart_0_ & ~pcount_1_ & ~pcount_0_;
  assign n2466 = pcount_2_ ? ~pencrypt_0_ : (~pstart_0_ & pencrypt_0_);
  assign n2467 = n1341 | ~n1330 | (~pcount_2_ & n1329);
  always @ (posedge clk) begin
    pksi_17_ <= n853;
    pksi_185_ <= n857;
    n_n2410 <= n861;
    pksi_170_ <= n866;
    pksi_155_ <= n870;
    pksi_147_ <= n874;
    pksi_109_ <= n878;
    n_n2513 <= n882;
    pksi_19_ <= n887;
    n_n2396 <= n891;
    n_n2412 <= n896;
    n_n121 <= n901;
    pksi_148_ <= n906;
    n_n2448 <= n910;
    pksi_107_ <= n915;
    pksi_110_ <= n919;
    pksi_9_ <= n923;
    pksi_176_ <= n927;
    pksi_180_ <= n931;
    pksi_178_ <= n935;
    pksi_135_ <= n939;
    pksi_129_ <= n943;
    pksi_100_ <= n947;
    pksi_117_ <= n951;
    pksi_118_ <= n955;
    pksi_5_ <= n959;
    pksi_169_ <= n963;
    n_n2408 <= n967;
    pksi_184_ <= n972;
    pksi_125_ <= n976;
    pksi_138_ <= n980;
    pksi_114_ <= n984;
    pksi_99_ <= n988;
    pksi_85_ <= n992;
    pksi_14_ <= n996;
    pksi_4_ <= n1000;
    pksi_186_ <= n1004;
    n_n2420 <= n1008;
    pksi_141_ <= n1013;
    pksi_113_ <= n1017;
    pksi_115_ <= n1021;
    pksi_98_ <= n1025;
    pksi_2_ <= n1029;
    pksi_23_ <= n1033;
    pksi_177_ <= n1037;
    pksi_189_ <= n1041;
    n_n2485 <= n1045;
    n_n2495 <= n1050;
    pksi_97_ <= n1055;
    pksi_102_ <= n1059;
    pksi_11_ <= n1063;
    pksi_173_ <= n1067;
    pksi_179_ <= n1071;
    pksi_171_ <= n1075;
    pksi_104_ <= n1079;
    pksi_103_ <= n1083;
    n_n2384 <= n1087;
    pksi_183_ <= n1092;
    pksi_172_ <= n1096;
    n_n2416 <= n1100;
    pksi_116_ <= n1105;
    pksi_96_ <= n1109;
    pksi_119_ <= n1113;
    pksi_84_ <= n1117;
    pksi_159_ <= n1121;
    n_n2440 <= n1125;
    pksi_160_ <= n1130;
    pksi_128_ <= n1134;
    pksi_127_ <= n1138;
    pksi_142_ <= n1142;
    n_n2272 <= n1146;
    pksi_149_ <= n1151;
    pksi_162_ <= n1155;
    pksi_154_ <= n1159;
    pksi_121_ <= n1163;
    pksi_134_ <= n1167;
    pksi_126_ <= n1171;
    pksi_82_ <= n1175;
    n_n2430 <= n1179;
    pksi_153_ <= n1184;
    pksi_165_ <= n1188;
    pksi_137_ <= n1192;
    n_n2481 <= n1196;
    pksi_101_ <= n1201;
    pksi_93_ <= n1205;
    pksi_161_ <= n1209;
    pksi_156_ <= n1213;
    n_n2452 <= n1217;
    n_n2462 <= n1222;
    pksi_123_ <= n1227;
    pksi_111_ <= n1231;
    pksi_92_ <= n1235;
    pksi_15_ <= n1239;
    n_n109 <= n1243;
    pksi_145_ <= n1248;
    pksi_144_ <= n1252;
    pksi_150_ <= n1256;
    pksi_124_ <= n1260;
    pksi_132_ <= n1264;
    pksi_130_ <= n1268;
    pksi_105_ <= n1272;
    pksi_112_ <= n1276;
    n_n10 <= n1280;
    pksi_6_ <= n1285;
    pksi_188_ <= n1289;
    pksi_152_ <= n1293;
    pksi_163_ <= n1297;
    pksi_166_ <= n1301;
    pksi_131_ <= n1305;
    n_n2474 <= n1309;
    pksi_136_ <= n1314;
    pksi_108_ <= n1318;
    n_n2517 <= n1322;
    n_n2268 <= n1327;
    pksi_175_ <= n1332;
    pksi_190_ <= n1336;
    pksi_164_ <= n1340;
    pksi_158_ <= n1344;
    pksi_167_ <= n1348;
    pksi_133_ <= n1352;
    n_n2476 <= n1356;
    pksi_122_ <= n1361;
    n_n2507 <= n1365;
    pksi_75_ <= n1370;
    pksi_182_ <= n1374;
    pksi_174_ <= n1378;
    pksi_157_ <= n1382;
    pksi_151_ <= n1386;
    pksi_146_ <= n1390;
    pksi_140_ <= n1394;
    pksi_120_ <= n1398;
    n_n168 <= n1402;
    pksi_106_ <= n1407;
    pksi_57_ <= n1411;
    pksi_36_ <= n1415;
    pksi_38_ <= n1419;
    pksi_28_ <= n1423;
    n_n2374 <= n1427;
    pksi_53_ <= n1432;
    pksi_27_ <= n1436;
    pksi_26_ <= n1440;
    pksi_47_ <= n1444;
    pksi_1_ <= n1448;
    pksi_63_ <= n1452;
    pksi_34_ <= n1456;
    pksi_24_ <= n1460;
    pksi_30_ <= n1464;
    pksi_18_ <= n1468;
    pksi_79_ <= n1472;
    pksi_54_ <= n1476;
    n_n2337 <= n1480;
    pksi_46_ <= n1485;
    pksi_39_ <= n1489;
    pksi_8_ <= n1493;
    n_n2277 <= n1497;
    pksi_91_ <= n1502;
    pksi_51_ <= n1506;
    pksi_70_ <= n1510;
    pksi_0_ <= n1514;
    pksi_73_ <= n1518;
    pksi_89_ <= n1522;
    pksi_60_ <= n1526;
    pksi_48_ <= n1530;
    pksi_22_ <= n1534;
    n_n2280 <= n1538;
    pksi_77_ <= n1543;
    pksi_64_ <= n1547;
    pksi_56_ <= n1551;
    pksi_80_ <= n1555;
    pksi_81_ <= n1559;
    n_n2301 <= n1563;
    pksi_66_ <= n1568;
    pksi_72_ <= n1572;
    pksi_78_ <= n1576;
    pksi_69_ <= n1580;
    n_n2320 <= n1584;
    pksi_40_ <= n1589;
    pksi_32_ <= n1593;
    pksi_94_ <= n1597;
    pksi_87_ <= n1601;
    pksi_61_ <= n1605;
    pksi_59_ <= n1609;
    n_n2333 <= n1613;
    pksi_42_ <= n1618;
    pksi_86_ <= n1622;
    pksi_76_ <= n1626;
    n_n2305 <= n1630;
    pksi_50_ <= n1635;
    pksi_33_ <= n1639;
    pksi_12_ <= n1643;
    pksi_74_ <= n1647;
    pksi_95_ <= n1651;
    pksi_58_ <= n1655;
    pksi_62_ <= n1659;
    pksi_29_ <= n1663;
    pksi_3_ <= n1667;
    pksi_83_ <= n1671;
    pksi_68_ <= n1675;
    pksi_71_ <= n1679;
    pksi_37_ <= n1683;
    pksi_41_ <= n1687;
    n_n2365 <= n1691;
    n_n2369 <= n1696;
    n_n2288 <= n1701;
    pksi_55_ <= n1706;
    pksi_52_ <= n1710;
    pksi_45_ <= n1714;
    pksi_43_ <= n1718;
    pksi_16_ <= n1722;
    pksi_10_ <= n1726;
    n_n2310 <= n1730;
    pksi_67_ <= n1735;
    pksi_31_ <= n1739;
    pksi_25_ <= n1743;
    pksi_35_ <= n1747;
    pksi_20_ <= n1751;
    pksi_21_ <= n1755;
    pksi_49_ <= n1759;
    pksi_65_ <= n1763;
    pksi_44_ <= n1767;
    n_n2342 <= n1771;
    n_n2352 <= n1776;
    pksi_7_ <= n1781;
    pksi_13_ <= n1785;
  end
endmodule


