// Benchmark "TOP" written by ABC on Tue Mar  5 09:56:12 2019

module des ( 
    Preset_0_, Poutreg_63_, Poutreg_62_, Poutreg_61_, Poutreg_60_,
    Poutreg_59_, Poutreg_58_, Poutreg_57_, Poutreg_56_, Poutreg_55_,
    Poutreg_54_, Poutreg_53_, Poutreg_52_, Poutreg_51_, Poutreg_50_,
    Poutreg_49_, Poutreg_48_, Poutreg_47_, Poutreg_46_, Poutreg_45_,
    Poutreg_44_, Poutreg_43_, Poutreg_42_, Poutreg_41_, Poutreg_40_,
    Poutreg_39_, Poutreg_38_, Poutreg_37_, Poutreg_36_, Poutreg_35_,
    Poutreg_34_, Poutreg_33_, Poutreg_32_, Poutreg_31_, Poutreg_30_,
    Poutreg_29_, Poutreg_28_, Poutreg_27_, Poutreg_26_, Poutreg_25_,
    Poutreg_24_, Poutreg_23_, Poutreg_22_, Poutreg_21_, Poutreg_20_,
    Poutreg_19_, Poutreg_18_, Poutreg_17_, Poutreg_16_, Poutreg_15_,
    Poutreg_14_, Poutreg_13_, Poutreg_12_, Poutreg_11_, Poutreg_10_,
    Poutreg_9_, Poutreg_8_, Poutreg_7_, Poutreg_6_, Poutreg_5_, Poutreg_4_,
    Poutreg_3_, Poutreg_2_, Poutreg_1_, Poutreg_0_, Pload_key_0_,
    Pinreg_55_, Pinreg_54_, Pinreg_53_, Pinreg_52_, Pinreg_51_, Pinreg_50_,
    Pinreg_49_, Pinreg_48_, Pinreg_47_, Pinreg_46_, Pinreg_45_, Pinreg_44_,
    Pinreg_43_, Pinreg_42_, Pinreg_41_, Pinreg_40_, Pinreg_39_, Pinreg_38_,
    Pinreg_37_, Pinreg_36_, Pinreg_35_, Pinreg_34_, Pinreg_33_, Pinreg_32_,
    Pinreg_31_, Pinreg_30_, Pinreg_29_, Pinreg_28_, Pinreg_27_, Pinreg_26_,
    Pinreg_25_, Pinreg_24_, Pinreg_23_, Pinreg_22_, Pinreg_21_, Pinreg_20_,
    Pinreg_19_, Pinreg_18_, Pinreg_17_, Pinreg_16_, Pinreg_15_, Pinreg_14_,
    Pinreg_13_, Pinreg_12_, Pinreg_11_, Pinreg_10_, Pinreg_9_, Pinreg_8_,
    Pinreg_7_, Pinreg_6_, Pinreg_5_, Pinreg_4_, Pinreg_3_, Pinreg_2_,
    Pinreg_1_, Pinreg_0_, Pencrypt_mode_0_, Pencrypt_0_, Pdata_in_7_,
    Pdata_in_6_, Pdata_in_5_, Pdata_in_4_, Pdata_in_3_, Pdata_in_2_,
    Pdata_in_1_, Pdata_in_0_, Pdata_63_, Pdata_62_, Pdata_61_, Pdata_60_,
    Pdata_59_, Pdata_58_, Pdata_57_, Pdata_56_, Pdata_55_, Pdata_54_,
    Pdata_53_, Pdata_52_, Pdata_51_, Pdata_50_, Pdata_49_, Pdata_48_,
    Pdata_47_, Pdata_46_, Pdata_45_, Pdata_44_, Pdata_43_, Pdata_42_,
    Pdata_41_, Pdata_40_, Pdata_39_, Pdata_38_, Pdata_37_, Pdata_36_,
    Pdata_35_, Pdata_34_, Pdata_33_, Pdata_32_, Pdata_31_, Pdata_30_,
    Pdata_29_, Pdata_28_, Pdata_27_, Pdata_26_, Pdata_25_, Pdata_24_,
    Pdata_23_, Pdata_22_, Pdata_21_, Pdata_20_, Pdata_19_, Pdata_18_,
    Pdata_17_, Pdata_16_, Pdata_15_, Pdata_14_, Pdata_13_, Pdata_12_,
    Pdata_11_, Pdata_10_, Pdata_9_, Pdata_8_, Pdata_7_, Pdata_6_, Pdata_5_,
    Pdata_4_, Pdata_3_, Pdata_2_, Pdata_1_, Pdata_0_, Pcount_3_, Pcount_2_,
    Pcount_1_, Pcount_0_, PD_27_, PD_26_, PD_25_, PD_24_, PD_23_, PD_22_,
    PD_21_, PD_20_, PD_19_, PD_18_, PD_17_, PD_16_, PD_15_, PD_14_, PD_13_,
    PD_12_, PD_11_, PD_10_, PD_9_, PD_8_, PD_7_, PD_6_, PD_5_, PD_4_,
    PD_3_, PD_2_, PD_1_, PD_0_, PC_27_, PC_26_, PC_25_, PC_24_, PC_23_,
    PC_22_, PC_21_, PC_20_, PC_19_, PC_18_, PC_17_, PC_16_, PC_15_, PC_14_,
    PC_13_, PC_12_, PC_11_, PC_10_, PC_9_, PC_8_, PC_7_, PC_6_, PC_5_,
    PC_4_, PC_3_, PC_2_, PC_1_, PC_0_,
    Poutreg_new_63_, Poutreg_new_62_, Poutreg_new_61_, Poutreg_new_60_,
    Poutreg_new_59_, Poutreg_new_58_, Poutreg_new_57_, Poutreg_new_56_,
    Poutreg_new_55_, Poutreg_new_54_, Poutreg_new_53_, Poutreg_new_52_,
    Poutreg_new_51_, Poutreg_new_50_, Poutreg_new_49_, Poutreg_new_48_,
    Poutreg_new_47_, Poutreg_new_46_, Poutreg_new_45_, Poutreg_new_44_,
    Poutreg_new_43_, Poutreg_new_42_, Poutreg_new_41_, Poutreg_new_40_,
    Poutreg_new_39_, Poutreg_new_38_, Poutreg_new_37_, Poutreg_new_36_,
    Poutreg_new_35_, Poutreg_new_34_, Poutreg_new_33_, Poutreg_new_32_,
    Poutreg_new_31_, Poutreg_new_30_, Poutreg_new_29_, Poutreg_new_28_,
    Poutreg_new_27_, Poutreg_new_26_, Poutreg_new_25_, Poutreg_new_24_,
    Poutreg_new_23_, Poutreg_new_22_, Poutreg_new_21_, Poutreg_new_20_,
    Poutreg_new_19_, Poutreg_new_18_, Poutreg_new_17_, Poutreg_new_16_,
    Poutreg_new_15_, Poutreg_new_14_, Poutreg_new_13_, Poutreg_new_12_,
    Poutreg_new_11_, Poutreg_new_10_, Poutreg_new_9_, Poutreg_new_8_,
    Poutreg_new_7_, Poutreg_new_6_, Poutreg_new_5_, Poutreg_new_4_,
    Poutreg_new_3_, Poutreg_new_2_, Poutreg_new_1_, Poutreg_new_0_,
    Pinreg_new_55_, Pinreg_new_54_, Pinreg_new_53_, Pinreg_new_52_,
    Pinreg_new_51_, Pinreg_new_50_, Pinreg_new_49_, Pinreg_new_48_,
    Pinreg_new_47_, Pinreg_new_46_, Pinreg_new_45_, Pinreg_new_44_,
    Pinreg_new_43_, Pinreg_new_42_, Pinreg_new_41_, Pinreg_new_40_,
    Pinreg_new_39_, Pinreg_new_38_, Pinreg_new_37_, Pinreg_new_36_,
    Pinreg_new_35_, Pinreg_new_34_, Pinreg_new_33_, Pinreg_new_32_,
    Pinreg_new_31_, Pinreg_new_30_, Pinreg_new_29_, Pinreg_new_28_,
    Pinreg_new_27_, Pinreg_new_26_, Pinreg_new_25_, Pinreg_new_24_,
    Pinreg_new_23_, Pinreg_new_22_, Pinreg_new_21_, Pinreg_new_20_,
    Pinreg_new_19_, Pinreg_new_18_, Pinreg_new_17_, Pinreg_new_16_,
    Pinreg_new_15_, Pinreg_new_14_, Pinreg_new_13_, Pinreg_new_12_,
    Pinreg_new_11_, Pinreg_new_10_, Pinreg_new_9_, Pinreg_new_8_,
    Pinreg_new_7_, Pinreg_new_6_, Pinreg_new_5_, Pinreg_new_4_,
    Pinreg_new_3_, Pinreg_new_2_, Pinreg_new_1_, Pinreg_new_0_,
    Pencrypt_mode_new_0_, Pdata_new_63_, Pdata_new_62_, Pdata_new_61_,
    Pdata_new_60_, Pdata_new_59_, Pdata_new_58_, Pdata_new_57_,
    Pdata_new_56_, Pdata_new_55_, Pdata_new_54_, Pdata_new_53_,
    Pdata_new_52_, Pdata_new_51_, Pdata_new_50_, Pdata_new_49_,
    Pdata_new_48_, Pdata_new_47_, Pdata_new_46_, Pdata_new_45_,
    Pdata_new_44_, Pdata_new_43_, Pdata_new_42_, Pdata_new_41_,
    Pdata_new_40_, Pdata_new_39_, Pdata_new_38_, Pdata_new_37_,
    Pdata_new_36_, Pdata_new_35_, Pdata_new_34_, Pdata_new_33_,
    Pdata_new_32_, Pdata_new_31_, Pdata_new_30_, Pdata_new_29_,
    Pdata_new_28_, Pdata_new_27_, Pdata_new_26_, Pdata_new_25_,
    Pdata_new_24_, Pdata_new_23_, Pdata_new_22_, Pdata_new_21_,
    Pdata_new_20_, Pdata_new_19_, Pdata_new_18_, Pdata_new_17_,
    Pdata_new_16_, Pdata_new_15_, Pdata_new_14_, Pdata_new_13_,
    Pdata_new_12_, Pdata_new_11_, Pdata_new_10_, Pdata_new_9_,
    Pdata_new_8_, Pdata_new_7_, Pdata_new_6_, Pdata_new_5_, Pdata_new_4_,
    Pdata_new_3_, Pdata_new_2_, Pdata_new_1_, Pdata_new_0_, Pcount_new_3_,
    Pcount_new_2_, Pcount_new_1_, Pcount_new_0_, PD_new_27_, PD_new_26_,
    PD_new_25_, PD_new_24_, PD_new_23_, PD_new_22_, PD_new_21_, PD_new_20_,
    PD_new_19_, PD_new_18_, PD_new_17_, PD_new_16_, PD_new_15_, PD_new_14_,
    PD_new_13_, PD_new_12_, PD_new_11_, PD_new_10_, PD_new_9_, PD_new_8_,
    PD_new_7_, PD_new_6_, PD_new_5_, PD_new_4_, PD_new_3_, PD_new_2_,
    PD_new_1_, PD_new_0_, PC_new_27_, PC_new_26_, PC_new_25_, PC_new_24_,
    PC_new_23_, PC_new_22_, PC_new_21_, PC_new_20_, PC_new_19_, PC_new_18_,
    PC_new_17_, PC_new_16_, PC_new_15_, PC_new_14_, PC_new_13_, PC_new_12_,
    PC_new_11_, PC_new_10_, PC_new_9_, PC_new_8_, PC_new_7_, PC_new_6_,
    PC_new_5_, PC_new_4_, PC_new_3_, PC_new_2_, PC_new_1_, PC_new_0_  );
  input  Preset_0_, Poutreg_63_, Poutreg_62_, Poutreg_61_, Poutreg_60_,
    Poutreg_59_, Poutreg_58_, Poutreg_57_, Poutreg_56_, Poutreg_55_,
    Poutreg_54_, Poutreg_53_, Poutreg_52_, Poutreg_51_, Poutreg_50_,
    Poutreg_49_, Poutreg_48_, Poutreg_47_, Poutreg_46_, Poutreg_45_,
    Poutreg_44_, Poutreg_43_, Poutreg_42_, Poutreg_41_, Poutreg_40_,
    Poutreg_39_, Poutreg_38_, Poutreg_37_, Poutreg_36_, Poutreg_35_,
    Poutreg_34_, Poutreg_33_, Poutreg_32_, Poutreg_31_, Poutreg_30_,
    Poutreg_29_, Poutreg_28_, Poutreg_27_, Poutreg_26_, Poutreg_25_,
    Poutreg_24_, Poutreg_23_, Poutreg_22_, Poutreg_21_, Poutreg_20_,
    Poutreg_19_, Poutreg_18_, Poutreg_17_, Poutreg_16_, Poutreg_15_,
    Poutreg_14_, Poutreg_13_, Poutreg_12_, Poutreg_11_, Poutreg_10_,
    Poutreg_9_, Poutreg_8_, Poutreg_7_, Poutreg_6_, Poutreg_5_, Poutreg_4_,
    Poutreg_3_, Poutreg_2_, Poutreg_1_, Poutreg_0_, Pload_key_0_,
    Pinreg_55_, Pinreg_54_, Pinreg_53_, Pinreg_52_, Pinreg_51_, Pinreg_50_,
    Pinreg_49_, Pinreg_48_, Pinreg_47_, Pinreg_46_, Pinreg_45_, Pinreg_44_,
    Pinreg_43_, Pinreg_42_, Pinreg_41_, Pinreg_40_, Pinreg_39_, Pinreg_38_,
    Pinreg_37_, Pinreg_36_, Pinreg_35_, Pinreg_34_, Pinreg_33_, Pinreg_32_,
    Pinreg_31_, Pinreg_30_, Pinreg_29_, Pinreg_28_, Pinreg_27_, Pinreg_26_,
    Pinreg_25_, Pinreg_24_, Pinreg_23_, Pinreg_22_, Pinreg_21_, Pinreg_20_,
    Pinreg_19_, Pinreg_18_, Pinreg_17_, Pinreg_16_, Pinreg_15_, Pinreg_14_,
    Pinreg_13_, Pinreg_12_, Pinreg_11_, Pinreg_10_, Pinreg_9_, Pinreg_8_,
    Pinreg_7_, Pinreg_6_, Pinreg_5_, Pinreg_4_, Pinreg_3_, Pinreg_2_,
    Pinreg_1_, Pinreg_0_, Pencrypt_mode_0_, Pencrypt_0_, Pdata_in_7_,
    Pdata_in_6_, Pdata_in_5_, Pdata_in_4_, Pdata_in_3_, Pdata_in_2_,
    Pdata_in_1_, Pdata_in_0_, Pdata_63_, Pdata_62_, Pdata_61_, Pdata_60_,
    Pdata_59_, Pdata_58_, Pdata_57_, Pdata_56_, Pdata_55_, Pdata_54_,
    Pdata_53_, Pdata_52_, Pdata_51_, Pdata_50_, Pdata_49_, Pdata_48_,
    Pdata_47_, Pdata_46_, Pdata_45_, Pdata_44_, Pdata_43_, Pdata_42_,
    Pdata_41_, Pdata_40_, Pdata_39_, Pdata_38_, Pdata_37_, Pdata_36_,
    Pdata_35_, Pdata_34_, Pdata_33_, Pdata_32_, Pdata_31_, Pdata_30_,
    Pdata_29_, Pdata_28_, Pdata_27_, Pdata_26_, Pdata_25_, Pdata_24_,
    Pdata_23_, Pdata_22_, Pdata_21_, Pdata_20_, Pdata_19_, Pdata_18_,
    Pdata_17_, Pdata_16_, Pdata_15_, Pdata_14_, Pdata_13_, Pdata_12_,
    Pdata_11_, Pdata_10_, Pdata_9_, Pdata_8_, Pdata_7_, Pdata_6_, Pdata_5_,
    Pdata_4_, Pdata_3_, Pdata_2_, Pdata_1_, Pdata_0_, Pcount_3_, Pcount_2_,
    Pcount_1_, Pcount_0_, PD_27_, PD_26_, PD_25_, PD_24_, PD_23_, PD_22_,
    PD_21_, PD_20_, PD_19_, PD_18_, PD_17_, PD_16_, PD_15_, PD_14_, PD_13_,
    PD_12_, PD_11_, PD_10_, PD_9_, PD_8_, PD_7_, PD_6_, PD_5_, PD_4_,
    PD_3_, PD_2_, PD_1_, PD_0_, PC_27_, PC_26_, PC_25_, PC_24_, PC_23_,
    PC_22_, PC_21_, PC_20_, PC_19_, PC_18_, PC_17_, PC_16_, PC_15_, PC_14_,
    PC_13_, PC_12_, PC_11_, PC_10_, PC_9_, PC_8_, PC_7_, PC_6_, PC_5_,
    PC_4_, PC_3_, PC_2_, PC_1_, PC_0_;
  output Poutreg_new_63_, Poutreg_new_62_, Poutreg_new_61_, Poutreg_new_60_,
    Poutreg_new_59_, Poutreg_new_58_, Poutreg_new_57_, Poutreg_new_56_,
    Poutreg_new_55_, Poutreg_new_54_, Poutreg_new_53_, Poutreg_new_52_,
    Poutreg_new_51_, Poutreg_new_50_, Poutreg_new_49_, Poutreg_new_48_,
    Poutreg_new_47_, Poutreg_new_46_, Poutreg_new_45_, Poutreg_new_44_,
    Poutreg_new_43_, Poutreg_new_42_, Poutreg_new_41_, Poutreg_new_40_,
    Poutreg_new_39_, Poutreg_new_38_, Poutreg_new_37_, Poutreg_new_36_,
    Poutreg_new_35_, Poutreg_new_34_, Poutreg_new_33_, Poutreg_new_32_,
    Poutreg_new_31_, Poutreg_new_30_, Poutreg_new_29_, Poutreg_new_28_,
    Poutreg_new_27_, Poutreg_new_26_, Poutreg_new_25_, Poutreg_new_24_,
    Poutreg_new_23_, Poutreg_new_22_, Poutreg_new_21_, Poutreg_new_20_,
    Poutreg_new_19_, Poutreg_new_18_, Poutreg_new_17_, Poutreg_new_16_,
    Poutreg_new_15_, Poutreg_new_14_, Poutreg_new_13_, Poutreg_new_12_,
    Poutreg_new_11_, Poutreg_new_10_, Poutreg_new_9_, Poutreg_new_8_,
    Poutreg_new_7_, Poutreg_new_6_, Poutreg_new_5_, Poutreg_new_4_,
    Poutreg_new_3_, Poutreg_new_2_, Poutreg_new_1_, Poutreg_new_0_,
    Pinreg_new_55_, Pinreg_new_54_, Pinreg_new_53_, Pinreg_new_52_,
    Pinreg_new_51_, Pinreg_new_50_, Pinreg_new_49_, Pinreg_new_48_,
    Pinreg_new_47_, Pinreg_new_46_, Pinreg_new_45_, Pinreg_new_44_,
    Pinreg_new_43_, Pinreg_new_42_, Pinreg_new_41_, Pinreg_new_40_,
    Pinreg_new_39_, Pinreg_new_38_, Pinreg_new_37_, Pinreg_new_36_,
    Pinreg_new_35_, Pinreg_new_34_, Pinreg_new_33_, Pinreg_new_32_,
    Pinreg_new_31_, Pinreg_new_30_, Pinreg_new_29_, Pinreg_new_28_,
    Pinreg_new_27_, Pinreg_new_26_, Pinreg_new_25_, Pinreg_new_24_,
    Pinreg_new_23_, Pinreg_new_22_, Pinreg_new_21_, Pinreg_new_20_,
    Pinreg_new_19_, Pinreg_new_18_, Pinreg_new_17_, Pinreg_new_16_,
    Pinreg_new_15_, Pinreg_new_14_, Pinreg_new_13_, Pinreg_new_12_,
    Pinreg_new_11_, Pinreg_new_10_, Pinreg_new_9_, Pinreg_new_8_,
    Pinreg_new_7_, Pinreg_new_6_, Pinreg_new_5_, Pinreg_new_4_,
    Pinreg_new_3_, Pinreg_new_2_, Pinreg_new_1_, Pinreg_new_0_,
    Pencrypt_mode_new_0_, Pdata_new_63_, Pdata_new_62_, Pdata_new_61_,
    Pdata_new_60_, Pdata_new_59_, Pdata_new_58_, Pdata_new_57_,
    Pdata_new_56_, Pdata_new_55_, Pdata_new_54_, Pdata_new_53_,
    Pdata_new_52_, Pdata_new_51_, Pdata_new_50_, Pdata_new_49_,
    Pdata_new_48_, Pdata_new_47_, Pdata_new_46_, Pdata_new_45_,
    Pdata_new_44_, Pdata_new_43_, Pdata_new_42_, Pdata_new_41_,
    Pdata_new_40_, Pdata_new_39_, Pdata_new_38_, Pdata_new_37_,
    Pdata_new_36_, Pdata_new_35_, Pdata_new_34_, Pdata_new_33_,
    Pdata_new_32_, Pdata_new_31_, Pdata_new_30_, Pdata_new_29_,
    Pdata_new_28_, Pdata_new_27_, Pdata_new_26_, Pdata_new_25_,
    Pdata_new_24_, Pdata_new_23_, Pdata_new_22_, Pdata_new_21_,
    Pdata_new_20_, Pdata_new_19_, Pdata_new_18_, Pdata_new_17_,
    Pdata_new_16_, Pdata_new_15_, Pdata_new_14_, Pdata_new_13_,
    Pdata_new_12_, Pdata_new_11_, Pdata_new_10_, Pdata_new_9_,
    Pdata_new_8_, Pdata_new_7_, Pdata_new_6_, Pdata_new_5_, Pdata_new_4_,
    Pdata_new_3_, Pdata_new_2_, Pdata_new_1_, Pdata_new_0_, Pcount_new_3_,
    Pcount_new_2_, Pcount_new_1_, Pcount_new_0_, PD_new_27_, PD_new_26_,
    PD_new_25_, PD_new_24_, PD_new_23_, PD_new_22_, PD_new_21_, PD_new_20_,
    PD_new_19_, PD_new_18_, PD_new_17_, PD_new_16_, PD_new_15_, PD_new_14_,
    PD_new_13_, PD_new_12_, PD_new_11_, PD_new_10_, PD_new_9_, PD_new_8_,
    PD_new_7_, PD_new_6_, PD_new_5_, PD_new_4_, PD_new_3_, PD_new_2_,
    PD_new_1_, PD_new_0_, PC_new_27_, PC_new_26_, PC_new_25_, PC_new_24_,
    PC_new_23_, PC_new_22_, PC_new_21_, PC_new_20_, PC_new_19_, PC_new_18_,
    PC_new_17_, PC_new_16_, PC_new_15_, PC_new_14_, PC_new_13_, PC_new_12_,
    PC_new_11_, PC_new_10_, PC_new_9_, PC_new_8_, PC_new_7_, PC_new_6_,
    PC_new_5_, PC_new_4_, PC_new_3_, PC_new_2_, PC_new_1_, PC_new_0_;
  wire n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
    n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
    n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
    n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
    n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
    n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
    n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
    n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
    n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
    n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
    n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
    n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
    n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
    n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
    n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
    n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
    n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
    n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
    n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
    n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
    n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
    n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
    n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
    n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
    n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
    n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
    n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
    n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
    n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
    n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
    n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
    n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
    n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
    n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
    n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
    n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
    n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
    n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
    n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
    n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
    n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
    n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
    n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
    n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
    n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
    n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
    n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
    n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
    n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
    n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
    n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
    n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
    n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
    n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
    n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
    n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
    n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
    n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
    n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
    n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
    n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
    n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
    n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
    n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
    n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
    n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
    n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
    n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
    n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
    n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
    n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
    n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
    n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
    n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
    n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
    n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
    n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
    n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
    n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
    n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
    n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
    n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
    n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
    n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
    n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
    n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
    n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
    n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
    n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
    n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
    n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
    n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
    n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
    n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
    n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
    n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
    n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
    n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
    n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
    n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
    n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
    n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
    n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
    n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
    n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
    n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
    n1997, n1998;
  assign Poutreg_new_63_ = ~n747;
  assign Poutreg_new_62_ = ~n849;
  assign Poutreg_new_61_ = ~n748;
  assign Poutreg_new_60_ = ~n845;
  assign Poutreg_new_59_ = ~n749;
  assign Poutreg_new_58_ = ~n841;
  assign Poutreg_new_57_ = ~n750;
  assign Poutreg_new_56_ = ~n836;
  assign Poutreg_new_55_ = ~n751;
  assign Poutreg_new_54_ = ~n868;
  assign Poutreg_new_53_ = ~n752;
  assign Poutreg_new_52_ = ~n838;
  assign Poutreg_new_51_ = ~n753;
  assign Poutreg_new_50_ = ~n867;
  assign Poutreg_new_49_ = ~n754;
  assign Poutreg_new_48_ = ~n866;
  assign Poutreg_new_47_ = ~n755;
  assign Poutreg_new_46_ = ~n865;
  assign Poutreg_new_45_ = ~n756;
  assign Poutreg_new_44_ = ~n864;
  assign Poutreg_new_43_ = ~n757;
  assign Poutreg_new_42_ = ~n863;
  assign Poutreg_new_41_ = ~n758;
  assign Poutreg_new_40_ = ~n862;
  assign Poutreg_new_39_ = ~n759;
  assign Poutreg_new_38_ = ~n861;
  assign Poutreg_new_37_ = ~n760;
  assign Poutreg_new_36_ = ~n860;
  assign Poutreg_new_35_ = ~n761;
  assign Poutreg_new_34_ = ~n859;
  assign Poutreg_new_33_ = ~n762;
  assign Poutreg_new_32_ = ~n858;
  assign Poutreg_new_31_ = ~n763;
  assign Poutreg_new_30_ = ~n857;
  assign Poutreg_new_29_ = ~n764;
  assign Poutreg_new_28_ = ~n856;
  assign Poutreg_new_27_ = ~n765;
  assign Poutreg_new_26_ = ~n855;
  assign Poutreg_new_25_ = ~n766;
  assign Poutreg_new_24_ = ~n854;
  assign Poutreg_new_23_ = ~n767;
  assign Poutreg_new_22_ = ~n853;
  assign Poutreg_new_21_ = ~n768;
  assign Poutreg_new_20_ = ~n852;
  assign Poutreg_new_19_ = ~n769;
  assign Poutreg_new_18_ = ~n851;
  assign Poutreg_new_17_ = ~n770;
  assign Poutreg_new_16_ = ~n850;
  assign Poutreg_new_15_ = ~n771;
  assign Poutreg_new_14_ = ~n848;
  assign Poutreg_new_13_ = ~n772;
  assign Poutreg_new_12_ = ~n847;
  assign Poutreg_new_11_ = ~n773;
  assign Poutreg_new_10_ = ~n846;
  assign Poutreg_new_9_ = ~n774;
  assign Poutreg_new_8_ = ~n844;
  assign Poutreg_new_7_ = ~n775;
  assign Poutreg_new_6_ = ~n843;
  assign Poutreg_new_5_ = ~n776;
  assign Poutreg_new_4_ = ~n842;
  assign Poutreg_new_3_ = ~n777;
  assign Poutreg_new_2_ = ~n840;
  assign Poutreg_new_1_ = ~n778;
  assign Poutreg_new_0_ = ~n839;
  assign Pinreg_new_55_ = ~n780;
  assign Pinreg_new_54_ = ~n781;
  assign Pinreg_new_53_ = ~n782;
  assign Pinreg_new_52_ = ~n783;
  assign Pinreg_new_51_ = ~n784;
  assign Pinreg_new_50_ = ~n785;
  assign Pinreg_new_49_ = ~n786;
  assign Pinreg_new_48_ = ~n787;
  assign Pinreg_new_47_ = ~n788;
  assign Pinreg_new_46_ = ~n789;
  assign Pinreg_new_45_ = ~n790;
  assign Pinreg_new_44_ = ~n791;
  assign Pinreg_new_43_ = ~n792;
  assign Pinreg_new_42_ = ~n793;
  assign Pinreg_new_41_ = ~n794;
  assign Pinreg_new_40_ = ~n795;
  assign Pinreg_new_39_ = ~n796;
  assign Pinreg_new_38_ = ~n797;
  assign Pinreg_new_37_ = ~n798;
  assign Pinreg_new_36_ = ~n799;
  assign Pinreg_new_35_ = ~n800;
  assign Pinreg_new_34_ = ~n801;
  assign Pinreg_new_33_ = ~n802;
  assign Pinreg_new_32_ = ~n803;
  assign Pinreg_new_31_ = ~n804;
  assign Pinreg_new_30_ = ~n805;
  assign Pinreg_new_29_ = ~n806;
  assign Pinreg_new_28_ = ~n807;
  assign Pinreg_new_27_ = ~n808;
  assign Pinreg_new_26_ = ~n809;
  assign Pinreg_new_25_ = ~n810;
  assign Pinreg_new_24_ = ~n811;
  assign Pinreg_new_23_ = ~n812;
  assign Pinreg_new_22_ = ~n813;
  assign Pinreg_new_21_ = ~n814;
  assign Pinreg_new_20_ = ~n815;
  assign Pinreg_new_19_ = ~n816;
  assign Pinreg_new_18_ = ~n817;
  assign Pinreg_new_17_ = ~n818;
  assign Pinreg_new_16_ = ~n819;
  assign Pinreg_new_15_ = ~n820;
  assign Pinreg_new_14_ = ~n821;
  assign Pinreg_new_13_ = ~n822;
  assign Pinreg_new_12_ = ~n823;
  assign Pinreg_new_11_ = ~n824;
  assign Pinreg_new_10_ = ~n825;
  assign Pinreg_new_9_ = ~n826;
  assign Pinreg_new_8_ = ~n827;
  assign Pinreg_new_7_ = ~n828;
  assign Pinreg_new_6_ = ~n829;
  assign Pinreg_new_5_ = ~n830;
  assign Pinreg_new_4_ = ~n831;
  assign Pinreg_new_3_ = ~n832;
  assign Pinreg_new_2_ = ~n833;
  assign Pinreg_new_1_ = ~n834;
  assign Pinreg_new_0_ = ~n835;
  assign Pencrypt_mode_new_0_ = ~n1799;
  assign Pdata_new_63_ = ~n1732;
  assign Pdata_new_62_ = ~n1733;
  assign Pdata_new_61_ = ~n1734;
  assign Pdata_new_60_ = ~n1735;
  assign Pdata_new_59_ = ~n1736;
  assign Pdata_new_58_ = ~n1737;
  assign Pdata_new_57_ = ~n1738;
  assign Pdata_new_56_ = ~n1739;
  assign Pdata_new_55_ = ~n1740;
  assign Pdata_new_54_ = ~n1741;
  assign Pdata_new_53_ = ~n1742;
  assign Pdata_new_52_ = ~n1743;
  assign Pdata_new_51_ = ~n1744;
  assign Pdata_new_50_ = ~n1745;
  assign Pdata_new_49_ = ~n1746;
  assign Pdata_new_48_ = ~n1747;
  assign Pdata_new_47_ = ~n1748;
  assign Pdata_new_46_ = ~n1749;
  assign Pdata_new_45_ = ~n1750;
  assign Pdata_new_44_ = ~n1751;
  assign Pdata_new_43_ = ~n1752;
  assign Pdata_new_42_ = ~n1753;
  assign Pdata_new_41_ = ~n1754;
  assign Pdata_new_40_ = ~n1755;
  assign Pdata_new_39_ = ~n1756;
  assign Pdata_new_38_ = ~n1757;
  assign Pdata_new_37_ = ~n1758;
  assign Pdata_new_36_ = ~n1759;
  assign Pdata_new_35_ = ~n1760;
  assign Pdata_new_34_ = ~n1761;
  assign Pdata_new_33_ = ~n1762;
  assign Pdata_new_32_ = ~n1763;
  assign Pdata_new_31_ = ~n1764;
  assign Pdata_new_30_ = ~n1765;
  assign Pdata_new_29_ = ~n1766;
  assign Pdata_new_28_ = ~n1767;
  assign Pdata_new_27_ = ~n1768;
  assign Pdata_new_26_ = ~n1769;
  assign Pdata_new_25_ = ~n1770;
  assign Pdata_new_24_ = ~n1771;
  assign Pdata_new_23_ = ~n1772;
  assign Pdata_new_22_ = ~n1773;
  assign Pdata_new_21_ = ~n1774;
  assign Pdata_new_20_ = ~n1775;
  assign Pdata_new_19_ = ~n1776;
  assign Pdata_new_18_ = ~n1777;
  assign Pdata_new_17_ = ~n1778;
  assign Pdata_new_16_ = ~n1779;
  assign Pdata_new_15_ = ~n1780;
  assign Pdata_new_14_ = ~n1781;
  assign Pdata_new_13_ = ~n1782;
  assign Pdata_new_12_ = ~n1783;
  assign Pdata_new_11_ = ~n1784;
  assign Pdata_new_10_ = ~n1785;
  assign Pdata_new_9_ = ~n1786;
  assign Pdata_new_8_ = ~n1787;
  assign Pdata_new_7_ = ~n1788;
  assign Pdata_new_6_ = ~n1789;
  assign Pdata_new_5_ = ~n1790;
  assign Pdata_new_4_ = ~n1791;
  assign Pdata_new_3_ = ~n1792;
  assign Pdata_new_2_ = ~n1793;
  assign Pdata_new_1_ = ~n1794;
  assign Pdata_new_0_ = ~n1795;
  assign Pcount_new_3_ = ~n779;
  assign Pcount_new_2_ = ~n1796;
  assign Pcount_new_1_ = ~n1797;
  assign Pcount_new_0_ = ~n1403;
  assign PD_new_27_ = ~n1524;
  assign PD_new_26_ = ~n1528;
  assign PD_new_25_ = ~n1532;
  assign PD_new_24_ = ~n1536;
  assign PD_new_23_ = ~n1540;
  assign PD_new_22_ = ~n1544;
  assign PD_new_21_ = ~n1548;
  assign PD_new_20_ = ~n1552;
  assign PD_new_19_ = ~n1556;
  assign PD_new_18_ = ~n1560;
  assign PD_new_17_ = ~n1564;
  assign PD_new_16_ = ~n1568;
  assign PD_new_15_ = ~n1572;
  assign PD_new_14_ = ~n1576;
  assign PD_new_13_ = ~n1580;
  assign PD_new_12_ = ~n1584;
  assign PD_new_11_ = ~n1588;
  assign PD_new_10_ = ~n1592;
  assign PD_new_9_ = ~n1596;
  assign PD_new_8_ = ~n1600;
  assign PD_new_7_ = ~n1604;
  assign PD_new_6_ = ~n1608;
  assign PD_new_5_ = ~n1612;
  assign PD_new_4_ = ~n1616;
  assign PD_new_3_ = ~n1620;
  assign PD_new_2_ = ~n1624;
  assign PD_new_1_ = ~n1628;
  assign PD_new_0_ = ~n1632;
  assign PC_new_27_ = ~n1412;
  assign PC_new_26_ = ~n1416;
  assign PC_new_25_ = ~n1420;
  assign PC_new_24_ = ~n1424;
  assign PC_new_23_ = ~n1428;
  assign PC_new_22_ = ~n1432;
  assign PC_new_21_ = ~n1436;
  assign PC_new_20_ = ~n1440;
  assign PC_new_19_ = ~n1444;
  assign PC_new_18_ = ~n1448;
  assign PC_new_17_ = ~n1452;
  assign PC_new_16_ = ~n1456;
  assign PC_new_15_ = ~n1460;
  assign PC_new_14_ = ~n1464;
  assign PC_new_13_ = ~n1468;
  assign PC_new_12_ = ~n1472;
  assign PC_new_11_ = ~n1476;
  assign PC_new_10_ = ~n1480;
  assign PC_new_9_ = ~n1484;
  assign PC_new_8_ = ~n1488;
  assign PC_new_7_ = ~n1492;
  assign PC_new_6_ = ~n1496;
  assign PC_new_5_ = ~n1500;
  assign PC_new_4_ = ~n1504;
  assign PC_new_3_ = ~n1508;
  assign PC_new_2_ = ~n1512;
  assign PC_new_1_ = ~n1516;
  assign PC_new_0_ = ~n1520;
  assign n746 = ~Pcount_3_ | n1648;
  assign n747 = (~Poutreg_63_ | Pcount_0_) & (n746 | n899);
  assign n748 = (~Poutreg_61_ | Pcount_0_) & (n746 | n931);
  assign n749 = (~Poutreg_59_ | Pcount_0_) & (n746 | n948);
  assign n750 = (~Poutreg_57_ | Pcount_0_) & (n746 | n976);
  assign n751 = (~Poutreg_55_ | Pcount_0_) & n986;
  assign n752 = (~Poutreg_53_ | Pcount_0_) & n1024;
  assign n753 = (~Poutreg_51_ | Pcount_0_) & n1037;
  assign n754 = (~Poutreg_49_ | Pcount_0_) & n1059;
  assign n755 = (~Poutreg_47_ | Pcount_0_) & n1099;
  assign n756 = (~Poutreg_45_ | Pcount_0_) & n1126;
  assign n757 = (~Poutreg_43_ | Pcount_0_) & n1135;
  assign n758 = (~Poutreg_41_ | Pcount_0_) & n1144;
  assign n759 = (~Poutreg_39_ | Pcount_0_) & n1157;
  assign n760 = (~Poutreg_37_ | Pcount_0_) & n1167;
  assign n761 = (~Poutreg_35_ | Pcount_0_) & n1197;
  assign n762 = (~Poutreg_33_ | Pcount_0_) & n1203;
  assign n763 = (~Poutreg_31_ | Pcount_0_) & n1216;
  assign n764 = (~Poutreg_29_ | Pcount_0_) & n1233;
  assign n765 = (~Poutreg_27_ | Pcount_0_) & n1242;
  assign n766 = (~Poutreg_25_ | Pcount_0_) & n1248;
  assign n767 = (~Poutreg_23_ | Pcount_0_) & n1290;
  assign n768 = (~Poutreg_21_ | Pcount_0_) & n1305;
  assign n769 = (~Poutreg_19_ | Pcount_0_) & n1313;
  assign n770 = (~Poutreg_17_ | Pcount_0_) & n1329;
  assign n771 = (~Poutreg_15_ | Pcount_0_) & n1336;
  assign n772 = (~Poutreg_13_ | Pcount_0_) & n1345;
  assign n773 = (~Poutreg_11_ | Pcount_0_) & n1354;
  assign n774 = (~Poutreg_9_ | Pcount_0_) & n1363;
  assign n775 = (~Poutreg_7_ | Pcount_0_) & n1374;
  assign n776 = (~Poutreg_5_ | Pcount_0_) & n1379;
  assign n777 = (~Poutreg_3_ | Pcount_0_) & n1392;
  assign n778 = (~Poutreg_1_ | Pcount_0_) & n1401;
  assign n779 = (n1404 | n1407) & (~Pcount_3_ | n1406);
  assign n780 = (~Pinreg_55_ | Pcount_0_) & (~Pinreg_47_ | n869);
  assign n781 = (~Pinreg_54_ | Pcount_0_) & (~Pinreg_46_ | n869);
  assign n782 = (~Pinreg_53_ | Pcount_0_) & (~Pinreg_45_ | n869);
  assign n783 = (~Pinreg_52_ | Pcount_0_) & (~Pinreg_44_ | n869);
  assign n784 = (~Pinreg_51_ | Pcount_0_) & (~Pinreg_43_ | n869);
  assign n785 = (~Pinreg_50_ | Pcount_0_) & (~Pinreg_42_ | n869);
  assign n786 = (~Pinreg_49_ | Pcount_0_) & (~Pinreg_41_ | n869);
  assign n787 = (~Pinreg_48_ | Pcount_0_) & (~Pinreg_40_ | n869);
  assign n788 = (~Pinreg_47_ | Pcount_0_) & (~Pinreg_39_ | n869);
  assign n789 = (~Pinreg_46_ | Pcount_0_) & (~Pinreg_38_ | n869);
  assign n790 = (~Pinreg_45_ | Pcount_0_) & (~Pinreg_37_ | n869);
  assign n791 = (~Pinreg_44_ | Pcount_0_) & (~Pinreg_36_ | n869);
  assign n792 = (~Pinreg_43_ | Pcount_0_) & (~Pinreg_35_ | n869);
  assign n793 = (~Pinreg_42_ | Pcount_0_) & (~Pinreg_34_ | n869);
  assign n794 = (~Pinreg_41_ | Pcount_0_) & (~Pinreg_33_ | n869);
  assign n795 = (~Pinreg_40_ | Pcount_0_) & (~Pinreg_32_ | n869);
  assign n796 = (~Pinreg_39_ | Pcount_0_) & (~Pinreg_31_ | n869);
  assign n797 = (~Pinreg_38_ | Pcount_0_) & (~Pinreg_30_ | n869);
  assign n798 = (~Pinreg_37_ | Pcount_0_) & (~Pinreg_29_ | n869);
  assign n799 = (~Pinreg_36_ | Pcount_0_) & (~Pinreg_28_ | n869);
  assign n800 = (~Pinreg_35_ | Pcount_0_) & (~Pinreg_27_ | n869);
  assign n801 = (~Pinreg_34_ | Pcount_0_) & (~Pinreg_26_ | n869);
  assign n802 = (~Pinreg_33_ | Pcount_0_) & (~Pinreg_25_ | n869);
  assign n803 = (~Pinreg_32_ | Pcount_0_) & (~Pinreg_24_ | n869);
  assign n804 = (~Pinreg_31_ | Pcount_0_) & (~Pinreg_23_ | n869);
  assign n805 = (~Pinreg_30_ | Pcount_0_) & (~Pinreg_22_ | n869);
  assign n806 = (~Pinreg_29_ | Pcount_0_) & (~Pinreg_21_ | n869);
  assign n807 = (~Pinreg_28_ | Pcount_0_) & (~Pinreg_20_ | n869);
  assign n808 = (~Pinreg_27_ | Pcount_0_) & (~Pinreg_19_ | n869);
  assign n809 = (~Pinreg_26_ | Pcount_0_) & (~Pinreg_18_ | n869);
  assign n810 = (~Pinreg_25_ | Pcount_0_) & (~Pinreg_17_ | n869);
  assign n811 = (~Pinreg_24_ | Pcount_0_) & (~Pinreg_16_ | n869);
  assign n812 = (~Pinreg_23_ | Pcount_0_) & (~Pinreg_15_ | n869);
  assign n813 = (~Pinreg_22_ | Pcount_0_) & (~Pinreg_14_ | n869);
  assign n814 = (~Pinreg_21_ | Pcount_0_) & (~Pinreg_13_ | n869);
  assign n815 = (~Pinreg_20_ | Pcount_0_) & (~Pinreg_12_ | n869);
  assign n816 = (~Pinreg_19_ | Pcount_0_) & (~Pinreg_11_ | n869);
  assign n817 = (~Pinreg_18_ | Pcount_0_) & (~Pinreg_10_ | n869);
  assign n818 = (~Pinreg_17_ | Pcount_0_) & (~Pinreg_9_ | n869);
  assign n819 = (~Pinreg_16_ | Pcount_0_) & (~Pinreg_8_ | n869);
  assign n820 = (~Pinreg_15_ | Pcount_0_) & (~Pinreg_7_ | n869);
  assign n821 = (~Pinreg_14_ | Pcount_0_) & (~Pinreg_6_ | n869);
  assign n822 = (~Pinreg_13_ | Pcount_0_) & (~Pinreg_5_ | n869);
  assign n823 = (~Pinreg_12_ | Pcount_0_) & (~Pinreg_4_ | n869);
  assign n824 = (~Pinreg_11_ | Pcount_0_) & (~Pinreg_3_ | n869);
  assign n825 = (~Pinreg_10_ | Pcount_0_) & (~Pinreg_2_ | n869);
  assign n826 = (~Pinreg_9_ | Pcount_0_) & (~Pinreg_1_ | n869);
  assign n827 = (~Pinreg_8_ | Pcount_0_) & (~Pinreg_0_ | n869);
  assign n828 = (~Pinreg_7_ | Pcount_0_) & (~Pdata_in_7_ | n869);
  assign n829 = (~Pinreg_6_ | Pcount_0_) & (~Pdata_in_6_ | n869);
  assign n830 = (~Pinreg_5_ | Pcount_0_) & (~Pdata_in_5_ | n869);
  assign n831 = (~Pinreg_4_ | Pcount_0_) & (~Pdata_in_4_ | n869);
  assign n832 = (~Pinreg_3_ | Pcount_0_) & (~Pdata_in_3_ | n869);
  assign n833 = (~Pinreg_2_ | Pcount_0_) & (~Pdata_in_2_ | n869);
  assign n834 = (~Pinreg_1_ | Pcount_0_) & (~Pdata_in_1_ | n869);
  assign n835 = (~Pinreg_0_ | Pcount_0_) & (~Pdata_in_0_ | n869);
  assign n836 = (~Poutreg_56_ | Pcount_0_) & (~Pdata_32_ | n746);
  assign n837 = Pload_key_0_ & ~n746;
  assign n838 = (~Pdata_49_ | n746) & n1025;
  assign n839 = (~Pdata_39_ | n746) & n1402;
  assign n840 = (~Pdata_47_ | n746) & n1393;
  assign n841 = (~Poutreg_58_ | Pcount_0_) & (~Pdata_40_ | n746);
  assign n842 = (~Pdata_55_ | n746) & n1380;
  assign n843 = (~Pdata_63_ | n746) & n1375;
  assign n844 = (~Pdata_38_ | n746) & n1364;
  assign n845 = (~Poutreg_60_ | Pcount_0_) & (~Pdata_48_ | n746);
  assign n846 = (~Pdata_46_ | n746) & n1355;
  assign n847 = (~Pdata_54_ | n746) & n1346;
  assign n848 = (~Pdata_62_ | n746) & n1337;
  assign n849 = (~Poutreg_62_ | Pcount_0_) & (~Pdata_56_ | n746);
  assign n850 = (~Pdata_37_ | n746) & n1330;
  assign n851 = (~Pdata_45_ | n746) & n1314;
  assign n852 = (~Pdata_53_ | n746) & n1306;
  assign n853 = (~Pdata_61_ | n746) & n1291;
  assign n854 = (~Pdata_36_ | n746) & n1249;
  assign n855 = (~Pdata_44_ | n746) & n1243;
  assign n856 = (~Pdata_52_ | n746) & n1234;
  assign n857 = (~Pdata_60_ | n746) & n1217;
  assign n858 = (~Pdata_35_ | n746) & n1204;
  assign n859 = (~Pdata_43_ | n746) & n1198;
  assign n860 = (~Pdata_51_ | n746) & n1168;
  assign n861 = (~Pdata_59_ | n746) & n1158;
  assign n862 = (~Pdata_34_ | n746) & n1145;
  assign n863 = (~Pdata_42_ | n746) & n1136;
  assign n864 = (~Pdata_50_ | n746) & n1127;
  assign n865 = (~Pdata_58_ | n746) & n1100;
  assign n866 = (~Pdata_33_ | n746) & n1060;
  assign n867 = (~Pdata_41_ | n746) & n1038;
  assign n868 = (~Pdata_57_ | n746) & n987;
  assign n869 = ~Pcount_0_ | ~n746;
  assign n870 = (~n893 | ~n1140) & (~n892 | ~n896);
  assign n871 = (~n878 | ~n892) & (~n1140 | ~n1649);
  assign n872 = ~Pdata_49_ ^ ~PD_2_;
  assign n873 = (n871 | ~n1394) & (n870 | n872);
  assign n874 = n1800 & (~n1651 | (~n877 & n885));
  assign n875 = n873 & n874 & (~n1394 | ~n1652);
  assign n876 = n1398 & ~n1633;
  assign n877 = n1394 & n1650;
  assign n878 = ~n887 & n1634;
  assign n879 = n876 & (n877 | (n878 & ~n890));
  assign n880 = ~n1651 | n890 | ~n1649;
  assign n881 = n1633 | n1653;
  assign n882 = ~n879 & n880 & (n881 | ~n1395);
  assign n883 = ~n1652 | n872 | n1397;
  assign n884 = (n1311 | ~n1650) & (~n878 | n1654);
  assign n885 = ~n872 | ~n896;
  assign n886 = n883 & n884 & (n885 | ~n1140);
  assign n887 = ~Pdata_50_ ^ ~PD_8_;
  assign n888 = ~n1397 ^ ~n1634;
  assign n889 = ~n1651 | n887 | n888;
  assign n890 = ~n872 | n1397;
  assign n891 = n890 | ~n1651;
  assign n892 = n1398 & n1633;
  assign n893 = ~n1397 & n1650;
  assign n894 = n1650 | n1649;
  assign n895 = n892 & (n893 | (n872 & n894));
  assign n896 = n1395 & ~n1397;
  assign n897 = n1140 | n876;
  assign n898 = ~n872 & (~n889 | (n896 & n897));
  assign n899 = ~Pdata_24_ ^ ~n1978;
  assign n900 = n914 & ~n920;
  assign n901 = ~n1338 & ~n912 & ~n916;
  assign n902 = n900 & ~n1926 & (n901 | ~n906);
  assign n903 = ~n902 & (~n912 | ~n918 | ~n1721);
  assign n904 = (~n934 | n938) & (~n1338 | ~n1720);
  assign n905 = n903 & n904 & (~n926 | ~n1656);
  assign n906 = ~Pdata_36_ ^ ~PC_4_;
  assign n907 = (~n926 | ~n1338) & (n906 | ~n1657);
  assign n908 = n1655 | ~n914 | ~n932;
  assign n909 = ~n934 | ~n1656;
  assign n910 = n908 & n909 & (n907 | ~n935);
  assign n911 = n906 | ~n912;
  assign n912 = ~Pdata_35_ ^ ~PC_0_;
  assign n913 = n911 & (~n906 | n912);
  assign n914 = ~Pdata_63_ ^ ~PC_13_;
  assign n915 = ~n900 & (n914 | ~n920);
  assign n916 = ~Pdata_32_ ^ ~PC_16_;
  assign n917 = ~n906 & n916;
  assign n918 = ~n916 & ~n920;
  assign n919 = ~n906 & n918 & (~n912 | ~n914);
  assign n920 = ~Pdata_34_ ^ ~PC_23_;
  assign n921 = ~n912 & n916;
  assign n922 = ~n914 & n920 & (n917 | n921);
  assign n923 = (~n920 | ~n921) & (n913 | ~n918);
  assign n924 = n1338 & n934;
  assign n925 = n924 & ~n912 & n918;
  assign n926 = ~n906 & ~n914;
  assign n927 = n901 & ~n920 & n926;
  assign n928 = ~n914 | n923 | ~n1338;
  assign n929 = (~n926 | n1659) & (~n932 | ~n1658);
  assign n930 = n929 & n928 & n905 & n910 & ~n1662 & ~n1924;
  assign n931 = ~n930 ^ ~Pdata_16_;
  assign n932 = n912 & n906;
  assign n933 = n932 & n900 & n916;
  assign n934 = n906 & ~n914;
  assign n935 = n920 & n916 & n912;
  assign n936 = ~n1338 & (n933 | (n934 & n935));
  assign n937 = n1655 | n911 | ~n914;
  assign n938 = n912 | n1655;
  assign n939 = ~n936 & n937 & (~n926 | n938);
  assign n940 = (n906 | ~n921) & (n913 | n916);
  assign n941 = n916 | ~n900 | ~n906;
  assign n942 = ~n926 | n1655;
  assign n943 = (n906 & (~n920 | ~n924)) | (n920 & ~n924);
  assign n944 = n941 & n942 & (~n916 | n943);
  assign n945 = n1803 & (~n920 | n940 | ~n1657);
  assign n946 = n905 & n1341 & (~n906 | n1659);
  assign n947 = n945 & (~n912 | n944) & n946;
  assign n948 = ~n947 ^ ~Pdata_8_;
  assign n949 = n980 | n1635;
  assign n950 = ~n956 | n1030;
  assign n951 = n957 | ~n980;
  assign n952 = (n949 | n950) & (n951 | ~n1163);
  assign n953 = (n983 | n1663) & (n952 | n958);
  assign n954 = n949 | n981;
  assign n955 = n953 & (n954 | ~n1161);
  assign n956 = ~Pdata_43_ ^ ~PC_15_;
  assign n957 = n956 | ~n1159;
  assign n958 = ~Pdata_48_ ^ ~PC_1_;
  assign n959 = (n956 | ~n961) & (n957 | n958);
  assign n960 = n956 & ~n958 & n1159;
  assign n961 = n958 & ~n1159;
  assign n962 = ~n1664 & (n960 | (n956 & n961));
  assign n963 = n955 & ~n962 & (n954 | n959);
  assign n964 = (~n960 | n1663) & (~n961 | n1667);
  assign n965 = n1805 & (n958 | ~n1635 | n1666);
  assign n966 = n964 & n965;
  assign n967 = n1804 & (n949 | ~n981 | n983);
  assign n968 = n1159 | n958;
  assign n969 = n967 & (n968 | ~n1724);
  assign n970 = ~n956 ^ ~n1635;
  assign n971 = n1030 | n958;
  assign n972 = n981 | ~n1635;
  assign n973 = (n970 | n971) & (n972 | ~n1161);
  assign n974 = ~n956 | n968;
  assign n975 = n974 & n950 & (n957 | n958);
  assign n976 = ~Pdata_0_ ^ ~n1979;
  assign n977 = (~n958 | n1669) & (n968 | n1667);
  assign n978 = n1809 & (~n960 | ~n981 | n1665);
  assign n979 = n977 & n978;
  assign n980 = ~Pdata_46_ ^ ~PC_19_;
  assign n981 = ~Pdata_44_ ^ ~PC_6_;
  assign n982 = n980 & (~n973 | (n981 & ~n983));
  assign n983 = n957 | ~n958;
  assign n984 = n954 | n983;
  assign n985 = n956 & (~n1808 | (~n1159 & ~n1663));
  assign n986 = (n746 | n1810) & (~Poutreg_63_ | n869);
  assign n987 = (~Poutreg_62_ | n869) & (~Poutreg_54_ | Pcount_0_);
  assign n988 = (n1017 | n1236) & (~n996 | ~n997);
  assign n989 = ~n1017 | n1149;
  assign n990 = n988 & (n989 | ~n1039);
  assign n991 = ~n993 | ~n1146;
  assign n992 = ~n1039 | n989 | n991;
  assign n993 = ~Pdata_36_ ^ ~PC_27_;
  assign n994 = n1004 | ~n1146;
  assign n995 = ~n997 | n993 | n994;
  assign n996 = ~n1054 & ~n1636;
  assign n997 = n1017 & n1149;
  assign n998 = n996 & (~n1022 | (n997 & ~n1670));
  assign n999 = ~n998 & n992 & n995;
  assign n1000 = n1813 & (~n1050 | ~n1146 | n1671);
  assign n1001 = n1670 | n1017;
  assign n1002 = n1004 | ~n1149;
  assign n1003 = n999 & n1000 & (n1001 | n1002);
  assign n1004 = ~n1054 | n1636;
  assign n1005 = n993 | ~n1146;
  assign n1006 = (n1005 | ~n1050) & (n1004 | ~n1049);
  assign n1007 = ~n993 | n1018 | n1056;
  assign n1008 = n1001 | n1236;
  assign n1009 = n1007 & n1008 & (n1006 | ~n1051);
  assign n1010 = (n1042 | ~n1049) & (n1004 | n1053);
  assign n1011 = n1811 & (~n993 | n1013 | n1056);
  assign n1012 = n1010 & n1011;
  assign n1013 = ~n996 | ~n1149;
  assign n1014 = n1012 & n1009 & (n1001 | n1013);
  assign n1015 = n1636 | n989 | ~n1146;
  assign n1016 = (~n997 | ~n1054) & (~n996 | ~n1051);
  assign n1017 = ~Pdata_37_ ^ ~PC_14_;
  assign n1018 = ~n1050 | ~n1149;
  assign n1019 = n1015 & n1016 & (n1017 | n1018);
  assign n1020 = n1814 & (n990 | n1005);
  assign n1021 = n1003 & n1014 & (~n993 | n1019);
  assign n1022 = n1149 | n1001;
  assign n1023 = n1020 & n1021 & (n1004 | n1022);
  assign n1024 = (n746 | n1815) & (~Poutreg_61_ | n869);
  assign n1025 = (~Poutreg_60_ | n869) & (~Poutreg_52_ | Pcount_0_);
  assign n1026 = ~n981 | ~n1159 | n970 | n980;
  assign n1027 = (n957 | n972) & (n950 | n1665);
  assign n1028 = n1026 & n1027 & (n951 | n981);
  assign n1029 = ~n1163 | n957 | n980;
  assign n1030 = ~n981 | n1159;
  assign n1031 = n1029 & (n970 | ~n980 | n1030);
  assign n1032 = (n958 & n1031) | (n1028 & (~n958 | n1031));
  assign n1033 = n969 & n966;
  assign n1034 = (n954 | ~n956) & (n951 | n972);
  assign n1035 = n1165 & (~n1161 | n1665);
  assign n1036 = n1035 & n955 & n1033 & n1032 & n979 & n1034;
  assign n1037 = (n746 | n1816) & (~Poutreg_59_ | n869);
  assign n1038 = (~Poutreg_58_ | n869) & (~Poutreg_50_ | Pcount_0_);
  assign n1039 = n1054 & n1636;
  assign n1040 = n1039 & (~n1022 | (n997 & ~n1670));
  assign n1041 = ~n1051 | n993 | n994;
  assign n1042 = ~n1017 | n1018;
  assign n1043 = ~n1040 & n1041 & (n991 | n1042);
  assign n1044 = n1004 & ~n1050;
  assign n1045 = n989 | n991 | n1044;
  assign n1046 = n1236 & ~n996 & n1146;
  assign n1047 = n1002 & ~n1146;
  assign n1048 = n1046 | n1047 | n993 | ~n1017;
  assign n1049 = n993 & ~n1146;
  assign n1050 = ~n1054 & n1636;
  assign n1051 = ~n1017 & ~n1149;
  assign n1052 = n1049 & (~n990 | (n1050 & n1051));
  assign n1053 = n1146 | n1671;
  assign n1054 = ~Pdata_39_ ^ ~PC_20_;
  assign n1055 = n1053 | n1054;
  assign n1056 = n1017 | ~n1146;
  assign n1057 = n1018 & ~n1637;
  assign n1058 = n1056 | n1057;
  assign n1059 = (n746 | n1817) & (~Poutreg_57_ | n869);
  assign n1060 = (~Poutreg_56_ | n869) & (~Poutreg_48_ | Pcount_0_);
  assign n1061 = ~Pdata_63_ ^ ~PD_0_;
  assign n1062 = ~Pdata_61_ ^ ~PD_21_;
  assign n1063 = ~n1087 | ~n1672;
  assign n1064 = n1063 | n1061 | n1062;
  assign n1065 = n1078 | n1076 | n1673;
  assign n1066 = n1078 | n1061 | ~n1062;
  assign n1067 = n1065 & ~n1929 & (n1063 | n1066);
  assign n1068 = n1930 & (n1078 | n1083 | ~n1352);
  assign n1069 = (~n1349 | n1676) & (n1073 | n1818);
  assign n1070 = n1069 & n1068 & n1067;
  assign n1071 = ~n1062 | n1087 | n1222;
  assign n1072 = n1061 | ~n1078;
  assign n1073 = n1062 | n1083;
  assign n1074 = n1078 | ~n1222;
  assign n1075 = (n1073 | n1074) & (n1071 | n1072);
  assign n1076 = ~Pdata_59_ ^ ~PD_17_;
  assign n1077 = ~n1078 | ~n1222;
  assign n1078 = ~Pdata_32_ ^ ~PD_3_;
  assign n1079 = (n1076 | n1077) & (n1078 | ~n1351);
  assign n1080 = ~n1061 | n1074 | ~n1076 | ~n1349;
  assign n1081 = n1674 | n1220;
  assign n1082 = n1080 & n1081 & (n1079 | n1073);
  assign n1083 = n1061 | n1087;
  assign n1084 = n1077 | n1076 | n1083;
  assign n1085 = ~n1076 | n1077 | ~n1675;
  assign n1086 = ~n1672 | n1073 | n1078;
  assign n1087 = ~Pdata_60_ ^ ~PD_13_;
  assign n1088 = n1062 & (~n1084 | (n1087 & ~n1676));
  assign n1089 = ~n1349 | n1061 | n1076;
  assign n1090 = (~n1061 | n1063) & n1089;
  assign n1091 = ~n1352 | n1061 | ~n1087;
  assign n1092 = n1066 | ~n1351;
  assign n1093 = ~n1061 | n1062 | n1063;
  assign n1094 = n1819 & (~n1078 | (n1090 & ~n1950));
  assign n1095 = (n1062 & n1680) | (n1676 & (~n1062 | n1680));
  assign n1096 = (n1075 | ~n1076) & (n1066 | ~n1087);
  assign n1097 = n1678 & n1082;
  assign n1098 = n1070 & n1094 & n1093 & n1091 & n1092 & n1095 & n1096 & n1097;
  assign n1099 = (n746 | n1820) & (~Poutreg_55_ | n869);
  assign n1100 = (~Poutreg_54_ | n869) & (~Poutreg_46_ | Pcount_0_);
  assign n1101 = ~n1102 | n1120;
  assign n1102 = ~Pdata_55_ ^ ~PD_4_;
  assign n1103 = n1101 & (n1102 | ~n1120);
  assign n1104 = ~n1638 & ~n1639;
  assign n1105 = ~n1102 & n1682;
  assign n1106 = n1104 & (n1105 | ~n1822);
  assign n1107 = ~n1932 & (~n1105 | ~n1132 | ~n1201);
  assign n1108 = n1823 & n1824 & (n1130 | n1117);
  assign n1109 = n1201 | n1207;
  assign n1110 = n1107 & n1108 & (n1109 | ~n1683);
  assign n1111 = n1821 & (n1130 | (~n1105 & n1822));
  assign n1112 = n1102 | n1119;
  assign n1113 = n1111 & (n1112 | n1109);
  assign n1114 = ~n1201 | n1207 | ~n1683;
  assign n1115 = (n1109 | n1685) & (n1130 | n1684);
  assign n1116 = n1201 | n1211;
  assign n1117 = n1133 | n1101;
  assign n1118 = n1114 & n1115 & (n1116 | n1117);
  assign n1119 = ~n1120 | n1133;
  assign n1120 = ~Pdata_51_ ^ ~PD_1_;
  assign n1121 = n1119 & (n1120 | ~n1133);
  assign n1122 = n1118 & n1113;
  assign n1123 = n1931 & (~n1201 | (n1825 & n1826));
  assign n1124 = n1828 & (n1211 | n1685);
  assign n1125 = n1124 & n1123 & n1110 & n1122;
  assign n1126 = (n746 | n1829) & (~Poutreg_53_ | n869);
  assign n1127 = (~Poutreg_52_ | n869) & (~Poutreg_44_ | Pcount_0_);
  assign n1128 = n1830 & (n1109 | (n1822 & n1684));
  assign n1129 = n1133 | ~n1681;
  assign n1130 = ~n1201 | n1211;
  assign n1131 = n1128 & (n1129 | n1130);
  assign n1132 = ~n1638 & n1639;
  assign n1133 = ~Pdata_54_ ^ ~PD_16_;
  assign n1134 = n1132 & (~n1684 | (~n1103 & n1133));
  assign n1135 = (n746 | n1834) & (~Poutreg_51_ | n869);
  assign n1136 = (~Poutreg_50_ | n869) & (~Poutreg_42_ | Pcount_0_);
  assign n1137 = ~n1649 | n890 | ~n1140;
  assign n1138 = (~n878 | n881) & (~n1650 | n1654);
  assign n1139 = n1137 & (~n876 | n885) & n1138;
  assign n1140 = ~n1398 & n1633;
  assign n1141 = n878 & n1140 & n890;
  assign n1142 = n1649 & n892;
  assign n1143 = n1142 & ~n1397;
  assign n1144 = (~Poutreg_49_ | n869) & (n746 | ~n1996);
  assign n1145 = (~Poutreg_48_ | n869) & (~Poutreg_40_ | Pcount_0_);
  assign n1146 = ~Pdata_35_ ^ ~PC_2_;
  assign n1147 = ~n1017 | ~n1039;
  assign n1148 = n994 & (n1146 | (~n996 & n1147));
  assign n1149 = ~Pdata_40_ ^ ~PC_9_;
  assign n1150 = (n989 | n1146) & (n1149 | n1056);
  assign n1151 = (n1148 | ~n1149) & (n1054 | n1150);
  assign n1152 = (~n1039 | n1056) & n1151;
  assign n1153 = n1001 | n1018;
  assign n1154 = (n1146 | n1687) & (~n993 | n1152);
  assign n1155 = n1835 & (n994 | n1671);
  assign n1156 = n1155 & n1153 & n1009 & n1043 & n1003 & n1154;
  assign n1157 = (n746 | n1836) & (~Poutreg_47_ | n869);
  assign n1158 = (~Poutreg_46_ | n869) & (~Poutreg_38_ | Pcount_0_);
  assign n1159 = ~Pdata_47_ ^ ~PC_12_;
  assign n1160 = n980 & (~n950 | (~n981 & n1159));
  assign n1161 = n1159 & n956 & n958;
  assign n1162 = n981 & (~n951 | (~n980 & n1161));
  assign n1163 = n981 & n1635;
  assign n1164 = n960 & (~n954 | (n980 & n1163));
  assign n1165 = ~n961 | n1663;
  assign n1166 = n1165 | n956;
  assign n1167 = (n746 | n1837) & (~Poutreg_45_ | n869);
  assign n1168 = (~Poutreg_44_ | n869) & (~Poutreg_36_ | Pcount_0_);
  assign n1169 = (~n1292 | ~n1726) & (n1177 | ~n1358);
  assign n1170 = n1367 | ~n1642;
  assign n1171 = n1169 & (n1170 | ~n1303);
  assign n1172 = ~n1190 & n1641;
  assign n1173 = ~n1299 & ~n1642;
  assign n1174 = ~n1292 & ~n1300;
  assign n1175 = n1172 & (~n1170 | (n1173 & n1174));
  assign n1176 = n1689 | ~n1296 | ~n1303;
  assign n1177 = n1689 | ~n1690;
  assign n1178 = ~n1175 & n1176 & (n1177 | ~n1295);
  assign n1179 = n1292 | ~n1300;
  assign n1180 = (~n1172 | ~n1174) & (n1179 | ~n1358);
  assign n1181 = ~n1292 | n1641 | ~n1691;
  assign n1182 = n1177 | ~n1303;
  assign n1183 = n1181 & n1182 & (n1180 | ~n1298);
  assign n1184 = (~n1296 | ~n1358) & (~n1295 | ~n1690);
  assign n1185 = ~n1690 | ~n1172 | ~n1302;
  assign n1186 = ~n1173 | n1692;
  assign n1187 = n1185 & n1186 & (n1184 | ~n1298);
  assign n1188 = ~n1302 | ~n1358;
  assign n1189 = n1694 | ~n1298 | ~n1300;
  assign n1190 = ~Pdata_57_ ^ ~PD_10_;
  assign n1191 = n1188 & n1189 & (n1190 | ~n1361);
  assign n1192 = n1942 & (n1694 | n1695);
  assign n1193 = n1178 & n1171;
  assign n1194 = (n1191 | ~n1292) & (~n1299 | n1692);
  assign n1195 = (n1370 | ~n1641) & (~n1295 | n1693);
  assign n1196 = n1195 & n1187 & n1183 & n1192 & n1193 & n1194;
  assign n1197 = (n746 | n1838) & (~Poutreg_43_ | n869);
  assign n1198 = (~Poutreg_42_ | n869) & (~Poutreg_34_ | Pcount_0_);
  assign n1199 = (~n1681 | ~n1696) & (n1103 | ~n1640);
  assign n1200 = ~n1102 | ~n1120;
  assign n1201 = ~Pdata_53_ ^ ~PD_22_;
  assign n1202 = n1200 & ~n1681 & (n1102 | n1201);
  assign n1203 = (n746 | n1840) & (~Poutreg_41_ | n869);
  assign n1204 = (~Poutreg_40_ | n869) & (~Poutreg_32_ | Pcount_0_);
  assign n1205 = n1639 | n1685;
  assign n1206 = n1841 & n1842 & (n1211 | ~n1683);
  assign n1207 = ~n1638 | ~n1639;
  assign n1208 = n1205 & n1206 & (n1112 | n1207);
  assign n1209 = ~n1132 | n1102 | n1121;
  assign n1210 = (~n1681 | n1686) & (n1638 | ~n1683);
  assign n1211 = ~n1638 | n1639;
  assign n1212 = n1209 & n1210 & (n1103 | n1211);
  assign n1213 = (~n1201 & n1212) | (n1208 & (n1201 | n1212));
  assign n1214 = n1118 & (n1129 | n1109);
  assign n1215 = n1110 & n1214 & n1213 & n1131;
  assign n1216 = (n746 | n1843) & (~Poutreg_39_ | n869);
  assign n1217 = (~Poutreg_38_ | n869) & (~Poutreg_30_ | Pcount_0_);
  assign n1218 = n1066 | n1076 | n1087 | ~n1222;
  assign n1219 = n1946 & (n1078 | ~n1672 | ~n1675);
  assign n1220 = ~n1078 | ~n1352;
  assign n1221 = n1218 & n1219 & (n1220 | ~n1677);
  assign n1222 = ~Pdata_62_ ^ ~PD_7_;
  assign n1223 = n1074 & (~n1078 | n1222);
  assign n1224 = n1073 | ~n1351;
  assign n1225 = n1061 | ~n1087 | ~n1222 | n1643;
  assign n1226 = n1224 & (~n1062 | n1063) & n1225;
  assign n1227 = n1643 | n1223 | n1674;
  assign n1228 = ~n1677 | n1222 | ~n1643;
  assign n1229 = (n1078 & n1226) | (n1091 & (~n1078 | n1226));
  assign n1230 = n1061 | n1679;
  assign n1231 = (~n1087 | n1092) & (n1074 | n1089);
  assign n1232 = n1067 & n1221 & n1229 & n1227 & n1228 & n1097 & n1230 & n1231;
  assign n1233 = (n746 | n1844) & (~Poutreg_37_ | n869);
  assign n1234 = (~Poutreg_36_ | n869) & (~Poutreg_28_ | Pcount_0_);
  assign n1235 = n1149 | n1044 | ~n1146;
  assign n1236 = ~n1039 | ~n1149;
  assign n1237 = n1235 & (~n996 | n1146) & n1236;
  assign n1238 = n1949 & (~n1017 | n1057 | n1146);
  assign n1239 = ~n993 | n1017 | n1237;
  assign n1240 = (n1022 | ~n1050) & (~n1670 | n1687);
  assign n1241 = n1240 & n1012 & n1238 & n1043 & n1003 & n1239;
  assign n1242 = (n746 | n1845) & (~Poutreg_35_ | n869);
  assign n1243 = (~Poutreg_34_ | n869) & (~Poutreg_26_ | Pcount_0_);
  assign n1244 = n1846 & (~n1078 | n1093) & ~n1951;
  assign n1245 = (n1222 | n1089) & (n1062 | n1680);
  assign n1246 = n1225 & n1679 & (n1083 | n1220);
  assign n1247 = n1246 & n1244 & n1221 & n1070 & n1082 & n1245;
  assign n1248 = (n746 | n1847) & (~Poutreg_33_ | n869);
  assign n1249 = (~Poutreg_32_ | n869) & (~Poutreg_24_ | Pcount_0_);
  assign n1250 = n1276 | n1382;
  assign n1251 = ~n1281 | ~n1285;
  assign n1252 = (~n1258 | ~n1259) & (n1250 | n1251);
  assign n1253 = n1697 | n1251 | ~n1276;
  assign n1254 = n1276 | n1265 | n1384;
  assign n1255 = n1253 & n1254 & (n1252 | ~n1317);
  assign n1256 = n1644 & n1271;
  assign n1257 = n1258 & ~n1276 & n1382;
  assign n1258 = ~n1281 & n1285;
  assign n1259 = n1276 & ~n1382;
  assign n1260 = n1256 & (n1257 | (n1258 & n1259));
  assign n1261 = n1268 | n1251 | ~n1259;
  assign n1262 = ~n1325 | ~n1382;
  assign n1263 = n1281 | n1268;
  assign n1264 = ~n1260 & n1261 & (n1262 | n1263);
  assign n1265 = ~n1271 | n1644;
  assign n1266 = ~n1276 | ~n1382;
  assign n1267 = ~n1258 | n1265 | n1266;
  assign n1268 = n1271 | ~n1644;
  assign n1269 = ~n1376 | n1268 | ~n1325;
  assign n1270 = ~n1256 | n1250 | n1251;
  assign n1271 = ~Pdata_44_ ^ ~PC_7_;
  assign n1272 = n1644 | ~n1315 | ~n1382;
  assign n1273 = ~n1281 | n1271 | n1272;
  assign n1274 = n1384 | n1268 | ~n1276;
  assign n1275 = n1952 & (n1265 | n1262 | n1281);
  assign n1276 = ~Pdata_39_ ^ ~PC_22_;
  assign n1277 = ~n1382 | n1263 | ~n1285;
  assign n1278 = n1274 & n1275 & (n1276 | n1277);
  assign n1279 = (~n1258 & n1276) | (n1251 & (~n1258 | ~n1276));
  assign n1280 = n1279 & (~n1281 | ~n1315);
  assign n1281 = ~Pdata_41_ ^ ~PC_11_;
  assign n1282 = ~n1376 & (n1281 | ~n1382);
  assign n1283 = ~n1317 | n1384;
  assign n1284 = n1283 & (~n1256 | n1282 | ~n1285);
  assign n1285 = ~Pdata_40_ ^ ~PC_18_;
  assign n1286 = (~n1258 | n1276) & (~n1281 | n1285);
  assign n1287 = (n1325 & ~n1644) | (~n1280 & (n1325 | n1644));
  assign n1288 = ~n1382 & ~n1271 & n1287;
  assign n1289 = n1272 | n1281;
  assign n1290 = (n746 | n1849) & (~Poutreg_31_ | n869);
  assign n1291 = (~Poutreg_30_ | n869) & (~Poutreg_22_ | Pcount_0_);
  assign n1292 = ~Pdata_59_ ^ ~PD_5_;
  assign n1293 = ~n1691 | n1292 | ~n1641;
  assign n1294 = ~n1690 | ~n1172 | ~n1173;
  assign n1295 = ~n1190 & ~n1641;
  assign n1296 = n1292 & ~n1300;
  assign n1297 = n1295 & (~n1170 | (n1173 & n1296));
  assign n1298 = n1299 & ~n1642;
  assign n1299 = ~Pdata_56_ ^ ~PD_20_;
  assign n1300 = ~Pdata_55_ ^ ~PD_15_;
  assign n1301 = ~n1190 & (n1298 | (n1299 & n1300));
  assign n1302 = n1299 & n1642;
  assign n1303 = n1190 & ~n1641;
  assign n1304 = n1302 & n1303;
  assign n1305 = (n746 | n1852) & (~Poutreg_29_ | n869);
  assign n1306 = (~Poutreg_28_ | n869) & (~Poutreg_20_ | Pcount_0_);
  assign n1307 = ~n1308 & (~n878 | ~n1397);
  assign n1308 = n887 & n888;
  assign n1309 = n1308 & n876;
  assign n1310 = ~n1398 & (~n1728 | (n896 & ~n1633));
  assign n1311 = ~n1633 | n1653;
  assign n1312 = n1311 | ~n1649;
  assign n1313 = (n746 | n1854) & (~Poutreg_27_ | n869);
  assign n1314 = (~Poutreg_26_ | n869) & (~Poutreg_18_ | Pcount_0_);
  assign n1315 = n1276 & ~n1285;
  assign n1316 = ~n1281 & ~n1382;
  assign n1317 = ~n1271 & ~n1644;
  assign n1318 = n1315 & n1316 & (n1317 | n1256);
  assign n1319 = n1697 | n1281 | ~n1325;
  assign n1320 = ~n1318 & n1319 & (~n1257 | ~n1317);
  assign n1321 = ~n1317 | n1251 | ~n1259;
  assign n1322 = ~n1315 | n1268 | n1282;
  assign n1323 = n1266 & n1250;
  assign n1324 = ~n1258 | n1323 | ~n1705;
  assign n1325 = ~n1276 & ~n1285;
  assign n1326 = ~n1382 & ~n1263 & n1325;
  assign n1327 = n1644 & ~n1276 & ~n1384;
  assign n1328 = n1327 & n1271;
  assign n1329 = (~Poutreg_25_ | n869) & (n746 | ~n1997);
  assign n1330 = (~Poutreg_24_ | n869) & (~Poutreg_16_ | Pcount_0_);
  assign n1331 = ~n914 | n1646;
  assign n1332 = ~n924 & n1331 & (n906 | ~n915);
  assign n1333 = ~n906 | n938;
  assign n1334 = (~n921 | n1332) & (~n1338 | ~n1658);
  assign n1335 = ~n1990 & n1333 & n939 & n905 & n910 & n1334;
  assign n1336 = (n746 | n1856) & (~Poutreg_23_ | n869);
  assign n1337 = (~Poutreg_22_ | n869) & (~Poutreg_14_ | Pcount_0_);
  assign n1338 = ~Pdata_33_ ^ ~PC_10_;
  assign n1339 = n921 & (n914 | n1338);
  assign n1340 = (n906 & ~n1729) | (n938 & (~n906 | ~n1729));
  assign n1341 = n939 & ~n1662;
  assign n1342 = n1961 | n1962 | n920 | ~n1338;
  assign n1343 = n903 & (~n914 | n1659);
  assign n1344 = ~n1963 & n1342 & n1341 & n910 & n1340 & n1343;
  assign n1345 = (n746 | n1857) & (~Poutreg_21_ | n869);
  assign n1346 = (~Poutreg_20_ | n869) & (~Poutreg_12_ | Pcount_0_);
  assign n1347 = ~n1061 | n1076 | ~n1222;
  assign n1348 = n1347 & (n1061 | ~n1076);
  assign n1349 = ~n1062 & n1087;
  assign n1350 = n1349 & ~n1061 & n1222;
  assign n1351 = ~n1076 & ~n1222;
  assign n1352 = n1076 & n1062 & n1222;
  assign n1353 = ~n1674 & (n1351 | n1352);
  assign n1354 = (n746 | n1860) & (~Poutreg_19_ | n869);
  assign n1355 = (~Poutreg_18_ | n869) & (~Poutreg_10_ | Pcount_0_);
  assign n1356 = n1302 & n1296 & n1303;
  assign n1357 = n1172 & ~n1174 & n1298;
  assign n1358 = n1641 & n1190;
  assign n1359 = (~n1642 & n1702) | (n1174 & (n1642 | n1702));
  assign n1360 = n1359 & ~n1299 & n1358;
  assign n1361 = n1298 & ~n1300 & ~n1641;
  assign n1362 = ~n1292 & (n1361 | ~n1370);
  assign n1363 = (~Poutreg_17_ | n869) & (n746 | ~n1998);
  assign n1364 = (~Poutreg_16_ | n869) & (~Poutreg_8_ | Pcount_0_);
  assign n1365 = n1702 | ~n1299 | ~n1694;
  assign n1366 = n1692 | n1299;
  assign n1367 = n1299 | n1179;
  assign n1368 = n1365 & n1366 & (~n1358 | n1367);
  assign n1369 = n1966 & (n1190 | ~n1300 | n1689);
  assign n1370 = ~n1299 | n1688;
  assign n1371 = ~n1361 & (~n1641 | (n1369 & n1370));
  assign n1372 = ~n1298 | n1179 | n1190;
  assign n1373 = n1303 & (~n1693 | ~n1695);
  assign n1374 = (n746 | n1863) & (~Poutreg_15_ | n869);
  assign n1375 = (~Poutreg_14_ | n869) & (~Poutreg_6_ | Pcount_0_);
  assign n1376 = n1281 & ~n1382;
  assign n1377 = ~n1285 & n1376;
  assign n1378 = n1263 | n1323;
  assign n1379 = (n746 | n1864) & (~Poutreg_13_ | n869);
  assign n1380 = (~Poutreg_12_ | n869) & (~Poutreg_4_ | Pcount_0_);
  assign n1381 = n1317 | ~n1382;
  assign n1382 = ~Pdata_43_ ^ ~PC_25_;
  assign n1383 = ~n1285 & n1381 & (~n1263 | n1382);
  assign n1384 = n1251 | ~n1382;
  assign n1385 = n1277 & ~n1383 & (~n1271 | n1384);
  assign n1386 = n1698 & n1321 & n1278 & n1320;
  assign n1387 = (n1276 & n1385) | (n1283 & (~n1276 | n1385));
  assign n1388 = n1705 | n1262 | ~n1281;
  assign n1389 = ~n1644 | n1250 | ~n1258;
  assign n1390 = (n1280 | n1697) & (n1382 | n1706);
  assign n1391 = n1390 & n1388 & n1387 & n1386 & n1264 & n1389;
  assign n1392 = (n746 | n1865) & (~Poutreg_11_ | n869);
  assign n1393 = (~Poutreg_10_ | n869) & (~Poutreg_2_ | Pcount_0_);
  assign n1394 = ~n872 & n1397;
  assign n1395 = n887 & ~n1634;
  assign n1396 = n897 & n1394 & (n1395 | n878);
  assign n1397 = ~Pdata_47_ ^ ~PD_12_;
  assign n1398 = ~Pdata_52_ ^ ~PD_26_;
  assign n1399 = ~n1972 | n1397 | n1398;
  assign n1400 = n881 | ~n894;
  assign n1401 = (n746 | n1866) & (~Poutreg_9_ | n869);
  assign n1402 = (~Poutreg_8_ | n869) & (~Poutreg_0_ | Pcount_0_);
  assign n1403 = Pcount_0_ | n1404;
  assign n1404 = n837 | Preset_0_;
  assign n1405 = n1403 & (Pcount_1_ | n1404);
  assign n1406 = n1405 & (Pcount_2_ | n1404);
  assign n1407 = Pcount_3_ | n1648;
  assign n1408 = n746 & n1407 & (Pcount_0_ | ~n1798);
  assign n1409 = (~PC_26_ | n1712) & (~PC_0_ | n1713);
  assign n1410 = (~PC_25_ | n1709) & (~PC_1_ | n1711);
  assign n1411 = (~PC_27_ | n1718) & n1867;
  assign n1412 = n1411 & n1409 & n1410;
  assign n1413 = (~PC_27_ | n1713) & (~PC_25_ | n1712);
  assign n1414 = (~PC_24_ | n1709) & (~PC_0_ | n1711);
  assign n1415 = (~PC_26_ | n1718) & n1868;
  assign n1416 = n1415 & n1413 & n1414;
  assign n1417 = (~PC_26_ | n1713) & (~PC_24_ | n1712);
  assign n1418 = (~PC_27_ | n1711) & (~PC_23_ | n1709);
  assign n1419 = (~PC_25_ | n1718) & n1869;
  assign n1420 = n1419 & n1417 & n1418;
  assign n1421 = (~PC_25_ | n1713) & (~PC_23_ | n1712);
  assign n1422 = (~PC_26_ | n1711) & (~PC_22_ | n1709);
  assign n1423 = (~PC_24_ | n1718) & n1870;
  assign n1424 = n1423 & n1421 & n1422;
  assign n1425 = (~PC_24_ | n1713) & (~PC_22_ | n1712);
  assign n1426 = (~PC_25_ | n1711) & (~PC_21_ | n1709);
  assign n1427 = (~PC_23_ | n1718) & n1871;
  assign n1428 = n1427 & n1425 & n1426;
  assign n1429 = (~PC_23_ | n1713) & (~PC_21_ | n1712);
  assign n1430 = (~PC_24_ | n1711) & (~PC_20_ | n1709);
  assign n1431 = (~PC_22_ | n1718) & n1872;
  assign n1432 = n1431 & n1429 & n1430;
  assign n1433 = (~PC_22_ | n1713) & (~PC_20_ | n1712);
  assign n1434 = (~PC_23_ | n1711) & (~PC_19_ | n1709);
  assign n1435 = (~PC_21_ | n1718) & n1873;
  assign n1436 = n1435 & n1433 & n1434;
  assign n1437 = (~PC_21_ | n1713) & (~PC_19_ | n1712);
  assign n1438 = (~PC_22_ | n1711) & (~PC_18_ | n1709);
  assign n1439 = (~PC_20_ | n1718) & n1874;
  assign n1440 = n1439 & n1437 & n1438;
  assign n1441 = (~PC_20_ | n1713) & (~PC_18_ | n1712);
  assign n1442 = (~PC_21_ | n1711) & (~PC_17_ | n1709);
  assign n1443 = (~PC_19_ | n1718) & n1875;
  assign n1444 = n1443 & n1441 & n1442;
  assign n1445 = (~PC_19_ | n1713) & (~PC_17_ | n1712);
  assign n1446 = (~PC_20_ | n1711) & (~PC_16_ | n1709);
  assign n1447 = (~PC_18_ | n1718) & n1876;
  assign n1448 = n1447 & n1445 & n1446;
  assign n1449 = (~PC_18_ | n1713) & (~PC_16_ | n1712);
  assign n1450 = (~PC_19_ | n1711) & (~PC_15_ | n1709);
  assign n1451 = (~PC_17_ | n1718) & n1877;
  assign n1452 = n1451 & n1449 & n1450;
  assign n1453 = (~PC_17_ | n1713) & (~PC_15_ | n1712);
  assign n1454 = (~PC_18_ | n1711) & (~PC_14_ | n1709);
  assign n1455 = (~PC_16_ | n1718) & n1878;
  assign n1456 = n1455 & n1453 & n1454;
  assign n1457 = (~PC_16_ | n1713) & (~PC_14_ | n1712);
  assign n1458 = (~PC_17_ | n1711) & (~PC_13_ | n1709);
  assign n1459 = (~PC_15_ | n1718) & n1879;
  assign n1460 = n1459 & n1457 & n1458;
  assign n1461 = (~PC_15_ | n1713) & (~PC_13_ | n1712);
  assign n1462 = (~PC_16_ | n1711) & (~PC_12_ | n1709);
  assign n1463 = (~PC_14_ | n1718) & n1880;
  assign n1464 = n1463 & n1461 & n1462;
  assign n1465 = (~PC_14_ | n1713) & (~PC_12_ | n1712);
  assign n1466 = (~PC_15_ | n1711) & (~PC_11_ | n1709);
  assign n1467 = (~PC_13_ | n1718) & n1881;
  assign n1468 = n1467 & n1465 & n1466;
  assign n1469 = (~PC_13_ | n1713) & (~PC_11_ | n1712);
  assign n1470 = (~PC_14_ | n1711) & (~PC_10_ | n1709);
  assign n1471 = (~PC_12_ | n1718) & n1882;
  assign n1472 = n1471 & n1469 & n1470;
  assign n1473 = (~PC_12_ | n1713) & (~PC_10_ | n1712);
  assign n1474 = (~PC_13_ | n1711) & (~PC_9_ | n1709);
  assign n1475 = (~PC_11_ | n1718) & n1883;
  assign n1476 = n1475 & n1473 & n1474;
  assign n1477 = (~PC_11_ | n1713) & (~PC_9_ | n1712);
  assign n1478 = (~PC_12_ | n1711) & (~PC_8_ | n1709);
  assign n1479 = (~PC_10_ | n1718) & n1884;
  assign n1480 = n1479 & n1477 & n1478;
  assign n1481 = (~PC_10_ | n1713) & (~PC_8_ | n1712);
  assign n1482 = (~PC_11_ | n1711) & (~PC_7_ | n1709);
  assign n1483 = (~PC_9_ | n1718) & n1885;
  assign n1484 = n1483 & n1481 & n1482;
  assign n1485 = (~PC_9_ | n1713) & (~PC_7_ | n1712);
  assign n1486 = (~PC_10_ | n1711) & (~PC_6_ | n1709);
  assign n1487 = (~PC_8_ | n1718) & n1886;
  assign n1488 = n1487 & n1485 & n1486;
  assign n1489 = (~PC_8_ | n1713) & (~PC_6_ | n1712);
  assign n1490 = (~PC_9_ | n1711) & (~PC_5_ | n1709);
  assign n1491 = (~PC_7_ | n1718) & n1887;
  assign n1492 = n1491 & n1489 & n1490;
  assign n1493 = (~PC_7_ | n1713) & (~PC_5_ | n1712);
  assign n1494 = (~PC_8_ | n1711) & (~PC_4_ | n1709);
  assign n1495 = (~PC_6_ | n1718) & n1888;
  assign n1496 = n1495 & n1493 & n1494;
  assign n1497 = (~PC_6_ | n1713) & (~PC_4_ | n1712);
  assign n1498 = (~PC_7_ | n1711) & (~PC_3_ | n1709);
  assign n1499 = (~PC_5_ | n1718) & n1889;
  assign n1500 = n1499 & n1497 & n1498;
  assign n1501 = (~PC_5_ | n1713) & (~PC_3_ | n1712);
  assign n1502 = (~PC_6_ | n1711) & (~PC_2_ | n1709);
  assign n1503 = (~PC_4_ | n1718) & n1890;
  assign n1504 = n1503 & n1501 & n1502;
  assign n1505 = (~PC_4_ | n1713) & (~PC_2_ | n1712);
  assign n1506 = (~PC_5_ | n1711) & (~PC_1_ | n1709);
  assign n1507 = (~PC_3_ | n1718) & n1891;
  assign n1508 = n1507 & n1505 & n1506;
  assign n1509 = (~PC_3_ | n1713) & (~PC_1_ | n1712);
  assign n1510 = (~PC_4_ | n1711) & (~PC_0_ | n1709);
  assign n1511 = (~PC_2_ | n1718) & n1892;
  assign n1512 = n1511 & n1509 & n1510;
  assign n1513 = (~PC_2_ | n1713) & (~PC_0_ | n1712);
  assign n1514 = (~PC_27_ | n1709) & (~PC_3_ | n1711);
  assign n1515 = (~PC_1_ | n1718) & n1893;
  assign n1516 = n1515 & n1513 & n1514;
  assign n1517 = (~PC_27_ | n1712) & (~PC_1_ | n1713);
  assign n1518 = (~PC_26_ | n1709) & (~PC_2_ | n1711);
  assign n1519 = (~PC_0_ | n1718) & n1894;
  assign n1520 = n1519 & n1517 & n1518;
  assign n1521 = (~PD_26_ | n1712) & (~PD_0_ | n1713);
  assign n1522 = (~PD_25_ | n1709) & (~PD_1_ | n1711);
  assign n1523 = (~PD_27_ | n1718) & n1895;
  assign n1524 = n1523 & n1521 & n1522;
  assign n1525 = (~PD_27_ | n1713) & (~PD_25_ | n1712);
  assign n1526 = (~PD_24_ | n1709) & (~PD_0_ | n1711);
  assign n1527 = (~PD_26_ | n1718) & n1896;
  assign n1528 = n1527 & n1525 & n1526;
  assign n1529 = (~PD_26_ | n1713) & (~PD_24_ | n1712);
  assign n1530 = (~PD_27_ | n1711) & (~PD_23_ | n1709);
  assign n1531 = (~PD_25_ | n1718) & n1897;
  assign n1532 = n1531 & n1529 & n1530;
  assign n1533 = (~PD_25_ | n1713) & (~PD_23_ | n1712);
  assign n1534 = (~PD_26_ | n1711) & (~PD_22_ | n1709);
  assign n1535 = (~PD_24_ | n1718) & n1898;
  assign n1536 = n1535 & n1533 & n1534;
  assign n1537 = (~PD_24_ | n1713) & (~PD_22_ | n1712);
  assign n1538 = (~PD_25_ | n1711) & (~PD_21_ | n1709);
  assign n1539 = (~PD_23_ | n1718) & n1899;
  assign n1540 = n1539 & n1537 & n1538;
  assign n1541 = (~PD_23_ | n1713) & (~PD_21_ | n1712);
  assign n1542 = (~PD_24_ | n1711) & (~PD_20_ | n1709);
  assign n1543 = (~PD_22_ | n1718) & n1900;
  assign n1544 = n1543 & n1541 & n1542;
  assign n1545 = (~PD_22_ | n1713) & (~PD_20_ | n1712);
  assign n1546 = (~PD_23_ | n1711) & (~PD_19_ | n1709);
  assign n1547 = (~PD_21_ | n1718) & n1901;
  assign n1548 = n1547 & n1545 & n1546;
  assign n1549 = (~PD_21_ | n1713) & (~PD_19_ | n1712);
  assign n1550 = (~PD_22_ | n1711) & (~PD_18_ | n1709);
  assign n1551 = (~PD_20_ | n1718) & n1902;
  assign n1552 = n1551 & n1549 & n1550;
  assign n1553 = (~PD_20_ | n1713) & (~PD_18_ | n1712);
  assign n1554 = (~PD_21_ | n1711) & (~PD_17_ | n1709);
  assign n1555 = (~PD_19_ | n1718) & n1903;
  assign n1556 = n1555 & n1553 & n1554;
  assign n1557 = (~PD_19_ | n1713) & (~PD_17_ | n1712);
  assign n1558 = (~PD_20_ | n1711) & (~PD_16_ | n1709);
  assign n1559 = (~PD_18_ | n1718) & n1904;
  assign n1560 = n1559 & n1557 & n1558;
  assign n1561 = (~PD_18_ | n1713) & (~PD_16_ | n1712);
  assign n1562 = (~PD_19_ | n1711) & (~PD_15_ | n1709);
  assign n1563 = (~PD_17_ | n1718) & n1905;
  assign n1564 = n1563 & n1561 & n1562;
  assign n1565 = (~PD_17_ | n1713) & (~PD_15_ | n1712);
  assign n1566 = (~PD_18_ | n1711) & (~PD_14_ | n1709);
  assign n1567 = (~PD_16_ | n1718) & n1906;
  assign n1568 = n1567 & n1565 & n1566;
  assign n1569 = (~PD_16_ | n1713) & (~PD_14_ | n1712);
  assign n1570 = (~PD_17_ | n1711) & (~PD_13_ | n1709);
  assign n1571 = (~PD_15_ | n1718) & n1907;
  assign n1572 = n1571 & n1569 & n1570;
  assign n1573 = (~PD_15_ | n1713) & (~PD_13_ | n1712);
  assign n1574 = (~PD_16_ | n1711) & (~PD_12_ | n1709);
  assign n1575 = (~PD_14_ | n1718) & n1908;
  assign n1576 = n1575 & n1573 & n1574;
  assign n1577 = (~PD_14_ | n1713) & (~PD_12_ | n1712);
  assign n1578 = (~PD_15_ | n1711) & (~PD_11_ | n1709);
  assign n1579 = (~PD_13_ | n1718) & n1909;
  assign n1580 = n1579 & n1577 & n1578;
  assign n1581 = (~PD_13_ | n1713) & (~PD_11_ | n1712);
  assign n1582 = (~PD_14_ | n1711) & (~PD_10_ | n1709);
  assign n1583 = (~PD_12_ | n1718) & n1910;
  assign n1584 = n1583 & n1581 & n1582;
  assign n1585 = (~PD_12_ | n1713) & (~PD_10_ | n1712);
  assign n1586 = (~PD_13_ | n1711) & (~PD_9_ | n1709);
  assign n1587 = (~PD_11_ | n1718) & n1911;
  assign n1588 = n1587 & n1585 & n1586;
  assign n1589 = (~PD_11_ | n1713) & (~PD_9_ | n1712);
  assign n1590 = (~PD_12_ | n1711) & (~PD_8_ | n1709);
  assign n1591 = (~PD_10_ | n1718) & n1912;
  assign n1592 = n1591 & n1589 & n1590;
  assign n1593 = (~PD_10_ | n1713) & (~PD_8_ | n1712);
  assign n1594 = (~PD_11_ | n1711) & (~PD_7_ | n1709);
  assign n1595 = (~PD_9_ | n1718) & n1913;
  assign n1596 = n1595 & n1593 & n1594;
  assign n1597 = (~PD_9_ | n1713) & (~PD_7_ | n1712);
  assign n1598 = (~PD_10_ | n1711) & (~PD_6_ | n1709);
  assign n1599 = (~PD_8_ | n1718) & n1914;
  assign n1600 = n1599 & n1597 & n1598;
  assign n1601 = (~PD_8_ | n1713) & (~PD_6_ | n1712);
  assign n1602 = (~PD_9_ | n1711) & (~PD_5_ | n1709);
  assign n1603 = (~PD_7_ | n1718) & n1915;
  assign n1604 = n1603 & n1601 & n1602;
  assign n1605 = (~PD_7_ | n1713) & (~PD_5_ | n1712);
  assign n1606 = (~PD_8_ | n1711) & (~PD_4_ | n1709);
  assign n1607 = (~PD_6_ | n1718) & n1916;
  assign n1608 = n1607 & n1605 & n1606;
  assign n1609 = (~PD_6_ | n1713) & (~PD_4_ | n1712);
  assign n1610 = (~PD_7_ | n1711) & (~PD_3_ | n1709);
  assign n1611 = (~PD_5_ | n1718) & n1917;
  assign n1612 = n1611 & n1609 & n1610;
  assign n1613 = (~PD_5_ | n1713) & (~PD_3_ | n1712);
  assign n1614 = (~PD_6_ | n1711) & (~PD_2_ | n1709);
  assign n1615 = (~PD_4_ | n1718) & n1918;
  assign n1616 = n1615 & n1613 & n1614;
  assign n1617 = (~PD_4_ | n1713) & (~PD_2_ | n1712);
  assign n1618 = (~PD_5_ | n1711) & (~PD_1_ | n1709);
  assign n1619 = (~PD_3_ | n1718) & n1919;
  assign n1620 = n1619 & n1617 & n1618;
  assign n1621 = (~PD_3_ | n1713) & (~PD_1_ | n1712);
  assign n1622 = (~PD_4_ | n1711) & (~PD_0_ | n1709);
  assign n1623 = (~PD_2_ | n1718) & n1920;
  assign n1624 = n1623 & n1621 & n1622;
  assign n1625 = (~PD_2_ | n1713) & (~PD_0_ | n1712);
  assign n1626 = (~PD_27_ | n1709) & (~PD_3_ | n1711);
  assign n1627 = (~PD_1_ | n1718) & n1921;
  assign n1628 = n1627 & n1625 & n1626;
  assign n1629 = (~PD_27_ | n1712) & (~PD_1_ | n1713);
  assign n1630 = (~PD_26_ | n1709) & (~PD_2_ | n1711);
  assign n1631 = (~PD_0_ | n1718) & n1922;
  assign n1632 = n1631 & n1629 & n1630;
  assign n1633 = ~Pdata_48_ ^ ~PD_23_;
  assign n1634 = ~Pdata_51_ ^ ~PD_18_;
  assign n1635 = ~Pdata_45_ ^ ~PC_26_;
  assign n1636 = ~Pdata_38_ ^ ~PC_5_;
  assign n1637 = n993 & (~n1002 | (n1039 & ~n1149));
  assign n1638 = ~Pdata_52_ ^ ~PD_11_;
  assign n1639 = ~Pdata_56_ ^ ~PD_19_;
  assign n1640 = ~n1639 ^ ~n1133;
  assign n1641 = ~Pdata_60_ ^ ~PD_24_;
  assign n1642 = ~Pdata_58_ ^ ~PD_27_;
  assign n1643 = ~n1062 ^ n1076;
  assign n1644 = ~Pdata_42_ ^ ~PC_3_;
  assign n1645 = ~n1649 & (~n887 | ~n1633);
  assign n1646 = ~n906 ^ n1338;
  assign n1647 = ~Pencrypt_mode_0_ ^ Pencrypt_0_;
  assign n1648 = ~Pcount_0_ | ~Pcount_2_ | ~Pcount_1_;
  assign n1649 = ~n887 & ~n1634;
  assign n1650 = n887 & n1634;
  assign n1651 = ~n1398 & ~n1633;
  assign n1652 = n1649 & n876;
  assign n1653 = n1398 | ~n872 | ~n1397;
  assign n1654 = ~n1397 | ~n872 | ~n876;
  assign n1655 = ~n1338 | n916 | ~n920;
  assign n1656 = n920 & n901;
  assign n1657 = n914 & ~n1338;
  assign n1658 = ~n920 & ~n914 & n916;
  assign n1659 = ~n1338 | n920 | ~n921;
  assign n1660 = n1656 & ~n906 & n914;
  assign n1661 = n906 & n1657 & n935;
  assign n1662 = n1660 | n1661 | n925 | n927;
  assign n1663 = n980 | n972;
  assign n1664 = n972 | ~n980;
  assign n1665 = ~n980 | n1635;
  assign n1666 = n956 | n1030 | n980;
  assign n1667 = n1665 | n956 | n981;
  assign n1668 = n1664 | n956 | n958;
  assign n1669 = n956 | ~n980 | n1030 | ~n1635;
  assign n1670 = n993 | n1146;
  assign n1671 = n989 | n993;
  assign n1672 = n1076 & ~n1222;
  assign n1673 = ~n1061 | n1071;
  assign n1674 = ~n1061 | n1087;
  assign n1675 = ~n1062 & ~n1674;
  assign n1676 = n1078 | n1347;
  assign n1677 = n1061 & n1087;
  assign n1678 = ~n1088 & n1085 & n1086;
  assign n1679 = n1078 | n1071 | ~n1076;
  assign n1680 = ~n1078 | n1087 | n1347;
  assign n1681 = ~n1102 & ~n1120;
  assign n1682 = n1120 & n1133;
  assign n1683 = n1102 & n1682;
  assign n1684 = ~n1102 | n1119;
  assign n1685 = ~n1133 | ~n1681;
  assign n1686 = ~n1104 | n1133;
  assign n1687 = n989 | ~n996;
  assign n1688 = ~n1642 | n1190 | n1300;
  assign n1689 = n1299 | ~n1642;
  assign n1690 = n1300 & n1292;
  assign n1691 = ~n1299 & ~n1688;
  assign n1692 = ~n1174 | ~n1303;
  assign n1693 = n1179 | ~n1302;
  assign n1694 = ~n1172 & ~n1303;
  assign n1695 = n1367 | n1642;
  assign n1696 = n1639 & n1133;
  assign n1697 = n1382 | n1265;
  assign n1698 = n1269 & n1267 & n1270 & n1273;
  assign n1699 = n1255 & n1698 & n1264;
  assign n1700 = n1303 & ~n1642 & n1690;
  assign n1701 = n1190 | n1695;
  assign n1702 = ~n1174 & ~n1690;
  assign n1703 = ~n1297 & n1294 & n1187 & n1293;
  assign n1704 = n886 & n1139;
  assign n1705 = n1317 | n1256;
  assign n1706 = ~n1705 | ~n1281 | ~n1325;
  assign n1707 = n1404 | ~n1717;
  assign n1708 = Pencrypt_mode_0_ | n1707;
  assign n1709 = ~n1408 | n1708;
  assign n1710 = ~Pencrypt_mode_0_ | n1707;
  assign n1711 = ~n1408 | n1710;
  assign n1712 = n1408 | n1708;
  assign n1713 = n1408 | n1710;
  assign n1714 = Preset_0_ | ~n837;
  assign n1715 = Pencrypt_0_ | n1714;
  assign n1716 = ~Pencrypt_0_ | n1714;
  assign n1717 = n1647 | n746;
  assign n1718 = n1404 | n1717;
  assign n1719 = n1923 & (~n900 | n913 | ~n916);
  assign n1720 = ~n1925 & (~n906 | (n914 & n935));
  assign n1721 = (n934 & ~n1338) | (n926 & (n934 | n1338));
  assign n1722 = n956 & (n961 | (~n958 & n981));
  assign n1723 = (~n980 & ~n1722) | (n975 & (n980 | ~n1722));
  assign n1724 = (~n954 & (~n956 | ~n1664)) | (n956 & ~n1664);
  assign n1725 = ~n1936 & (n887 | ~n892 | n1397);
  assign n1726 = (n1641 & n1691) | (~n1370 & (~n1641 | n1691));
  assign n1727 = n1943 & (n1199 | ~n1201);
  assign n1728 = (n1397 & n1645) | (~n878 & (~n1397 | n1645));
  assign n1729 = n920 & (n1339 | (n1657 & n912));
  assign n1730 = n892 & (n896 | (~n887 & n888));
  assign n1731 = n1650 & (n892 | (~n1397 & n1398));
  assign n1732 = (n746 & n1863) | (~Pdata_in_6_ & (~n746 | n1863));
  assign n1733 = (n746 & n1856) | (~Pinreg_6_ & (~n746 | n1856));
  assign n1734 = (n746 & n1849) | (~Pinreg_14_ & (~n746 | n1849));
  assign n1735 = (n746 & n1843) | (~Pinreg_22_ & (~n746 | n1843));
  assign n1736 = (n746 & n1836) | (~Pinreg_30_ & (~n746 | n1836));
  assign n1737 = (n746 & n1820) | (~Pinreg_38_ & (~n746 | n1820));
  assign n1738 = (n746 & n1810) | (~Pinreg_46_ & (~n746 | n1810));
  assign n1739 = (n746 & n899) | (~Pinreg_54_ & (~n746 | n899));
  assign n1740 = (n746 & n1864) | (~Pdata_in_4_ & (~n746 | n1864));
  assign n1741 = (n746 & n1857) | (~Pinreg_4_ & (~n746 | n1857));
  assign n1742 = (n746 & n1852) | (~Pinreg_12_ & (~n746 | n1852));
  assign n1743 = (n746 & n1844) | (~Pinreg_20_ & (~n746 | n1844));
  assign n1744 = (n746 & n1837) | (~Pinreg_28_ & (~n746 | n1837));
  assign n1745 = (n746 & n1829) | (~Pinreg_36_ & (~n746 | n1829));
  assign n1746 = (n746 & n1815) | (~Pinreg_44_ & (~n746 | n1815));
  assign n1747 = (n746 & n931) | (~Pinreg_52_ & (~n746 | n931));
  assign n1748 = (n746 & n1865) | (~Pdata_in_2_ & (~n746 | n1865));
  assign n1749 = (n746 & n1860) | (~Pinreg_2_ & (~n746 | n1860));
  assign n1750 = (n746 & n1854) | (~Pinreg_10_ & (~n746 | n1854));
  assign n1751 = (n746 & n1845) | (~Pinreg_18_ & (~n746 | n1845));
  assign n1752 = (n746 & n1838) | (~Pinreg_26_ & (~n746 | n1838));
  assign n1753 = (n746 & n1834) | (~Pinreg_34_ & (~n746 | n1834));
  assign n1754 = (n746 & n1816) | (~Pinreg_42_ & (~n746 | n1816));
  assign n1755 = (n746 & n948) | (~Pinreg_50_ & (~n746 | n948));
  assign n1756 = (n746 & n1866) | (~Pdata_in_0_ & (~n746 | n1866));
  assign n1757 = (~Pinreg_0_ & (~n746 | ~n1998)) | (n746 & ~n1998);
  assign n1758 = (~Pinreg_8_ & (~n746 | ~n1997)) | (n746 & ~n1997);
  assign n1759 = (n746 & n1847) | (~Pinreg_16_ & (~n746 | n1847));
  assign n1760 = (n746 & n1840) | (~Pinreg_24_ & (~n746 | n1840));
  assign n1761 = (~Pinreg_32_ & (~n746 | ~n1996)) | (n746 & ~n1996);
  assign n1762 = (n746 & n1817) | (~Pinreg_40_ & (~n746 | n1817));
  assign n1763 = (n746 & n976) | (~Pinreg_48_ & (~n746 | n976));
  assign n1764 = (~Pdata_63_ & n746) | (~Pdata_in_7_ & (~Pdata_63_ | ~n746));
  assign n1765 = (~Pdata_62_ & n746) | (~Pinreg_7_ & (~Pdata_62_ | ~n746));
  assign n1766 = (~Pdata_61_ & n746) | (~Pinreg_15_ & (~Pdata_61_ | ~n746));
  assign n1767 = (~Pdata_60_ & n746) | (~Pinreg_23_ & (~Pdata_60_ | ~n746));
  assign n1768 = (~Pdata_59_ & n746) | (~Pinreg_31_ & (~Pdata_59_ | ~n746));
  assign n1769 = (~Pdata_58_ & n746) | (~Pinreg_39_ & (~Pdata_58_ | ~n746));
  assign n1770 = (~Pdata_57_ & n746) | (~Pinreg_47_ & (~Pdata_57_ | ~n746));
  assign n1771 = (~Pdata_56_ & n746) | (~Pinreg_55_ & (~Pdata_56_ | ~n746));
  assign n1772 = (~Pdata_55_ & n746) | (~Pdata_in_5_ & (~Pdata_55_ | ~n746));
  assign n1773 = (~Pdata_54_ & n746) | (~Pinreg_5_ & (~Pdata_54_ | ~n746));
  assign n1774 = (~Pdata_53_ & n746) | (~Pinreg_13_ & (~Pdata_53_ | ~n746));
  assign n1775 = (~Pdata_52_ & n746) | (~Pinreg_21_ & (~Pdata_52_ | ~n746));
  assign n1776 = (~Pdata_51_ & n746) | (~Pinreg_29_ & (~Pdata_51_ | ~n746));
  assign n1777 = (~Pdata_50_ & n746) | (~Pinreg_37_ & (~Pdata_50_ | ~n746));
  assign n1778 = (~Pdata_49_ & n746) | (~Pinreg_45_ & (~Pdata_49_ | ~n746));
  assign n1779 = (~Pdata_48_ & n746) | (~Pinreg_53_ & (~Pdata_48_ | ~n746));
  assign n1780 = (~Pdata_47_ & n746) | (~Pdata_in_3_ & (~Pdata_47_ | ~n746));
  assign n1781 = (~Pdata_46_ & n746) | (~Pinreg_3_ & (~Pdata_46_ | ~n746));
  assign n1782 = (~Pdata_45_ & n746) | (~Pinreg_11_ & (~Pdata_45_ | ~n746));
  assign n1783 = (~Pdata_44_ & n746) | (~Pinreg_19_ & (~Pdata_44_ | ~n746));
  assign n1784 = (~Pdata_43_ & n746) | (~Pinreg_27_ & (~Pdata_43_ | ~n746));
  assign n1785 = (~Pdata_42_ & n746) | (~Pinreg_35_ & (~Pdata_42_ | ~n746));
  assign n1786 = (~Pdata_41_ & n746) | (~Pinreg_43_ & (~Pdata_41_ | ~n746));
  assign n1787 = (~Pdata_40_ & n746) | (~Pinreg_51_ & (~Pdata_40_ | ~n746));
  assign n1788 = (~Pdata_39_ & n746) | (~Pdata_in_1_ & (~Pdata_39_ | ~n746));
  assign n1789 = (~Pdata_38_ & n746) | (~Pinreg_1_ & (~Pdata_38_ | ~n746));
  assign n1790 = (~Pdata_37_ & n746) | (~Pinreg_9_ & (~Pdata_37_ | ~n746));
  assign n1791 = (~Pdata_36_ & n746) | (~Pinreg_17_ & (~Pdata_36_ | ~n746));
  assign n1792 = (~Pdata_35_ & n746) | (~Pinreg_25_ & (~Pdata_35_ | ~n746));
  assign n1793 = (~Pdata_34_ & n746) | (~Pinreg_33_ & (~Pdata_34_ | ~n746));
  assign n1794 = (~Pdata_33_ & n746) | (~Pinreg_41_ & (~Pdata_33_ | ~n746));
  assign n1795 = (~Pdata_32_ & n746) | (~Pinreg_49_ & (~Pdata_32_ | ~n746));
  assign n1796 = (~Pcount_2_ | n1405) & n1974;
  assign n1797 = (~Pcount_1_ | n1403) & n1975;
  assign n1798 = ~n1976 & (~Pcount_1_ | (Pcount_3_ & Pcount_2_));
  assign n1799 = (~Pencrypt_0_ & ~n746) | (~Pencrypt_mode_0_ & (~Pencrypt_0_ | n746));
  assign n1800 = n872 | ~n876 | ~n878 | n1397;
  assign n1801 = (~n1395 | n1654) & (n887 | n1311);
  assign n1802 = (~n1142 | ~n1397) & (~n1649 | n1653);
  assign n1803 = ~n916 | n1338 | n913 | n914;
  assign n1804 = ~n1163 | n980 | ~n1161;
  assign n1805 = n1665 | ~n981 | ~n1161;
  assign n1806 = (n973 | n980) & (n1159 | n1668);
  assign n1807 = n968 | n1635 | n981;
  assign n1808 = n1807 & (~n958 | n980 | n1030);
  assign n1809 = ~n1163 | ~n980 | ~n1161;
  assign n1810 = ~Pdata_25_ ^ ~n1980;
  assign n1811 = ~n1051 | n1005 | ~n1039;
  assign n1812 = ~n1051 | ~n1039 | ~n1049;
  assign n1813 = n1812 & (n1013 | n993 | n1056);
  assign n1814 = n1146 | n989 | ~n1050;
  assign n1815 = ~n1023 ^ ~Pdata_17_;
  assign n1816 = ~n1036 ^ ~Pdata_9_;
  assign n1817 = ~Pdata_1_ ^ ~n1981;
  assign n1818 = ~n1076 | n1077;
  assign n1819 = ~n1061 | n1679;
  assign n1820 = ~n1098 ^ ~Pdata_26_;
  assign n1821 = n1207 | n1117 | ~n1201;
  assign n1822 = n1101 | ~n1133;
  assign n1823 = n1116 | n1112;
  assign n1824 = ~n1201 | n1129 | ~n1132;
  assign n1825 = (~n1638 | n1685) & (n1112 | n1211);
  assign n1826 = (n1121 | ~n1132) & (~n1681 | n1686);
  assign n1827 = ~n1640 | n1200 | n1638;
  assign n1828 = n1827 & (n1109 | (~n1105 & n1117));
  assign n1829 = ~n1125 ^ ~Pdata_18_;
  assign n1830 = n1686 | n1200 | n1201;
  assign n1831 = n1207 | n1121 | n1102;
  assign n1832 = n1831 & (n1103 | n1686);
  assign n1833 = (n1211 | ~n1683) & (n1205 | n1638);
  assign n1834 = ~Pdata_10_ ^ ~n1982;
  assign n1835 = (~n1039 | n1053) & (n1005 | n1042);
  assign n1836 = ~n1156 ^ ~Pdata_27_;
  assign n1837 = ~Pdata_19_ ^ ~n1984;
  assign n1838 = ~n1196 ^ ~Pdata_11_;
  assign n1839 = (n1202 | n1686) & (n1116 | ~n1683);
  assign n1840 = ~Pdata_3_ ^ ~n1985;
  assign n1841 = n1682 | ~n1102 | ~n1132;
  assign n1842 = ~n1133 | n1102 | ~n1104;
  assign n1843 = ~n1215 ^ ~Pdata_28_;
  assign n1844 = ~n1232 ^ ~Pdata_20_;
  assign n1845 = ~n1241 ^ ~Pdata_12_;
  assign n1846 = (n1076 & n1673) | (n1075 & (~n1076 | n1673));
  assign n1847 = ~n1247 ^ ~Pdata_4_;
  assign n1848 = (~n1276 | n1284) & (n1286 | n1697);
  assign n1849 = ~Pdata_29_ ^ ~n1986;
  assign n1850 = n1694 | ~n1296 | ~n1298;
  assign n1851 = n1850 & (n1299 | ~n1700);
  assign n1852 = ~Pdata_21_ ^ ~n1987;
  assign n1853 = (~n892 | n1307) & (n1397 | ~n1652);
  assign n1854 = ~Pdata_13_ ^ ~n1988;
  assign n1855 = (n1271 | n1262) & (n1265 | n1266);
  assign n1856 = ~n1335 ^ ~Pdata_30_;
  assign n1857 = ~n1344 ^ ~Pdata_22_;
  assign n1858 = n1673 & (~n1062 | ~n1087 | n1348);
  assign n1859 = (n1071 | n1076) & (n1089 | ~n1222);
  assign n1860 = ~Pdata_14_ ^ ~n1991;
  assign n1861 = (n1641 | n1701) & (~n1190 | n1693);
  assign n1862 = (~n1292 | n1371) & (n1368 | ~n1642);
  assign n1863 = ~Pdata_31_ ^ ~n1993;
  assign n1864 = ~Pdata_23_ ^ ~n1994;
  assign n1865 = ~n1391 ^ ~Pdata_15_;
  assign n1866 = ~Pdata_7_ ^ ~n1995;
  assign n1867 = (~Pinreg_48_ | n1716) & (~Pinreg_27_ | n1715);
  assign n1868 = (~Pinreg_35_ | n1715) & (~Pinreg_27_ | n1716);
  assign n1869 = (~Pinreg_43_ | n1715) & (~Pinreg_35_ | n1716);
  assign n1870 = (~Pinreg_51_ | n1715) & (~Pinreg_43_ | n1716);
  assign n1871 = (~Pinreg_51_ | n1716) & (~Pdata_in_2_ | n1715);
  assign n1872 = (~Pinreg_2_ | n1715) & (~Pdata_in_2_ | n1716);
  assign n1873 = (~Pinreg_10_ | n1715) & (~Pinreg_2_ | n1716);
  assign n1874 = (~Pinreg_18_ | n1715) & (~Pinreg_10_ | n1716);
  assign n1875 = (~Pinreg_26_ | n1715) & (~Pinreg_18_ | n1716);
  assign n1876 = (~Pinreg_34_ | n1715) & (~Pinreg_26_ | n1716);
  assign n1877 = (~Pinreg_42_ | n1715) & (~Pinreg_34_ | n1716);
  assign n1878 = (~Pinreg_50_ | n1715) & (~Pinreg_42_ | n1716);
  assign n1879 = (~Pinreg_50_ | n1716) & (~Pdata_in_1_ | n1715);
  assign n1880 = (~Pinreg_1_ | n1715) & (~Pdata_in_1_ | n1716);
  assign n1881 = (~Pinreg_9_ | n1715) & (~Pinreg_1_ | n1716);
  assign n1882 = (~Pinreg_17_ | n1715) & (~Pinreg_9_ | n1716);
  assign n1883 = (~Pinreg_25_ | n1715) & (~Pinreg_17_ | n1716);
  assign n1884 = (~Pinreg_33_ | n1715) & (~Pinreg_25_ | n1716);
  assign n1885 = (~Pinreg_41_ | n1715) & (~Pinreg_33_ | n1716);
  assign n1886 = (~Pinreg_49_ | n1715) & (~Pinreg_41_ | n1716);
  assign n1887 = (~Pinreg_49_ | n1716) & (~Pdata_in_0_ | n1715);
  assign n1888 = (~Pinreg_0_ | n1715) & (~Pdata_in_0_ | n1716);
  assign n1889 = (~Pinreg_8_ | n1715) & (~Pinreg_0_ | n1716);
  assign n1890 = (~Pinreg_16_ | n1715) & (~Pinreg_8_ | n1716);
  assign n1891 = (~Pinreg_24_ | n1715) & (~Pinreg_16_ | n1716);
  assign n1892 = (~Pinreg_32_ | n1715) & (~Pinreg_24_ | n1716);
  assign n1893 = (~Pinreg_40_ | n1715) & (~Pinreg_32_ | n1716);
  assign n1894 = (~Pinreg_48_ | n1715) & (~Pinreg_40_ | n1716);
  assign n1895 = (~Pinreg_54_ | n1716) & (~Pdata_in_3_ | n1715);
  assign n1896 = (~Pinreg_3_ | n1715) & (~Pdata_in_3_ | n1716);
  assign n1897 = (~Pinreg_11_ | n1715) & (~Pinreg_3_ | n1716);
  assign n1898 = (~Pinreg_19_ | n1715) & (~Pinreg_11_ | n1716);
  assign n1899 = (~Pinreg_19_ | n1716) & (~Pdata_in_4_ | n1715);
  assign n1900 = (~Pinreg_4_ | n1715) & (~Pdata_in_4_ | n1716);
  assign n1901 = (~Pinreg_12_ | n1715) & (~Pinreg_4_ | n1716);
  assign n1902 = (~Pinreg_20_ | n1715) & (~Pinreg_12_ | n1716);
  assign n1903 = (~Pinreg_28_ | n1715) & (~Pinreg_20_ | n1716);
  assign n1904 = (~Pinreg_36_ | n1715) & (~Pinreg_28_ | n1716);
  assign n1905 = (~Pinreg_44_ | n1715) & (~Pinreg_36_ | n1716);
  assign n1906 = (~Pinreg_52_ | n1715) & (~Pinreg_44_ | n1716);
  assign n1907 = (~Pinreg_52_ | n1716) & (~Pdata_in_5_ | n1715);
  assign n1908 = (~Pinreg_5_ | n1715) & (~Pdata_in_5_ | n1716);
  assign n1909 = (~Pinreg_13_ | n1715) & (~Pinreg_5_ | n1716);
  assign n1910 = (~Pinreg_21_ | n1715) & (~Pinreg_13_ | n1716);
  assign n1911 = (~Pinreg_29_ | n1715) & (~Pinreg_21_ | n1716);
  assign n1912 = (~Pinreg_37_ | n1715) & (~Pinreg_29_ | n1716);
  assign n1913 = (~Pinreg_45_ | n1715) & (~Pinreg_37_ | n1716);
  assign n1914 = (~Pinreg_53_ | n1715) & (~Pinreg_45_ | n1716);
  assign n1915 = (~Pinreg_53_ | n1716) & (~Pdata_in_6_ | n1715);
  assign n1916 = (~Pinreg_6_ | n1715) & (~Pdata_in_6_ | n1716);
  assign n1917 = (~Pinreg_14_ | n1715) & (~Pinreg_6_ | n1716);
  assign n1918 = (~Pinreg_22_ | n1715) & (~Pinreg_14_ | n1716);
  assign n1919 = (~Pinreg_30_ | n1715) & (~Pinreg_22_ | n1716);
  assign n1920 = (~Pinreg_38_ | n1715) & (~Pinreg_30_ | n1716);
  assign n1921 = (~Pinreg_46_ | n1715) & (~Pinreg_38_ | n1716);
  assign n1922 = (~Pinreg_54_ | n1715) & (~Pinreg_46_ | n1716);
  assign n1923 = ~n932 | n915 | n916;
  assign n1924 = ~n1338 & (n919 | n922 | ~n1719);
  assign n1925 = ~n906 & (~n900 | n912 | n916);
  assign n1926 = ~n906 & (~n921 | n1338);
  assign n1927 = ~n1635 & (~n1723 | (~n951 & ~n981));
  assign n1928 = n958 & n1635 & (~n951 | ~n1666);
  assign n1929 = n1078 & (~n1064 | (n1351 & n1675));
  assign n1930 = ~n1062 | ~n1078 | ~n1351 | ~n1677;
  assign n1931 = n1201 | n1103 | n1686;
  assign n1932 = ~n1201 & (n1106 | (~n1117 & n1132));
  assign n1933 = n1201 & (~n1832 | (~n1638 & n1683));
  assign n1934 = ~n1201 & (n1134 | (n1640 & n1681));
  assign n1935 = (n1308 & ~n1633) | (n896 & (n1308 | n1633));
  assign n1936 = n1397 & (n1652 | (n892 & n887));
  assign n1937 = n872 & (~n1725 | (n893 & n897));
  assign n1938 = n1935 & ~n872 & ~n1398;
  assign n1939 = n1160 | ~n1666;
  assign n1940 = ~n1635 & (n1162 | (n958 & n1939));
  assign n1941 = ~n1635 | n975 | n980;
  assign n1942 = n1702 | ~n1173 | ~n1694;
  assign n1943 = n1696 | n1201 | ~n1681;
  assign n1944 = ~n1638 & (~n1727 | (n1639 & n1683));
  assign n1945 = ~n1638 | ~n1696 | n1103 | ~n1201;
  assign n1946 = ~n1078 | n1347 | ~n1349;
  assign n1947 = n993 & ~n1039;
  assign n1948 = ~n993 & (n1017 | n1044);
  assign n1949 = n1947 | n1948 | ~n1146 | ~n1149;
  assign n1950 = n1351 & n1349;
  assign n1951 = ~n1078 & (n1950 | (n1352 & n1677));
  assign n1952 = ~n1256 | ~n1281 | ~n1315 | ~n1382;
  assign n1953 = ~n1702 & (n1304 | (n1298 & n1358));
  assign n1954 = ~n1702 | ~n1358 | ~n1642;
  assign n1955 = ~n1292 & ~n1641 & (n1301 | n1691);
  assign n1956 = ~n1641 | n1701;
  assign n1957 = n872 & (~n1853 | (n893 & n1651));
  assign n1958 = ~n872 & (n1142 | n1309 | n1310);
  assign n1959 = n1281 & (~n1855 | (n1325 & ~n1697));
  assign n1960 = ~n1281 & (~n1977 | (n1315 & ~n1697));
  assign n1961 = n914 & n911;
  assign n1962 = ~n914 & (~n913 | n916);
  assign n1963 = ~n1338 & (n1658 | (n921 & n926));
  assign n1964 = n1078 & (~n1858 | (~n1073 & n1672));
  assign n1965 = ~n1078 & (~n1090 | n1350 | n1353);
  assign n1966 = ~n1190 | n1299 | n1300;
  assign n1967 = n1265 | n1276 | n1282 | ~n1285;
  assign n1968 = n1276 & n1705 & (n1377 | ~n1384);
  assign n1969 = ~n1271 | n1272;
  assign n1970 = ~n1271 & (n1327 | (n1316 & n1325));
  assign n1971 = (n872 & n1650) | (n1649 & (~n872 | n1650));
  assign n1972 = (n1633 & n1971) | (n878 & (~n1633 | n1971));
  assign n1973 = (~n872 & ~n1731) | (~n1730 & (n872 | ~n1731));
  assign n1974 = Pcount_2_ | ~Pcount_1_ | ~Pcount_0_ | n1404;
  assign n1975 = n1404 | Pcount_1_ | ~Pcount_0_;
  assign n1976 = ~Pcount_1_ & (Pcount_3_ | Pcount_2_);
  assign n1977 = ~n1256 | n1262;
  assign n1978 = n1802 & n891 & n886 & n875 & n882 & ~n895 & ~n898 & n1801;
  assign n1979 = ~n1928 & ~n1927 & n1806 & n963 & n1033;
  assign n1980 = n1668 & n1029 & ~n985 & n984 & ~n982 & n979 & n963 & n966;
  assign n1981 = n1058 & n1055 & ~n1052 & n1045 & n1043 & n999 & n1014 & n1048;
  assign n1982 = n1833 & n1131 & n1110 & n1113 & ~n1933 & ~n1934;
  assign n1983 = ~n875 | n877 | ~n882 | ~n1139 | n1937 | n1938 | n1141 | n1143;
  assign n1984 = n1941 & ~n1940 & n1669 & n1166 & ~n1164 & n979 & n963 & n969;
  assign n1985 = n1839 & n1131 & n1107 & n1122 & ~n1944 & n1945;
  assign n1986 = n1848 & n1706 & n1699 & n1278 & ~n1288 & n1289;
  assign n1987 = n1956 & ~n1955 & n1851 & n1703 & n1171 & n1183 & ~n1953 & n1954;
  assign n1988 = n1704 & n1312 & n873 & n882 & ~n1957 & ~n1958;
  assign n1989 = n1959 | n1960 | n1328 | ~n1386 | ~n1255 | ~n1322 | ~n1324 | n1326;
  assign n1990 = n1646 & n912 & ~n915 & ~n916;
  assign n1991 = n1859 & n1678 & n1070 & n1221 & ~n1964 & ~n1965;
  assign n1992 = n1362 | n1700 | ~n1703 | ~n1861 | ~n1193 | n1356 | n1357 | n1360;
  assign n1993 = n1862 & n1703 & ~n1373 & n1372 & n1178 & n1183;
  assign n1994 = n1977 & ~n1970 & n1967 & n1699 & n1320 & n1378 & ~n1968 & n1969;
  assign n1995 = n1973 & n1704 & n1400 & n875 & ~n1396 & n1399;
  assign n1996 = ~Pdata_2_ ^ ~n1983;
  assign n1997 = ~Pdata_5_ ^ ~n1989;
  assign n1998 = ~Pdata_6_ ^ ~n1992;
endmodule


