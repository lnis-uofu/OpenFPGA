*****************************
*     FPGA SPICE Netlist    *
* Description: Channel X-direction  [1][0] in FPGA *
*    Author: Xifan TANG     *
* Organization: EPFL/IC/LSI *
* Date: Thu Nov 15 14:26:08 2018
 *
*****************************
***** Subckt for Channel X [1][0] *****
.subckt chanx[1][0] 
+ in0 out1 in2 out3 in4 out5 in6 out7 in8 out9 in10 out11 in12 out13 in14 out15 in16 out17 in18 out19 in20 out21 in22 out23 in24 out25 in26 out27 in28 out29 in30 out31 in32 out33 in34 out35 in36 out37 in38 out39 in40 out41 in42 out43 in44 out45 in46 out47 in48 out49 in50 out51 in52 out53 in54 out55 in56 out57 in58 out59 in60 out61 in62 out63 in64 out65 in66 out67 in68 out69 in70 out71 in72 out73 in74 out75 in76 out77 in78 out79 in80 out81 in82 out83 in84 out85 in86 out87 in88 out89 in90 out91 in92 out93 in94 out95 in96 out97 in98 out99 
+ out0 in1 out2 in3 out4 in5 out6 in7 out8 in9 out10 in11 out12 in13 out14 in15 out16 in17 out18 in19 out20 in21 out22 in23 out24 in25 out26 in27 out28 in29 out30 in31 out32 in33 out34 in35 out36 in37 out38 in39 out40 in41 out42 in43 out44 in45 out46 in47 out48 in49 out50 in51 out52 in53 out54 in55 out56 in57 out58 in59 out60 in61 out62 in63 out64 in65 out66 in67 out68 in69 out70 in71 out72 in73 out74 in75 out76 in77 out78 in79 out80 in81 out82 in83 out84 in85 out86 in87 out88 in89 out90 in91 out92 in93 out94 in95 out96 in97 out98 in99 
+ mid_out0 mid_out1 mid_out2 mid_out3 mid_out4 mid_out5 mid_out6 mid_out7 mid_out8 mid_out9 mid_out10 mid_out11 mid_out12 mid_out13 mid_out14 mid_out15 mid_out16 mid_out17 mid_out18 mid_out19 mid_out20 mid_out21 mid_out22 mid_out23 mid_out24 mid_out25 mid_out26 mid_out27 mid_out28 mid_out29 mid_out30 mid_out31 mid_out32 mid_out33 mid_out34 mid_out35 mid_out36 mid_out37 mid_out38 mid_out39 mid_out40 mid_out41 mid_out42 mid_out43 mid_out44 mid_out45 mid_out46 mid_out47 mid_out48 mid_out49 mid_out50 mid_out51 mid_out52 mid_out53 mid_out54 mid_out55 mid_out56 mid_out57 mid_out58 mid_out59 mid_out60 mid_out61 mid_out62 mid_out63 mid_out64 mid_out65 mid_out66 mid_out67 mid_out68 mid_out69 mid_out70 mid_out71 mid_out72 mid_out73 mid_out74 mid_out75 mid_out76 mid_out77 mid_out78 mid_out79 mid_out80 mid_out81 mid_out82 mid_out83 mid_out84 mid_out85 mid_out86 mid_out87 mid_out88 mid_out89 mid_out90 mid_out91 mid_out92 mid_out93 mid_out94 mid_out95 mid_out96 mid_out97 mid_out98 mid_out99 
+ svdd sgnd
Xtrack_seg[0] in0 out0 mid_out0 svdd sgnd chan_segment_seg0
Xtrack_seg[1] in1 out1 mid_out1 svdd sgnd chan_segment_seg0
Xtrack_seg[2] in2 out2 mid_out2 svdd sgnd chan_segment_seg0
Xtrack_seg[3] in3 out3 mid_out3 svdd sgnd chan_segment_seg0
Xtrack_seg[4] in4 out4 mid_out4 svdd sgnd chan_segment_seg0
Xtrack_seg[5] in5 out5 mid_out5 svdd sgnd chan_segment_seg0
Xtrack_seg[6] in6 out6 mid_out6 svdd sgnd chan_segment_seg0
Xtrack_seg[7] in7 out7 mid_out7 svdd sgnd chan_segment_seg0
Xtrack_seg[8] in8 out8 mid_out8 svdd sgnd chan_segment_seg0
Xtrack_seg[9] in9 out9 mid_out9 svdd sgnd chan_segment_seg0
Xtrack_seg[10] in10 out10 mid_out10 svdd sgnd chan_segment_seg0
Xtrack_seg[11] in11 out11 mid_out11 svdd sgnd chan_segment_seg0
Xtrack_seg[12] in12 out12 mid_out12 svdd sgnd chan_segment_seg0
Xtrack_seg[13] in13 out13 mid_out13 svdd sgnd chan_segment_seg0
Xtrack_seg[14] in14 out14 mid_out14 svdd sgnd chan_segment_seg0
Xtrack_seg[15] in15 out15 mid_out15 svdd sgnd chan_segment_seg0
Xtrack_seg[16] in16 out16 mid_out16 svdd sgnd chan_segment_seg0
Xtrack_seg[17] in17 out17 mid_out17 svdd sgnd chan_segment_seg0
Xtrack_seg[18] in18 out18 mid_out18 svdd sgnd chan_segment_seg0
Xtrack_seg[19] in19 out19 mid_out19 svdd sgnd chan_segment_seg0
Xtrack_seg[20] in20 out20 mid_out20 svdd sgnd chan_segment_seg0
Xtrack_seg[21] in21 out21 mid_out21 svdd sgnd chan_segment_seg0
Xtrack_seg[22] in22 out22 mid_out22 svdd sgnd chan_segment_seg0
Xtrack_seg[23] in23 out23 mid_out23 svdd sgnd chan_segment_seg0
Xtrack_seg[24] in24 out24 mid_out24 svdd sgnd chan_segment_seg0
Xtrack_seg[25] in25 out25 mid_out25 svdd sgnd chan_segment_seg0
Xtrack_seg[26] in26 out26 mid_out26 svdd sgnd chan_segment_seg0
Xtrack_seg[27] in27 out27 mid_out27 svdd sgnd chan_segment_seg0
Xtrack_seg[28] in28 out28 mid_out28 svdd sgnd chan_segment_seg0
Xtrack_seg[29] in29 out29 mid_out29 svdd sgnd chan_segment_seg0
Xtrack_seg[30] in30 out30 mid_out30 svdd sgnd chan_segment_seg0
Xtrack_seg[31] in31 out31 mid_out31 svdd sgnd chan_segment_seg0
Xtrack_seg[32] in32 out32 mid_out32 svdd sgnd chan_segment_seg0
Xtrack_seg[33] in33 out33 mid_out33 svdd sgnd chan_segment_seg0
Xtrack_seg[34] in34 out34 mid_out34 svdd sgnd chan_segment_seg0
Xtrack_seg[35] in35 out35 mid_out35 svdd sgnd chan_segment_seg0
Xtrack_seg[36] in36 out36 mid_out36 svdd sgnd chan_segment_seg0
Xtrack_seg[37] in37 out37 mid_out37 svdd sgnd chan_segment_seg0
Xtrack_seg[38] in38 out38 mid_out38 svdd sgnd chan_segment_seg0
Xtrack_seg[39] in39 out39 mid_out39 svdd sgnd chan_segment_seg0
Xtrack_seg[40] in40 out40 mid_out40 svdd sgnd chan_segment_seg1
Xtrack_seg[41] in41 out41 mid_out41 svdd sgnd chan_segment_seg1
Xtrack_seg[42] in42 out42 mid_out42 svdd sgnd chan_segment_seg1
Xtrack_seg[43] in43 out43 mid_out43 svdd sgnd chan_segment_seg1
Xtrack_seg[44] in44 out44 mid_out44 svdd sgnd chan_segment_seg1
Xtrack_seg[45] in45 out45 mid_out45 svdd sgnd chan_segment_seg1
Xtrack_seg[46] in46 out46 mid_out46 svdd sgnd chan_segment_seg1
Xtrack_seg[47] in47 out47 mid_out47 svdd sgnd chan_segment_seg1
Xtrack_seg[48] in48 out48 mid_out48 svdd sgnd chan_segment_seg1
Xtrack_seg[49] in49 out49 mid_out49 svdd sgnd chan_segment_seg1
Xtrack_seg[50] in50 out50 mid_out50 svdd sgnd chan_segment_seg1
Xtrack_seg[51] in51 out51 mid_out51 svdd sgnd chan_segment_seg1
Xtrack_seg[52] in52 out52 mid_out52 svdd sgnd chan_segment_seg1
Xtrack_seg[53] in53 out53 mid_out53 svdd sgnd chan_segment_seg1
Xtrack_seg[54] in54 out54 mid_out54 svdd sgnd chan_segment_seg1
Xtrack_seg[55] in55 out55 mid_out55 svdd sgnd chan_segment_seg1
Xtrack_seg[56] in56 out56 mid_out56 svdd sgnd chan_segment_seg1
Xtrack_seg[57] in57 out57 mid_out57 svdd sgnd chan_segment_seg1
Xtrack_seg[58] in58 out58 mid_out58 svdd sgnd chan_segment_seg1
Xtrack_seg[59] in59 out59 mid_out59 svdd sgnd chan_segment_seg1
Xtrack_seg[60] in60 out60 mid_out60 svdd sgnd chan_segment_seg1
Xtrack_seg[61] in61 out61 mid_out61 svdd sgnd chan_segment_seg1
Xtrack_seg[62] in62 out62 mid_out62 svdd sgnd chan_segment_seg1
Xtrack_seg[63] in63 out63 mid_out63 svdd sgnd chan_segment_seg1
Xtrack_seg[64] in64 out64 mid_out64 svdd sgnd chan_segment_seg1
Xtrack_seg[65] in65 out65 mid_out65 svdd sgnd chan_segment_seg1
Xtrack_seg[66] in66 out66 mid_out66 svdd sgnd chan_segment_seg1
Xtrack_seg[67] in67 out67 mid_out67 svdd sgnd chan_segment_seg1
Xtrack_seg[68] in68 out68 mid_out68 svdd sgnd chan_segment_seg1
Xtrack_seg[69] in69 out69 mid_out69 svdd sgnd chan_segment_seg1
Xtrack_seg[70] in70 out70 mid_out70 svdd sgnd chan_segment_seg2
Xtrack_seg[71] in71 out71 mid_out71 svdd sgnd chan_segment_seg2
Xtrack_seg[72] in72 out72 mid_out72 svdd sgnd chan_segment_seg2
Xtrack_seg[73] in73 out73 mid_out73 svdd sgnd chan_segment_seg2
Xtrack_seg[74] in74 out74 mid_out74 svdd sgnd chan_segment_seg2
Xtrack_seg[75] in75 out75 mid_out75 svdd sgnd chan_segment_seg2
Xtrack_seg[76] in76 out76 mid_out76 svdd sgnd chan_segment_seg2
Xtrack_seg[77] in77 out77 mid_out77 svdd sgnd chan_segment_seg2
Xtrack_seg[78] in78 out78 mid_out78 svdd sgnd chan_segment_seg2
Xtrack_seg[79] in79 out79 mid_out79 svdd sgnd chan_segment_seg2
Xtrack_seg[80] in80 out80 mid_out80 svdd sgnd chan_segment_seg2
Xtrack_seg[81] in81 out81 mid_out81 svdd sgnd chan_segment_seg2
Xtrack_seg[82] in82 out82 mid_out82 svdd sgnd chan_segment_seg2
Xtrack_seg[83] in83 out83 mid_out83 svdd sgnd chan_segment_seg2
Xtrack_seg[84] in84 out84 mid_out84 svdd sgnd chan_segment_seg2
Xtrack_seg[85] in85 out85 mid_out85 svdd sgnd chan_segment_seg2
Xtrack_seg[86] in86 out86 mid_out86 svdd sgnd chan_segment_seg2
Xtrack_seg[87] in87 out87 mid_out87 svdd sgnd chan_segment_seg2
Xtrack_seg[88] in88 out88 mid_out88 svdd sgnd chan_segment_seg2
Xtrack_seg[89] in89 out89 mid_out89 svdd sgnd chan_segment_seg2
Xtrack_seg[90] in90 out90 mid_out90 svdd sgnd chan_segment_seg2
Xtrack_seg[91] in91 out91 mid_out91 svdd sgnd chan_segment_seg2
Xtrack_seg[92] in92 out92 mid_out92 svdd sgnd chan_segment_seg2
Xtrack_seg[93] in93 out93 mid_out93 svdd sgnd chan_segment_seg2
Xtrack_seg[94] in94 out94 mid_out94 svdd sgnd chan_segment_seg2
Xtrack_seg[95] in95 out95 mid_out95 svdd sgnd chan_segment_seg2
Xtrack_seg[96] in96 out96 mid_out96 svdd sgnd chan_segment_seg2
Xtrack_seg[97] in97 out97 mid_out97 svdd sgnd chan_segment_seg2
Xtrack_seg[98] in98 out98 mid_out98 svdd sgnd chan_segment_seg2
Xtrack_seg[99] in99 out99 mid_out99 svdd sgnd chan_segment_seg2
.eom
