// Benchmark "TOP" written by ABC on Tue Mar  5 10:05:28 2019

module s38584 ( clk, 
    Pg6753, Pg6752, Pg6751, Pg6750, Pg6749, Pg6748, Pg6747, Pg6746, Pg6745,
    Pg6744, Pg135, Pg134, Pg127, Pg126, Pg125, Pg124, Pg120, Pg116, Pg115,
    Pg114, Pg113, Pg100, Pg99, Pg92, Pg91, Pg90, Pg84, Pg73, Pg72, Pg64,
    Pg57, Pg56, Pg54, Pg53, Pg44, Pg36, Pg35, Pg5, 
    Pg34972, Pg34956, Pg34927, Pg34925, Pg34923, Pg34921, Pg34919, Pg34917,
    Pg34915, Pg34913, Pg34839, Pg34788, Pg34597, Pg34437, Pg34436, Pg34435,
    Pg34425, Pg34383, Pg34240, Pg34239, Pg34238, Pg34237, Pg34236, Pg34235,
    Pg34234, Pg34233, Pg34232, Pg34221, Pg34201, Pg33959, Pg33950, Pg33949,
    Pg33948, Pg33947, Pg33946, Pg33945, Pg33935, Pg33894, Pg33874, Pg33659,
    Pg33636, Pg33533, Pg33435, Pg33079, Pg32975, Pg32454, Pg32429, Pg32185,
    Pg31863, Pg31862, Pg31861, Pg31860, Pg31793, Pg31665, Pg31656, Pg31521,
    Pg30332, Pg30331, Pg30330, Pg30329, Pg30327, Pg29221, Pg29220, Pg29219,
    Pg29218, Pg29217, Pg29216, Pg29215, Pg29214, Pg29213, Pg29212, Pg29211,
    Pg29210, Pg28753, Pg28042, Pg28041, Pg28030, Pg27831, Pg26877, Pg26876,
    Pg26875, Pg26801, Pg25590, Pg25589, Pg25588, Pg25587, Pg25586, Pg25585,
    Pg25584, Pg25583, Pg25582, Pg25259, Pg25219, Pg25167, Pg25114, Pg24185,
    Pg24184, Pg24183, Pg24182, Pg24181, Pg24180, Pg24179, Pg24178, Pg24177,
    Pg24176, Pg24175, Pg24174, Pg24173, Pg24172, Pg24171, Pg24170, Pg24169,
    Pg24168, Pg24167, Pg24166, Pg24165, Pg24164, Pg24163, Pg24162, Pg24161,
    Pg24151, Pg23759, Pg23683, Pg23652, Pg23612, Pg23190, Pg23002, Pg21727,
    Pg21698, Pg21292, Pg21270, Pg21245, Pg21176, Pg20901, Pg20899, Pg20763,
    Pg20654, Pg20652, Pg20557, Pg20049, Pg19357, Pg19334, Pg18881, Pg18101,
    Pg18100, Pg18099, Pg18098, Pg18097, Pg18096, Pg18095, Pg18094, Pg18092,
    Pg17871, Pg17845, Pg17819, Pg17813, Pg17787, Pg17778, Pg17764, Pg17760,
    Pg17743, Pg17739, Pg17722, Pg17715, Pg17711, Pg17688, Pg17685, Pg17678,
    Pg17674, Pg17649, Pg17646, Pg17639, Pg17607, Pg17604, Pg17580, Pg17577,
    Pg17519, Pg17423, Pg17404, Pg17400, Pg17320, Pg17316, Pg17291, Pg16955,
    Pg16924, Pg16874, Pg16775, Pg16748, Pg16744, Pg16722, Pg16718, Pg16693,
    Pg16686, Pg16659, Pg16656, Pg16627, Pg16624, Pg16603, Pg14828, Pg14779,
    Pg14749, Pg14738, Pg14705, Pg14694, Pg14673, Pg14662, Pg14635, Pg14597,
    Pg14518, Pg14451, Pg14421, Pg14217, Pg14201, Pg14189, Pg14167, Pg14147,
    Pg14125, Pg14096, Pg13966, Pg13926, Pg13906, Pg13895, Pg13881, Pg13865,
    Pg13272, Pg13259, Pg13099, Pg13085, Pg13068, Pg13049, Pg13039, Pg12923,
    Pg12919, Pg12833, Pg12832, Pg12470, Pg12422, Pg12368, Pg12350, Pg12300,
    Pg12238, Pg12184, Pg11770, Pg11678, Pg11447, Pg11418, Pg11388, Pg11349,
    Pg10527, Pg10500, Pg10306, Pg10122, Pg9817, Pg9743, Pg9741, Pg9682,
    Pg9680, Pg9617, Pg9615, Pg9555, Pg9553, Pg9497, Pg9251, Pg9048, Pg9019,
    Pg8920, Pg8919, Pg8918, Pg8917, Pg8916, Pg8915, Pg8870, Pg8839, Pg8789,
    Pg8788, Pg8787, Pg8786, Pg8785, Pg8784, Pg8783, Pg8719, Pg8475, Pg8416,
    Pg8403, Pg8398, Pg8358, Pg8353, Pg8344, Pg8342, Pg8291, Pg8283, Pg8279,
    Pg8277, Pg8235, Pg8215, Pg8178, Pg8132, Pg7946, Pg7916, Pg7540, Pg7260,
    Pg7257, Pg7245, Pg7243  );
  input  Pg6753, Pg6752, Pg6751, Pg6750, Pg6749, Pg6748, Pg6747, Pg6746,
    Pg6745, Pg6744, Pg135, Pg134, Pg127, Pg126, Pg125, Pg124, Pg120, Pg116,
    Pg115, Pg114, Pg113, Pg100, Pg99, Pg92, Pg91, Pg90, Pg84, Pg73, Pg72,
    Pg64, Pg57, Pg56, Pg54, Pg53, Pg44, Pg36, Pg35, Pg5, clk;
  output Pg34972, Pg34956, Pg34927, Pg34925, Pg34923, Pg34921, Pg34919,
    Pg34917, Pg34915, Pg34913, Pg34839, Pg34788, Pg34597, Pg34437, Pg34436,
    Pg34435, Pg34425, Pg34383, Pg34240, Pg34239, Pg34238, Pg34237, Pg34236,
    Pg34235, Pg34234, Pg34233, Pg34232, Pg34221, Pg34201, Pg33959, Pg33950,
    Pg33949, Pg33948, Pg33947, Pg33946, Pg33945, Pg33935, Pg33894, Pg33874,
    Pg33659, Pg33636, Pg33533, Pg33435, Pg33079, Pg32975, Pg32454, Pg32429,
    Pg32185, Pg31863, Pg31862, Pg31861, Pg31860, Pg31793, Pg31665, Pg31656,
    Pg31521, Pg30332, Pg30331, Pg30330, Pg30329, Pg30327, Pg29221, Pg29220,
    Pg29219, Pg29218, Pg29217, Pg29216, Pg29215, Pg29214, Pg29213, Pg29212,
    Pg29211, Pg29210, Pg28753, Pg28042, Pg28041, Pg28030, Pg27831, Pg26877,
    Pg26876, Pg26875, Pg26801, Pg25590, Pg25589, Pg25588, Pg25587, Pg25586,
    Pg25585, Pg25584, Pg25583, Pg25582, Pg25259, Pg25219, Pg25167, Pg25114,
    Pg24185, Pg24184, Pg24183, Pg24182, Pg24181, Pg24180, Pg24179, Pg24178,
    Pg24177, Pg24176, Pg24175, Pg24174, Pg24173, Pg24172, Pg24171, Pg24170,
    Pg24169, Pg24168, Pg24167, Pg24166, Pg24165, Pg24164, Pg24163, Pg24162,
    Pg24161, Pg24151, Pg23759, Pg23683, Pg23652, Pg23612, Pg23190, Pg23002,
    Pg21727, Pg21698, Pg21292, Pg21270, Pg21245, Pg21176, Pg20901, Pg20899,
    Pg20763, Pg20654, Pg20652, Pg20557, Pg20049, Pg19357, Pg19334, Pg18881,
    Pg18101, Pg18100, Pg18099, Pg18098, Pg18097, Pg18096, Pg18095, Pg18094,
    Pg18092, Pg17871, Pg17845, Pg17819, Pg17813, Pg17787, Pg17778, Pg17764,
    Pg17760, Pg17743, Pg17739, Pg17722, Pg17715, Pg17711, Pg17688, Pg17685,
    Pg17678, Pg17674, Pg17649, Pg17646, Pg17639, Pg17607, Pg17604, Pg17580,
    Pg17577, Pg17519, Pg17423, Pg17404, Pg17400, Pg17320, Pg17316, Pg17291,
    Pg16955, Pg16924, Pg16874, Pg16775, Pg16748, Pg16744, Pg16722, Pg16718,
    Pg16693, Pg16686, Pg16659, Pg16656, Pg16627, Pg16624, Pg16603, Pg14828,
    Pg14779, Pg14749, Pg14738, Pg14705, Pg14694, Pg14673, Pg14662, Pg14635,
    Pg14597, Pg14518, Pg14451, Pg14421, Pg14217, Pg14201, Pg14189, Pg14167,
    Pg14147, Pg14125, Pg14096, Pg13966, Pg13926, Pg13906, Pg13895, Pg13881,
    Pg13865, Pg13272, Pg13259, Pg13099, Pg13085, Pg13068, Pg13049, Pg13039,
    Pg12923, Pg12919, Pg12833, Pg12832, Pg12470, Pg12422, Pg12368, Pg12350,
    Pg12300, Pg12238, Pg12184, Pg11770, Pg11678, Pg11447, Pg11418, Pg11388,
    Pg11349, Pg10527, Pg10500, Pg10306, Pg10122, Pg9817, Pg9743, Pg9741,
    Pg9682, Pg9680, Pg9617, Pg9615, Pg9555, Pg9553, Pg9497, Pg9251, Pg9048,
    Pg9019, Pg8920, Pg8919, Pg8918, Pg8917, Pg8916, Pg8915, Pg8870, Pg8839,
    Pg8789, Pg8788, Pg8787, Pg8786, Pg8785, Pg8784, Pg8783, Pg8719, Pg8475,
    Pg8416, Pg8403, Pg8398, Pg8358, Pg8353, Pg8344, Pg8342, Pg8291, Pg8283,
    Pg8279, Pg8277, Pg8235, Pg8215, Pg8178, Pg8132, Pg7946, Pg7916, Pg7540,
    Pg7260, Pg7257, Pg7245, Pg7243;
  reg Ng5057, Ng2771, Ng1882, Ng2299, Ng4040, Ng2547, Ng559, Ng3243, Ng452,
    Ng3542, Ng5232, Ng5813, Ng2907, Ng1744, Ng5909, Ng1802, Ng3554, Ng6219,
    Ng807, Ng6031, Ng847, Ng976, Ng4172, Ng4372, Ng3512, Ng749, Ng3490,
    Pg12350, Ng4235, Ng1600, Ng1714, Pg14451, Ng3155, Ng2236, Ng4555,
    Ng3698, Ng1736, Ng1968, Ng4621, Ng5607, Ng2657, Pg12300, Ng490, Ng311,
    Ng772, Ng5587, Ng6177, Ng6377, Ng3167, Ng5615, Ng4567, Ng3457, Ng6287,
    Pg7946, Ng2563, Ng4776, Ng4593, Ng6199, Ng2295, Ng1384, Ng1339, Ng5180,
    Ng2844, Ng1024, Ng5591, Ng3598, Ng4264, Ng767, Ng5853, Pg13865, Ng2089,
    Ng4933, Ng4521, Ng5507, Pg16656, Ng6291, Ng294, Ng5559, Pg9617, Pg9741,
    Ng3813, Ng562, Ng608, Ng1205, Ng3909, Ng6259, Ng5905, Ng921, Ng2955,
    Ng203, Ng1099, Ng4878, Ng5204, Pg17604, Ng3606, Ng1926, Ng6215, Ng3586,
    Ng291, Ng4674, Ng3570, Pg9048, Pg17607, Ng1862, Ng676, Ng843, Ng4332,
    Ng4153, Pg17711, Ng6336, Ng622, Ng3506, Ng4558, Pg17685, Ng3111,
    \[4430] , Ng26936, Ng939, Ng278, Ng4492, Ng4864, Ng1036, \[4427] ,
    Ng1178, Ng3239, Ng718, Ng6195, Ng1135, Ng6395, \[4415] , Ng554, Ng496,
    Ng3853, Ng5134, Pg17404, Pg8344, Ng2485, Ng925, Ng48, Ng5555, Pg14096,
    Ng1798, Ng4076, Ng2941, Ng3905, Ng763, Ng6255, Ng4375, Ng4871, Ng4722,
    Ng590, Pg13099, Ng1632, Pg12238, Ng3100, Ng1495, Ng1437, Ng6154,
    Ng1579, Ng5567, Ng1752, Ng1917, Ng744, Ng4737, \[4661] , Ng6267,
    Pg16659, Ng1442, Ng5965, Ng4477, Pg10500, Ng4643, Ng5264, Pg14779,
    Ng2610, Ng5160, Ng5933, Ng1454, Ng753, Ng1296, Ng3151, Ng2980, Ng6727,
    Ng3530, Ng4104, Ng1532, Pg9251, Ng2177, Ng52, Ng4754, Ng1189, Ng2287,
    Ng4273, Ng1389, Ng1706, Ng5835, Ng1171, Ng4269, Ng2399, Ng4983, Ng5611,
    Pg16627, Ng4572, Ng3143, Ng2898, Ng3343, Ng3235, Ng4543, Ng3566,
    Ng4534, Ng4961, Ng4927, Ng2259, Ng2819, Pg7257, Ng5802, Ng2852, Ng417,
    Ng681, Ng437, Ng351, Ng5901, Ng2886, Ng3494, Ng5511, Ng3518, Ng1604,
    Ng5092, Ng4831, Ng4382, Ng6386, Ng479, Ng3965, Ng4749, Ng2008, Ng736,
    Ng3933, Ng222, Ng3050, Ng1052, Pg17580, Ng2122, Ng2465, Ng5889, Ng4495,
    Pg8719, Ng4653, Ng3179, Ng1728, Ng2433, Ng3835, Ng6187, Ng4917, Ng1070,
    Ng822, Pg17715, Ng914, Ng5339, Ng4164, Ng969, Ng2807, Ng4054, Ng6191,
    Ng5077, Ng5523, Ng3680, Ng6637, Ng174, Ng1682, Ng355, Ng1087, Ng1105,
    Ng2342, Ng6307, Ng3802, Ng6159, Ng2255, Ng2815, Ng911, Ng43, Pg16775,
    Ng1748, Ng5551, Ng3558, Ng5499, Ng2960, Ng3901, Ng4888, Ng6251,
    Pg17649, Ng1373, Pg8215, Ng157, Ng2783, Ng4281, Ng3574, Ng2112, Ng1283,
    Ng433, Ng4297, Pg14738, Pg13272, Ng758, Ng4639, Ng6537, Ng5543, Pg8475,
    Ng5961, Ng6243, Ng632, Pg12919, Ng3889, Ng3476, Ng1664, Ng1246, Ng6629,
    Ng246, Ng4049, Pg7260, Ng2932, Ng4575, Ng4098, Ng4498, Ng528, Ng16,
    Ng3139, \[4432] , Ng4584, Ng142, Pg17639, Ng5831, Ng239, Ng1216,
    Ng2848, Ng5022, Pg16955, Ng1030, Pg13881, Ng3231, Pg9817, Ng1430,
    Ng4452, Ng2241, Ng1564, Pg9680, Ng6148, Ng6649, Ng110, Pg14147, Ng225,
    Ng4486, Ng4504, Ng5873, Ng5037, Ng2319, Ng5495, Pg11770, Ng5208,
    Ng5579, Ng5869, Ng1589, Ng5752, Ng6279, Ng5917, Ng2975, Ng6167,
    Pg13966, Ng2599, Ng1448, Pg14125, Ng2370, Ng5164, Ng1333, Ng153,
    Ng6549, Ng4087, Ng4801, Ng2984, Ng3961, Ng962, Ng101, Pg8918, Ng6625,
    Ng51, Ng1018, Pg17320, Ng4045, Ng1467, Ng2461, Ng2756, Ng5990, Ng1256,
    Ng5029, Ng6519, Ng1816, Ng4369, Ng4578, Ng4459, Ng3831, Ng2514, Ng3288,
    Ng2403, Ng2145, Ng1700, Ng513, Ng2841, Ng5297, Ng2763, Ng4793, Ng952,
    Ng1263, Ng1950, Ng5138, Ng2307, Ng5109, Pg8398, Ng4664, Ng2223, Ng5808,
    Ng6645, Ng2016, Ng3873, Pg13926, Ng2315, Ng2811, Ng5957, Ng2047,
    Ng3869, Pg17760, Ng5575, Ng46, Ng3752, Ng3917, Pg8783, Ng1585, Ng4388,
    Ng6275, Ng6311, Pg8916, Ng1041, Ng2595, Ng2537, \[4426] , Ng4430,
    Ng4564, Ng4826, Ng6239, Ng232, Ng5268, Ng6545, Ng2417, Ng1772, Ng5052,
    Pg9615, Ng1890, Ng2629, Ng572, Ng2130, Ng4108, Ng4308, Ng475, Ng990,
    Ng45, Pg12184, Ng3990, Ng5881, Ng1992, Ng3171, Ng812, Ng832, Ng5897,
    Ng4571, Pg13895, Ng4455, Ng2902, Ng333, Ng168, Ng2823, Ng3684, Ng3639,
    Pg14597, Ng3338, Ng5406, Ng269, Ng401, Ng6040, Ng441, Pg9553, Ng3808,
    Ng10384, Ng3957, Ng4093, Ng1760, Pg12422, Ng160, Ng2279, Ng3498, Ng586,
    Pg14201, Ng2619, Ng1183, Ng1608, Pg8785, Pg17577, Ng1779, Ng2652,
    Ng2193, Ng2393, Ng661, Ng4950, Ng5535, Ng2834, Ng1361, Ng6235, Ng1146,
    Ng2625, Ng150, Ng1696, Ng6555, Pg14189, Ng3881, Ng6621, Ng3470, Ng3897,
    Ng518, Ng538, Ng2606, Ng1472, Ng542, Ng5188, Ng5689, Pg13259, Ng405,
    Ng5216, Ng6494, Ng4669, Ng996, Ng4531, Ng2860, Ng4743, Ng6593, Pg8291,
    Ng4411, Ng1413, Ng26960, Pg13039, Ng6641, Ng1936, Ng55, Ng504, Ng2587,
    Ng4480, Ng2311, Ng3602, Ng5571, Ng3578, Pg9555, Ng5827, Ng3582, Ng6271,
    Ng4688, Ng2380, Ng5196, Ng3227, Ng2020, Pg14518, Pg17316, Ng6541,
    Ng3203, Ng1668, Ng4760, Ng262, Ng1840, Ng5467, Ng460, Ng6209, \[4436] ,
    Pg14662, Ng655, Ng3502, Ng2204, Ng5256, Ng4608, Ng794, Pg13906, Ng4423,
    Ng3689, Ng5685, Ng703, Ng862, Ng3247, Ng2040, Ng4146, Ng4633, Pg7916,
    Ng4732, Pg9497, Ng5817, Ng2351, Ng2648, Ng6736, Ng4944, Ng4072, Pg7540,
    Ng4443, Ng3466, Ng4116, Ng5041, Ng4434, Ng3827, Ng6500, Pg17813,
    Ng3133, Ng3333, Ng979, Ng4681, Ng298, Ng2667, Pg8789, Ng1894, Ng2988,
    Ng3538, Ng301, Ng341, Ng827, Pg17291, Ng2555, Ng5011, Ng199, Ng6523,
    Ng1526, Ng4601, Ng854, Ng1484, Ng4922, Ng5080, Ng5863, Ng4581, Ng2518,
    Ng2567, Ng568, Ng3263, Ng6613, Ng6044, Ng6444, Ng2965, Ng5857, Ng1616,
    Ng890, Pg17646, Ng3562, Pg10122, Ng1404, Ng3817, Ng93, Ng4501, Ng287,
    Ng2724, Ng4704, Ng22, Ng2878, Ng5220, Ng617, Pg12368, Ng316, Ng1277,
    Ng6513, Ng336, Ng2882, Ng933, Ng1906, Ng305, Ng8, Ng2799, Pg14167,
    Pg17787, Ng4912, Ng4157, Ng2541, Ng2153, Ng550, Ng255, Ng1945, Ng5240,
    Ng1478, Ng3863, Ng1959, Ng3480, Ng6653, Pg17764, Ng2864, Ng4894,
    Pg17678, Ng3857, Pg16693, Ng499, Ng1002, Ng776, Ng1236, Ng4646, Ng2476,
    Ng1657, Ng2375, Ng63, Pg17739, Ng358, Ng896, Ng283, Ng3161, Ng2384,
    Pg14828, Ng4616, Ng4561, Ng2024, Ng3451, Ng2795, Ng613, Ng4527, Ng1844,
    Ng5937, Ng4546, Ng2523, Pg11349, Ng2643, Ng1489, Pg8358, Ng2551,
    Ng5156, \[4421] , Pg8279, Pg8839, Ng1955, Ng6049, Ng2273, Pg14749,
    Ng4771, Ng6098, Ng3147, Ng3347, Ng2269, Ng191, Ng2712, Ng626, Ng2729,
    Ng5357, Ng4991, Pg17819, Ng4709, Ng2927, Ng4340, Ng5929, Ng4907,
    Pg16874, Ng4035, Ng2946, Ng918, Ng4082, Pg9743, Ng2036, Ng577, Ng1620,
    Ng2831, Ng667, Ng930, Ng3937, Ng817, Ng1249, Ng837, Pg16924, Ng599,
    Ng5475, Ng739, Ng5949, Ng6682, Ng904, Ng2873, Ng1854, Ng5084, Ng5603,
    Pg8870, Ng2495, Ng2437, Ng2102, Ng2208, Ng2579, Ng4064, Ng4899, Ng2719,
    Ng4785, Ng5583, Ng781, Ng6173, Pg17743, Ng2917, Ng686, Ng1252, Ng671,
    Ng2265, Ng6283, Pg14705, Pg17519, Pg8784, Ng5527, Ng4489, Ng1974,
    Ng1270, Ng4966, Ng6227, Ng3929, Ng5503, Ng4242, Ng5925, Ng1124, Ng4955,
    Ng5224, Ng2012, Ng6203, Ng5120, Pg17674, Ng2389, Ng4438, Ng2429,
    Ng2787, Ng1287, Ng2675, \[4507] , Ng4836, Ng1199, Pg19357, Ng5547,
    Ng2138, Pg16744, Ng2338, Pg8919, Ng6247, Ng2791, Ng3949, Ng1291,
    Ng5945, Ng5244, Ng2759, Ng6741, Ng785, Ng1259, Ng3484, Ng209, Ng6609,
    Ng5517, Ng2449, Ng2575, Ng65, Ng2715, Ng936, Ng2098, Ng4462, Ng604,
    Ng6589, Ng1886, Pg17845, Pg17871, Ng429, Ng1870, Ng4249, Ng1825,
    Ng1008, Ng4392, Ng3546, Ng5236, Ng1768, Ng4854, Ng3925, Ng6509, Ng732,
    Ng2504, Ng1322, Ng4520, Pg8917, Ng2185, Ng37, Ng4031, Ng2070, \[4658] ,
    Ng4176, Pg11418, Ng4405, Ng872, Ng6181, Ng6381, Ng4765, Ng5563, Ng1395,
    Ng1913, Ng2331, Ng6263, Ng50, Ng3945, Ng347, Ng4473, Ng1266, Ng5489,
    Ng714, Ng2748, Ng5471, Ng4540, Ng6723, Ng6605, Ng2445, Ng2173, Pg9019,
    Ng2491, Ng4849, Ng2169, Ng2283, Ng6585, \[4428] , Ng2407, Ng2868,
    Ng2767, Ng1783, Pg16718, Ng1312, Ng5212, Ng4245, Ng645, Ng4291,
    \[4435] , Ng182, Ng1129, Ng2227, Pg8788, Ng2246, Ng1830, Ng3590, Ng392,
    Ng1592, Ng6505, Ng1221, Ng5921, \[4431] , Ng146, Ng218, Ng1932, Ng1624,
    Ng5062, Ng5462, Ng2689, Ng6573, Ng1677, Ng2028, Ng2671, Pg10527,
    Pg7243, Ng1848, \[4434] , Ng5485, Ng2741, Pg11678, Ng2638, Ng4122,
    Ng4322, Ng5941, Ng2108, Pg13068, Ng25, Ng1644, Ng595, Ng2217, Ng1319,
    Ng2066, Ng1152, Ng5252, Ng2165, Ng2571, Ng5176, Pg14673, Ng1211,
    Ng2827, Pg14217, Ng4859, Ng424, Ng1274, Pg17423, Ng85, Ng2803, Ng1821,
    Ng2509, Ng5073, Ng1280, \[4651] , Pg13085, Ng6633, Ng5124, Pg17400,
    Ng6303, Ng5069, Ng2994, Ng650, Ng1636, Ng3921, Ng2093, Ng6732, Ng1306,
    Ng1061, Ng3462, Ng2181, Ng956, Ng1756, Ng5849, Ng4112, Ng2685, Ng2197,
    Ng2421, Ng1046, Ng482, Ng4401, Ng1514, Ng329, Ng6565, Ng2950, Ng1345,
    Ng6533, Pg14421, Ng4727, Pg12470, Ng1536, Ng3941, Ng370, Ng5694,
    Ng1858, Ng446, Ng3219, Ng1811, Ng6601, Ng2441, Ng1874, Ng4349, Ng6581,
    Ng6597, Ng3610, Ng2890, Ng1978, Ng1612, Ng112, Ng2856, Ng1982, Pg17722,
    Ng5228, Ng4119, Ng6390, Ng1542, Ng4258, Ng4818, Ng5033, Ng4717, Ng1554,
    Ng3849, Pg17778, Ng3199, Ng5845, Ng4975, Ng790, Ng5913, Ng1902, Ng6163,
    Ng4125, Ng4821, Ng4939, Pg19334, Ng3207, Ng4483, Ng3259, Ng5142,
    Ng5248, Ng2126, Ng3694, Ng5481, Ng1964, Ng5097, Ng3215, Pg16748, Ng111,
    Ng4427, Ng2779, Pg8786, Pg7245, Ng1720, Ng1367, Ng5112, Ng4145, Ng2161,
    Ng376, Ng2361, Pg11447, Ng582, Ng2051, Ng1193, Ng2327, Ng907, Ng947,
    Ng1834, Ng3594, Ng2999, Ng2303, Pg17688, Ng699, Ng723, Ng5703, Ng546,
    Ng2472, Ng5953, Pg8277, Ng1740, Ng3550, Ng3845, Ng2116, Pg14635,
    Ng3195, Ng3913, Pg10306, Ng1687, Ng2681, Ng2533, Ng324, Ng2697, Ng4417,
    Ng6561, Ng1141, Pg12923, Ng2413, Ng1710, Ng6527, Ng3255, Ng1691,
    Ng2936, Ng5644, Ng5152, Ng5352, Pg8915, Ng2775, Ng2922, Ng1111, Ng5893,
    Pg16603, Ng6617, Ng2060, Ng4512, Ng5599, Ng3401, Ng4366, Pg16722,
    \[4433] , Ng3129, Ng3329, Ng5170, Ng26959, Ng5821, Ng6299, Pg8416,
    Ng2079, Ng4698, Ng3703, Ng1559, Ng943, Ng411, Pg9682, Ng3953, Ng2704,
    Ng6035, Ng1300, Ng4057, Ng5200, Ng4843, Ng5046, Ng2250, Ng26885,
    Ng4549, Ng2453, Ng5841, Pg14694, Ng2912, Ng2357, Pg8920, Ng164, Ng4253,
    Ng5016, Ng3119, Ng1351, Ng1648, Ng6972, Ng5115, Ng3352, Ng6657, Ng4552,
    Ng3893, Ng3211, Pg13049, Pg16624, Ng5595, Ng3614, Ng2894, Ng3125,
    Pg16686, Ng3821, Ng4141, Ng6974, Ng5272, Ng2735, Ng728, Ng6295, Ng2661,
    Ng1988, Ng5128, Ng1548, Ng3106, Ng4659, Ng4358, Ng1792, Ng2084, Ng3187,
    Ng4311, Ng2583, Ng3003, Ng1094, Ng3841, Ng4284, Ng3191, Ng4239, Ng4180,
    Ng691, Ng534, Ng385, Ng2004, Ng2527, Ng5456, Ng4420, Ng5148, Ng4507,
    Ng5348, Ng3223, Ng2970, Ng5698, Ng5260, Ng1521, Ng3522, Ng3115, Ng3251,
    Pg12832, Ng4628, Ng1996, Pg8342, Ng4515, Pg8787, Ng4300, Ng1724,
    Ng1379, Pg11388, Ng1878, Ng5619, Ng71, \[4437] ;
  wire n4124_1, n4133, n4135, n4136, n4151_1, n4162, n4205, n4206_1, n4207,
    n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216_1, n4217,
    n4218, n4219, n4220, n4221, n4223, n4225, n4227, n4229, n4231, n4233,
    n4235, n4237, n4239, n4241, n4243, n4245, n4247, n4249_1, n4251, n4252,
    n4254_1, n4256, n4258, n4260, n4262, n4265, n4267, n4269, n4271, n4273,
    n4275, n4277, n4279, n4281, n4283, n4285, n4287, n4289, n4291, n4293,
    n4295, n4297, n4299, n4301, n4303, n4305, n4307, n4309, n4311, n4313,
    n4315, n4317, n4319, n4321, n4323, n4325, n4327, n4329, n4331, n4333,
    n4335, n4337, n4339, n4341, n4343, n4345, n4347, n4349, n4351, n4353,
    n4355, n4357, n4359, n4361, n4363, n4365, n4367, n4369_1, n4371, n4373,
    n4375, n4377, n4379, n4382, n4384, n4385, n4388, n4390, n4392, n4394,
    n4396, n4398, n4400, n4402, n4404, n4406, n4408, n4410, n4412, n4414,
    n4416, n4418, n4420, n4423, n4425, n4427, n4429, n4431, n4433, n4435,
    n4437_1, n4439, n4441, n4443, n4445, n4448, n4450, n4452_1, n4454,
    n4456_1, n4458, n4460_1, n4462, n4464, n4466, n4468, n4470_1, n4472,
    n4474, n4475_1, n4477, n4479, n4481, n4483, n4485_1, n4487, n4489_1,
    n4491, n4493, n4495_1, n4497, n4499_1, n4501, n4503, n4505, n4507,
    n4509, n4512, n4514_1, n4516, n4518, n4520, n4521, n4522, n4524_1,
    n4526, n4528, n4530, n4532, n4534_1, n4536, n4538, n4541, n4543, n4545,
    n4547, n4549_1, n4551, n4553, n4555, n4557, n4558, n4560, n4562, n4564,
    n4567, n4569, n4571, n4573, n4575, n4577, n4579, n4581, n4583, n4585,
    n4587, n4589, n4591, n4593, n4595, n4597, n4599, n4601, n4603, n4605,
    n4607_1, n4609, n4611, n4613, n4615, n4617_1, n4619, n4621, n4623,
    n4625, n4627_1, n4629, n4631_1, n4633, n4635, n4637, n4639, n4641,
    n4643, n4645, n4647, n4649, n4651, n4653, n4655, n4657, n4659, n4661,
    n4663, n4665, n4667, n4669, n4671, n4673, n4675, n4677, n4679, n4681,
    n4683, n4685, n4687_1, n4689, n4692, n4695, n4697, n4699, n4701, n4703,
    n4705, n4707, n4709, n4711, n4713, n4715, n4717, n4719, n4722, n4724,
    n4726, n4728, n4730, n4732, n4734, n4736, n4738, n4740, n4742, n4744,
    n4746_1, n4748, n4750, n4752, n4754, n4756_1, n4758, n4760, n4762,
    n4764, n4766_1, n4768, n4770, n4772, n4774, n4776, n4778, n4780,
    n4782_1, n4784, n4786, n4788, n4790, n4792, n4794, n4796, n4798, n4800,
    n4802_1, n4804, n4806, n4808, n4810, n4812_1, n4814, n4816, n4818,
    n4820, n4822_1, n4824, n4826, n4828, n4830, n4832, n4834, n4836, n4838,
    n4840, n4842, n4844, n4846, n4848, n4850, n4852, n4854, n4856, n4858,
    n4860, n4862, n4864, n4866, n4868, n4870, n4872, n4874, n4876, n4878,
    n4880, n4882_1, n4884, n4886, n4887, n4889, n4891, n4893, n4895, n4898,
    n4900, n4902, n4904_1, n4906, n4908, n4909, n4911, n4913, n4915, n4917,
    n4919, n4921, n4923, n4925, n4927, n4929, n4931, n4933, n4935, n4937,
    n4939_1, n4941, n4943, n4945, n4947, n4949, n4951, n4953, n4955, n4958,
    n4960, n4962, n4964, n4966, n4968, n4970, n4972, n4974, n4976, n4978_1,
    n4980, n4982, n4984, n4986, n4988, n4990, n4992_1, n4994, n4996, n4998,
    n5000, n5002_1, n5004, n5006, n5008, n5010, n5012, n5014, n5016_1,
    n5018, n5020, n5022, n5025, n5027, n5029, n5031, n5034, n5036_1, n5038,
    n5040, n5042, n5044, n5046, n5048, n5049, n5050, n5052, n5054, n5057,
    n5059, n5061, n5063, n5065, n5067, n5069_1, n5072, n5074, n5076, n5078,
    n5080, n5082, n5084, n5086, n5088, n5090, n5091, n5093, n5095, n5097,
    n5099, n5102, n5104, n5106, n5108, n5110, n5112, n5114, n5116_1, n5118,
    n5120, n5122, n5124, n5126_1, n5128, n5131_1, n5132, n5134, n5136,
    n5139, n5141_1, n5143, n5145, n5147, n5149, n5151, n5153, n5155, n5157,
    n5159, n5161, n5163, n5165, n5167, n5169, n5170, n5172, n5174, n5176,
    n5178, n5180, n5182, n5184, n5186, n5188, n5190, n5192, n5194, n5196,
    n5198, n5200, n5202, n5204, n5206, n5208, n5210, n5212, n5214, n5216,
    n5218, n5220, n5222, n5224, n5226, n5228, n5230, n5232, n5234, n5236,
    n5238, n5240, n5242, n5244, n5246, n5248, n5250, n5252, n5254, n5256,
    n5258, n5260, n5262, n5264, n5266, n5268, n5270, n5272, n5274, n5276,
    n5278, n5280, n5283, n5285, n5287, n5289, n5291, n5293, n5296, n5298_1,
    n5300, n5302, n5304, n5306, n5308, n5310, n5312, n5314, n5316, n5318_1,
    n5320, n5322_1, n5324, n5326, n5328, n5330, n5332, n5334, n5336, n5338,
    n5340, n5342, n5344, n5346, n5348, n5350, n5352, n5354, n5356, n5358,
    n5360, n5362, n5365, n5367, n5370, n5372, n5374, n5376, n5378, n5380,
    n5382, n5384, n5386, n5388, n5390, n5392, n5394, n5396, n5398, n5400,
    n5402, n5404, n5406, n5408, n5410, n5412, n5414, n5416_1, n5418, n5420,
    n5422, n5424, n5425, n5427, n5429, n5431, n5433, n5435, n5437, n5439,
    n5441, n5443, n5445, n5447, n5449, n5451, n5453, n5455, n5457, n5459,
    n5461_1, n5463, n5465, n5467, n5469, n5471, n5473, n5475, n5477, n5479,
    n5481, n5483, n5485, n5487, n5489, n5491, n5493, n5495, n5497, n5499,
    n5501, n5503, n5505, n5507, n5509, n5511, n5513, n5515, n5517, n5519,
    n5521, n5523, n5525, n5527, n5529, n5531, n5533, n5535, n5537, n5539,
    n5541, n5543, n5545, n5547, n5549, n5551, n5553, n5555, n5557, n5559,
    n5560, n5562, n5564, n5566, n5568, n5570, n5572, n5574, n5576, n5578,
    n5580, n5582, n5584, n5586, n5588, n5590, n5592, n5594, n5596, n5598_1,
    n5600, n5602, n5604, n5606, n5608, n5610, n5612, n5614, n5616, n5618,
    n5620, n5622, n5624, n5626, n5628_1, n5630, n5632, n5634, n5636,
    n5638_1, n5640, n5642, n5644, n5646, n5648, n5650, n5652, n5654, n5656,
    n5658, n5660, n5662_1, n5664, n5666, n5668, n5669, n5671_1, n5673,
    n5675, n5677, n5679, n5681, n5683, n5685, n5687, n5689, n5691, n5693,
    n5695_1, n5697, n5699, n5701, n5703, n5705, n5707, n5709, n5711, n5713,
    n5715, n5717, n5719, n5721, n5723, n5725, n5727, n5729, n5730, n5731,
    n5733, n5735, n5737, n5739, n5741, n5743, n5745, n5747, n5749, n5751,
    n5753_1, n5755, n5757, n5759, n5761, n5763_1, n5765, n5767, n5769,
    n5771, n5773, n5775, n5777, n5779, n5781, n5783, n5785, n5787, n5789,
    n5791_1, n5793, n5795, n5797, n5799, n5801_1, n5803, n5805, n5807,
    n5809, n5811_1, n5813, n5815, n5817, n5819, n5821, n5823, n5825, n5827,
    n5829, n5831, n5833, n5835, n5837, n5839, n5841, n5843, n5845, n5847,
    n5849, n5851, n5853, n5855, n5857, n5859_1, n5861, n5863, n5865, n5866,
    n5867, n5868, n5869_1, n5871, n5872, n5873, n5874_1, n5875, n5876,
    n5877, n5878, n5880, n5881, n5882, n5883, n5884_1, n5885, n5886, n5887,
    n5888, n5889, n5892, n5894, n5895, n5897, n5898_1, n5899, n5901, n5902,
    n5903, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5914,
    n5915, n5916, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
    n5926, n5927, n5929, n5930, n5931, n5933, n5934, n5935, n5936, n5938,
    n5939, n5940, n5941, n5942, n5944, n5945, n5947, n5948, n5949, n5950,
    n5951, n5952, n5953, n5954, n5956_1, n5957, n5958, n5959, n5960, n5961,
    n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
    n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
    n5982, n5983, n5984, n5985, n5988, n5989, n5990_1, n5991, n5992, n5993,
    n5994, n5995, n5996, n5997, n5998_1, n5999, n6000, n6001, n6002, n6003,
    n6004, n6005, n6006, n6007, n6008_1, n6009, n6010, n6011, n6012_1,
    n6013, n6014, n6015, n6016, n6017_1, n6018, n6019, n6020, n6021, n6022,
    n6023, n6024, n6025, n6026, n6027_1, n6028, n6029, n6030, n6031, n6032,
    n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042_1,
    n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
    n6053, n6054, n6055, n6056_1, n6057, n6058, n6059, n6060, n6061_1,
    n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
    n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081_1,
    n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091_1,
    n6092, n6093, n6094, n6095, n6096_1, n6097, n6098, n6099, n6100, n6101,
    n6102, n6103, n6104_1, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
    n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
    n6122, n6123, n6124, n6125, n6126, n6127_1, n6128, n6129, n6130, n6131,
    n6132, n6133, n6134, n6135, n6136, n6137_1, n6138, n6139, n6140, n6141,
    n6142_1, n6143, n6144, n6145, n6146, n6147_1, n6148, n6149, n6150,
    n6151, n6152_1, n6153, n6154, n6155, n6156_1, n6157, n6158, n6159,
    n6160_1, n6161, n6162, n6163, n6164, n6165_1, n6166, n6167, n6168,
    n6169_1, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
    n6179_1, n6180, n6181, n6182, n6183_1, n6184, n6185, n6186, n6187,
    n6188, n6189, n6190, n6191, n6192_1, n6193, n6194, n6195, n6196_1,
    n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206_1,
    n6207, n6208, n6209, n6210, n6211_1, n6212, n6213, n6214, n6215,
    n6216_1, n6217, n6218, n6219, n6220, n6221_1, n6222, n6223, n6224,
    n6225, n6226_1, n6227, n6228, n6229, n6230_1, n6231, n6232, n6233,
    n6234, n6235_1, n6236, n6237, n6238, n6239, n6240_1, n6241, n6242,
    n6243, n6244, n6245_1, n6246, n6247, n6248, n6249, n6250_1, n6251,
    n6252, n6253, n6254, n6255_1, n6256, n6257, n6258, n6259, n6260_1,
    n6261, n6262, n6263, n6264, n6265_1, n6266, n6267, n6268, n6269,
    n6270_1, n6271, n6272, n6273, n6274, n6275_1, n6276, n6277, n6278,
    n6279_1, n6280, n6281, n6282, n6283, n6284_1, n6285, n6286, n6287,
    n6288, n6289_1, n6290, n6291, n6292, n6293_1, n6294, n6295, n6296,
    n6297_1, n6298, n6299, n6300, n6301, n6302_1, n6303, n6304, n6305,
    n6306, n6307, n6308, n6309, n6310_1, n6311, n6312, n6313, n6314,
    n6315_1, n6316, n6317, n6318, n6319, n6320_1, n6321, n6322, n6323,
    n6324, n6325, n6326, n6327, n6328, n6329, n6330_1, n6331, n6332, n6333,
    n6334, n6335_1, n6336, n6337, n6338, n6339, n6340_1, n6341, n6342,
    n6343, n6344, n6345, n6346, n6347, n6348, n6349_1, n6350, n6351, n6352,
    n6353, n6354_1, n6355, n6356, n6357, n6358, n6359_1, n6360, n6361,
    n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369_1, n6370, n6371,
    n6372, n6373_1, n6374, n6375, n6376_1, n6377, n6378, n6379, n6380_1,
    n6381, n6382, n6383, n6384, n6385_1, n6386, n6387, n6388, n6389,
    n6390_1, n6391, n6392, n6393, n6394, n6395_1, n6396, n6397, n6398,
    n6399_1, n6400, n6401, n6402, n6403_1, n6404, n6405, n6406, n6407,
    n6408, n6409, n6410, n6411, n6412, n6413_1, n6414, n6415, n6416,
    n6417_1, n6418, n6419, n6420, n6421, n6422_1, n6423, n6424, n6425,
    n6426, n6427_1, n6428, n6429, n6430, n6431, n6432_1, n6433, n6434,
    n6435, n6436, n6437_1, n6438, n6439, n6440, n6441, n6442_1, n6443,
    n6444, n6445, n6446, n6447_1, n6448, n6449, n6450, n6451, n6452_1,
    n6453, n6454, n6455, n6456, n6457_1, n6458, n6459, n6460, n6461,
    n6462_1, n6463, n6464, n6465, n6466, n6467_1, n6468, n6469, n6470,
    n6471, n6472_1, n6473, n6474, n6475, n6476, n6477_1, n6478, n6479,
    n6480, n6481, n6482_1, n6483, n6484, n6485, n6486, n6487_1, n6488,
    n6489, n6490, n6491, n6492_1, n6493, n6494, n6495, n6496, n6497_1,
    n6498, n6499, n6500, n6501, n6502_1, n6503, n6504, n6505, n6506,
    n6507_1, n6508, n6509, n6510, n6511, n6512_1, n6513, n6514, n6515,
    n6516, n6517_1, n6518, n6519, n6520, n6521, n6522_1, n6523, n6524,
    n6525, n6526_1, n6527, n6528, n6529, n6530, n6531_1, n6532, n6533,
    n6534, n6535, n6536_1, n6537, n6538, n6539, n6540, n6541_1, n6542,
    n6543, n6544, n6545, n6546_1, n6547, n6548, n6549, n6550, n6551_1,
    n6552, n6553, n6554, n6555_1, n6556, n6557, n6558, n6559, n6560_1,
    n6561, n6562, n6563, n6564, n6565_1, n6566, n6567, n6568, n6569,
    n6570_1, n6571, n6572, n6573, n6574, n6575_1, n6576, n6577, n6578,
    n6579, n6580_1, n6581, n6582, n6583, n6584, n6585_1, n6586, n6587,
    n6588, n6589, n6590_1, n6591, n6592, n6593, n6594, n6595_1, n6596,
    n6597, n6598, n6599, n6600_1, n6601, n6602, n6603, n6604, n6605_1,
    n6606, n6607, n6608, n6609, n6610_1, n6611, n6612, n6613, n6614,
    n6615_1, n6616, n6617, n6618, n6619, n6620_1, n6621, n6622, n6623,
    n6624_1, n6625, n6626, n6627, n6628, n6629_1, n6630, n6631, n6632,
    n6633, n6634_1, n6635, n6636, n6637, n6638_1, n6639, n6640, n6641,
    n6642_1, n6643, n6644, n6645, n6646_1, n6647, n6648, n6649, n6650,
    n6651_1, n6652, n6653, n6654, n6655, n6656_1, n6657, n6658, n6659,
    n6660, n6661_1, n6662, n6663, n6664, n6665_1, n6666, n6667, n6668,
    n6669, n6670_1, n6671, n6672, n6673, n6674, n6675_1, n6676, n6677,
    n6678, n6679, n6680_1, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
    n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
    n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
    n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
    n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
    n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
    n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
    n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
    n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
    n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
    n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
    n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
    n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
    n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
    n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
    n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
    n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
    n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
    n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
    n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
    n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
    n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
    n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
    n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
    n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
    n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
    n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
    n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
    n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
    n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
    n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
    n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
    n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
    n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
    n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
    n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
    n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
    n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
    n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
    n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
    n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
    n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
    n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
    n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
    n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
    n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
    n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
    n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
    n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
    n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
    n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
    n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
    n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
    n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
    n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
    n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
    n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
    n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
    n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
    n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
    n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
    n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
    n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
    n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
    n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
    n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
    n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
    n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
    n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
    n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
    n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
    n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
    n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
    n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
    n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
    n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
    n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
    n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
    n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
    n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
    n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
    n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
    n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
    n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
    n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
    n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
    n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
    n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
    n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
    n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
    n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
    n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
    n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
    n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
    n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
    n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
    n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
    n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
    n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
    n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
    n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
    n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
    n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
    n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
    n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
    n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
    n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
    n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
    n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
    n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
    n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
    n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
    n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
    n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
    n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
    n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
    n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
    n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
    n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
    n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
    n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
    n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
    n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
    n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
    n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
    n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
    n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
    n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
    n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
    n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
    n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
    n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
    n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
    n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
    n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
    n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
    n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
    n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
    n8058, n8059, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
    n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
    n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
    n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
    n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
    n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
    n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
    n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
    n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
    n8149, n8150, n8151, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
    n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
    n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
    n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
    n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
    n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
    n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
    n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
    n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
    n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
    n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
    n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
    n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
    n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
    n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
    n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
    n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
    n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
    n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
    n8340, n8341, n8342, n8343, n8344, n8346, n8347, n8348, n8350, n8351,
    n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
    n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
    n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
    n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
    n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
    n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
    n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
    n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
    n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
    n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
    n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
    n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
    n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
    n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
    n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
    n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
    n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
    n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8533, n8534,
    n8535, n8540, n8541, n8542, n8543, n8544, n8546, n8548, n8550, n8552,
    n8554, n8556, n8558, n8560, n8562, n8563, n8565, n8566, n8568, n8569,
    n8571, n8572, n8574, n8576, n8577, n8579, n8580, n8582, n8584, n8586,
    n8587, n8589, n8590, n8592, n8593, n8595, n8596, n8598, n8599, n8601,
    n8602, n8604, n8605, n8607, n8608, n8610, n8614, n8616, n8618, n8620,
    n8622, n8624, n8626, n8628, n8630, n8632, n8634, n8636, n8637, n8639,
    n8641, n8642, n8644, n8645, n8647, n8648, n8649, n8650, n8651, n8652,
    n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
    n8663, n8664, n8665, n8667, n8668, n8669, n8670, n8671, n8673, n8674,
    n8676, n8678, n8680, n8681, n8683, n8685, n8686, n8688, n8690, n8691,
    n8693, n8695, n8696, n8698, n8700, n8701, n8703, n8705, n8706, n8708,
    n8710, n8711, n8713, n8715, n8716, n8718, n8720, n8722, n8723, n8724,
    n8726, n8728, n8730, n8732, n8734, n8736, n8738, n8740, n8742, n8744,
    n8745, n8747, n8748, n8750, n8752, n8754, n8756, n8758, n8760, n8761,
    n8762, n8764, n8766, n8768, n8770, n8771, n8772, n8774, n8776, n8778,
    n8779, n8780, n8782, n8784, n8786, n8788, n8790, n8792, n8794, n8796,
    n8798, n8800, n8802, n8804, n8806, n8808, n8810, n8812, n8814, n8816,
    n8818, n8820, n8822, n8824, n8826, n8828, n8830, n8832, n8834, n8836,
    n8838, n8839, n8841, n8842, n8844, n8845, n8847, n8849, n8851, n8853,
    n8855, n8857, n8859, n8861, n8863, n8864, n8866, n8867, n8869, n8871,
    n8873, n8874, n8876, n8877, n8879, n8881, n8883, n8884, n8886, n8887,
    n8889, n8891, n8893, n8894, n8896, n8897, n8899, n8901, n8903, n8904,
    n8906, n8907, n8909, n8910, n8912, n8914, n8915, n8917, n8919, n8920,
    n8922, n8923, n8925, n8927, n8929, n8930, n8932, n8933, n8935, n8937,
    n8939, n8940, n8942, n8943, n8945, n8947, n8949, n8950, n8952, n8954,
    n8956, n8957, n8959, n8961, n8962, n8964, n8966, n8968, n8970, n8972,
    n8974, n8976, n8978, n8980, n8982, n8984, n8986, n8988, n8990, n8992,
    n8994, n8996, n8998, n9000, n9002, n9004, n9006, n9008, n9010, n9012,
    n9014, n9016, n9018, n9020, n9022, n9024, n9026, n9028, n9030, n9032,
    n9034, n9036, n9038, n9040, n9042, n9044, n9046, n9048, n9050, n9052,
    n9054, n9056, n9058, n9060, n9062, n9064, n9066, n9068, n9070, n9071,
    n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
    n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
    n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
    n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
    n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
    n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
    n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
    n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
    n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
    n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
    n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
    n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
    n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
    n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
    n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
    n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
    n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
    n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
    n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
    n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
    n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
    n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
    n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
    n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
    n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
    n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
    n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
    n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
    n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
    n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
    n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
    n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
    n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
    n9402, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
    n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
    n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
    n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
    n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
    n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n687,
    n692_1, n697_1, n702_1, n707_1, n712, n716, n721_1, n726_1, n731_1,
    n736_1, n741_1, n746_1, n751_1, n756_1, n761_1, n766_1, n771_1, n776_1,
    n780_1, n785_1, n790_1, n795_1, n800_1, n805_1, n810_1, n815_1, n820_1,
    n823_1, n828_1, n833_1, n837_1, n841_1, n846_1, n851_1, n856_1, n861_1,
    n866_1, n871_1, n876_1, n881_1, n886_1, n890_1, n895_1, n900_1, n905_1,
    n910_1, n914_1, n919_1, n924_1, n929, n934_1, n939_1, n944_1, n948_1,
    n953_1, n958_1, n963_1, n968_1, n973_1, n978_1, n983_1, n988_1, n993_1,
    n998_1, n1003_1, n1008_1, n1013_1, n1018_1, n1022_1, n1026_1, n1031_1,
    n1036_1, n1041_1, n1045_1, n1049_1, n1054_1, n1059_1, n1064_1, n1068_1,
    n1072_1, n1077_1, n1082, n1087_1, n1092_1, n1097_1, n1102, n1107_1,
    n1112_1, n1117, n1122_1, n1127, n1132_1, n1136_1, n1140_1, n1145_1,
    n1150_1, n1155_1, n1160_1, n1165_1, n1170_1, n1174, n1177, n1181,
    n1186, n1191_1, n1196_1, n1201_1, n1205_1, n1209_1, n1214, n1219_1,
    n1224_1, n1228_1, n1232_1, n1237_1, n1242_1, n1247, n1252, n1257_1,
    n1262, n1267_1, n1272_1, n1277_1, n1282_1, n1287_1, n1292_1, n1297_1,
    n1302, n1307_1, n1312_1, n1317_1, n1322_1, n1327_1, n1331_1, n1335_1,
    n1339_1, n1344, n1349_1, n1354_1, n1358_1, n1362_1, n1367, n1372_1,
    n1377_1, n1382_1, n1387_1, n1392_1, n1397_1, n1402_1, n1407_1, n1411_1,
    n1415_1, n1420, n1423, n1428_1, n1433_1, n1438_1, n1442, n1447,
    n1452_1, n1457, n1462_1, n1467, n1472_1, n1477, n1481, n1485_1, n1490,
    n1495_1, n1500, n1504, n1509, n1513, n1517, n1522_1, n1527, n1532_1,
    n1537_1, n1542_1, n1547_1, n1552_1, n1557_1, n1562_1, n1567, n1572_1,
    n1577_1, n1581, n1586, n1591_1, n1596_1, n1601_1, n1606_1, n1611_1,
    n1616, n1621_1, n1626_1, n1631_1, n1636_1, n1641_1, n1646_1, n1650,
    n1654, n1659, n1664_1, n1669_1, n1674, n1679_1, n1684_1, n1689_1,
    n1694_1, n1699_1, n1704_1, n1709_1, n1714, n1717_1, n1722_1, n1727_1,
    n1732_1, n1737_1, n1742_1, n1747_1, n1752, n1757_1, n1762_1, n1767_1,
    n1772, n1777, n1782_1, n1787_1, n1792, n1797, n1802, n1807_1, n1812_1,
    n1816_1, n1821_1, n1826_1, n1831_1, n1836_1, n1840, n1844_1, n1849_1,
    n1854, n1859_1, n1864_1, n1868, n1873_1, n1878_1, n1883_1, n1888_1,
    n1893_1, n1898_1, n1903_1, n1908_1, n1912_1, n1916_1, n1920_1, n1925_1,
    n1930_1, n1935_1, n1940_1, n1945_1, n1950_1, n1955, n1959, n1964,
    n1969_1, n1974_1, n1979_1, n1983_1, n1988, n1993_1, n1998_1, n2002_1,
    n2007_1, n2012_1, n2017_1, n2022_1, n2027_1, n2031, n2035, n2040,
    n2045, n2050, n2055_1, n2060, n2065_1, n2070, n2074, n2078_1, n2083,
    n2087, n2092, n2096_1, n2101_1, n2106_1, n2111, n2116, n2120_1, n2124,
    n2127_1, n2131_1, n2136, n2141_1, n2146, n2150, n2154, n2159_1,
    n2164_1, n2169_1, n2173_1, n2178, n2183_1, n2188_1, n2193, n2198,
    n2203_1, n2208_1, n2212, n2217_1, n2222, n2227, n2232_1, n2237_1,
    n2242_1, n2247, n2252, n2257, n2261_1, n2265, n2270_1, n2275, n2280_1,
    n2285_1, n2289_1, n2293_1, n2297_1, n2301_1, n2306, n2309_1, n2313,
    n2318_1, n2323_1, n2328_1, n2331_1, n2336_1, n2341_1, n2345_1, n2349_1,
    n2354_1, n2359_1, n2364_1, n2369_1, n2374_1, n2379_1, n2384_1, n2388_1,
    n2393_1, n2398_1, n2403_1, n2408_1, n2413, n2418, n2423, n2428_1,
    n2432, n2436_1, n2441_1, n2445, n2449_1, n2454_1, n2458, n2463_1,
    n2468_1, n2473_1, n2478_1, n2483, n2488_1, n2493, n2498_1, n2502,
    n2506, n2511_1, n2516, n2521_1, n2525, n2530, n2535_1, n2540, n2545_1,
    n2550_1, n2555_1, n2560_1, n2565_1, n2570, n2575, n2580_1, n2585_1,
    n2590_1, n2595_1, n2600_1, n2605_1, n2610_1, n2615_1, n2619_1, n2624_1,
    n2629_1, n2634_1, n2639_1, n2644_1, n2649_1, n2654, n2659_1, n2663,
    n2668_1, n2672_1, n2677_1, n2682_1, n2687_1, n2692_1, n2697, n2701_1,
    n2705_1, n2710_1, n2715_1, n2720_1, n2725_1, n2729_1, n2733_1, n2738_1,
    n2743, n2748_1, n2752_1, n2755_1, n2760_1, n2765_1, n2770, n2774_1,
    n2778_1, n2783_1, n2788_1, n2793_1, n2798_1, n2803_1, n2808_1, n2813_1,
    n2818_1, n2823_1, n2828, n2833_1, n2838_1, n2843_1, n2848_1, n2852_1,
    n2857_1, n2862_1, n2867_1, n2872_1, n2876_1, n2881_1, n2885_1, n2890_1,
    n2895_1, n2899_1, n2904_1, n2909_1, n2914_1, n2919_1, n2924_1, n2929_1,
    n2934_1, n2937_1, n2941_1, n2946_1, n2951_1, n2956_1, n2961_1, n2966_1,
    n2971_1, n2975_1, n2979_1, n2984_1, n2989_1, n2994_1, n2999_1, n3004_1,
    n3009_1, n3013_1, n3018_1, n3023_1, n3028_1, n3033_1, n3038_1, n3042_1,
    n3047, n3052, n3057, n3061, n3065_1, n3070, n3075, n3079, n3082,
    n3086_1, n3091, n3096_1, n3101_1, n3106, n3111, n3116_1, n3121, n3126,
    n3131_1, n3136, n3141_1, n3146, n3151_1, n3156_1, n3161, n3165,
    n3170_1, n3175_1, n3180_1, n3185_1, n3190, n3195, n3200, n3205,
    n3210_1, n3215, n3219_1, n3223_1, n3228, n3232_1, n3237, n3242_1,
    n3247_1, n3252, n3257_1, n3262_1, n3267, n3270, n3275_1, n3279_1,
    n3282_1, n3286_1, n3291_1, n3296_1, n3301, n3306_1, n3311, n3316_1,
    n3321, n3326_1, n3331_1, n3336, n3340_1, n3345, n3350_1, n3355_1,
    n3360, n3365_1, n3370_1, n3375, n3379, n3382_1, n3386_1, n3391_1,
    n3396_1, n3401_1, n3406_1, n3411, n3416, n3421_1, n3426_1, n3431_1,
    n3435_1, n3439, n3444_1, n3449, n3454, n3459_1, n3464_1, n3468_1,
    n3471, n3476_1, n3480_1, n3485_1, n3490, n3495_1, n3500_1, n3505,
    n3510_1, n3515, n3519_1, n3524, n3528_1, n3533, n3538, n3543, n3548,
    n3553, n3558, n3561, n3566_1, n3571_1, n3576, n3581_1, n3586_1,
    n3591_1, n3595, n3599, n3604, n3608_1, n3613_1, n3618_1, n3623, n3627,
    n3631, n3636_1, n3641, n3646_1, n3651_1, n3656_1, n3661, n3665_1,
    n3670_1, n3675, n3680_1, n3685_1, n3690_1, n3695, n3700, n3705,
    n3710_1, n3715_1, n3720_1, n3725, n3730, n3735, n3740, n3745, n3750_1,
    n3755_1, n3760, n3765_1, n3770_1, n3775, n3779, n3783_1, n3788_1,
    n3792, n3797_1, n3802_1, n3807_1, n3812_1, n3817_1, n3822_1, n3827_1,
    n3832_1, n3837_1, n3842_1, n3847_1, n3851_1, n3856, n3861_1, n3866_1,
    n3871_1, n3876_1, n3881_1, n3886, n3891_1, n3896, n3900_1, n3903_1,
    n3907_1, n3912, n3917, n3922, n3927, n3932, n3937_1, n3942_1, n3947,
    n3952_1, n3957_1, n3962, n3967_1, n3971_1, n3975, n3980_1, n3984_1,
    n3988, n3992, n3996_1, n4001, n4006, n4010_1, n4015, n4020, n4025_1,
    n4030, n4035_1, n4039_1, n4042, n4047_1, n4052_1, n4057, n4062, n4066,
    n4070_1, n4075, n4080, n4084, n4089_1, n4094_1, n4099, n4104, n4109,
    n4114_1, n4119, n4124, n4128, n4133_1, n4138_1, n4142_1, n4147, n4151,
    n4156_1, n4160_1, n4164, n4169_1, n4174, n4178_1, n4182_1, n4187,
    n4192_1, n4197, n4202_1, n4206, n4211_1, n4216, n4221_1, n4226_1,
    n4231_1, n4235_1, n4239_1, n4244, n4249, n4254, n4259_1, n4263_1,
    n4267_1, n4272_1, n4277_1, n4282, n4287_1, n4291_1, n4296_1, n4301_1,
    n4306, n4311_1, n4316_1, n4321_1, n4326_1, n4331_1, n4336_1, n4340_1,
    n4344_1, n4349_1, n4354_1, n4359_1, n4364_1, n4369, n4374_1, n4379_1,
    n4384_1, n4389_1, n4393_1, n4397_1, n4402_1, n4407_1, n4412_1, n4417_1,
    n4422, n4427_1, n4432_1, n4437, n4442_1, n4447, n4452, n4456, n4460,
    n4465_1, n4470, n4475, n4480, n4485, n4489, n4492_1, n4495, n4499,
    n4504, n4509_1, n4514, n4519, n4524, n4529, n4534, n4539, n4544_1,
    n4549, n4554, n4559_1, n4564_1, n4569_1, n4574, n4578, n4582_1,
    n4587_1, n4592, n4597_1, n4602, n4607, n4612, n4617, n4622, n4627,
    n4631, n4636, n4640_1, n4644, n4648, n4652_1, n4657_1, n4662, n4667_1,
    n4672_1, n4677_1, n4682, n4687, n4692_1, n4697_1, n4702_1, n4707_1,
    n4712_1, n4717_1, n4722_1, n4727_1, n4731_1, n4736_1, n4741_1, n4746,
    n4751_1, n4756, n4761_1, n4766, n4770_1, n4773_1, n4777_1, n4782,
    n4787_1, n4792_1, n4797, n4802, n4807_1, n4812, n4817, n4822, n4827,
    n4832_1, n4837_1, n4842_1, n4846_1, n4851_1, n4855_1, n4859_1, n4864_1,
    n4868_1, n4873_1, n4877, n4882, n4887_1, n4890, n4894_1, n4899, n4904,
    n4909_1, n4914_1, n4919_1, n4924_1, n4929_1, n4934_1, n4939, n4944,
    n4948_1, n4953_1, n4958_1, n4963_1, n4968_1, n4973, n4978, n4983_1,
    n4987, n4992, n4997, n5002, n5007, n5011_1, n5016, n5021, n5026,
    n5031_1, n5036, n5041, n5046_1, n5051_1, n5056_1, n5060, n5064, n5069,
    n5074_1, n5079_1, n5083_1, n5088_1, n5093_1, n5098, n5103, n5107,
    n5111, n5116, n5121, n5126, n5131, n5136_1, n5141, n5146, n5151_1,
    n5156, n5160_1, n5165_1, n5170_1, n5175_1, n5180_1, n5185_1, n5190_1,
    n5195_1, n5200_1, n5205_1, n5210_1, n5214_1, n5218_1, n5223_1, n5228_1,
    n5233_1, n5237_1, n5241_1, n5246_1, n5251, n5256_1, n5261, n5265_1,
    n5269_1, n5273, n5278_1, n5283_1, n5288_1, n5293_1, n5298, n5303_1,
    n5308_1, n5313_1, n5318, n5322, n5326_1, n5331_1, n5335_1, n5339_1,
    n5344_1, n5349, n5353_1, n5356_1, n5361_1, n5366_1, n5371_1, n5376_1,
    n5381_1, n5385_1, n5389_1, n5393_1, n5398_1, n5402_1, n5406_1, n5411_1,
    n5416, n5421_1, n5426_1, n5431_1, n5436, n5441_1, n5446_1, n5451_1,
    n5456_1, n5461, n5466_1, n5471_1, n5476_1, n5481_1, n5486_1, n5491_1,
    n5496_1, n5501_1, n5506_1, n5511_1, n5516_1, n5521_1, n5526_1, n5531_1,
    n5536_1, n5541_1, n5545_1, n5549_1, n5554_1, n5558_1, n5563_1, n5568_1,
    n5573_1, n5578_1, n5583_1, n5588_1, n5593_1, n5598, n5603_1, n5608_1,
    n5613_1, n5618_1, n5623_1, n5628, n5633, n5638, n5643_1, n5648_1,
    n5653, n5658_1, n5662, n5666_1, n5671, n5676_1, n5681_1, n5686, n5690,
    n5695, n5700_1, n5705_1, n5710_1, n5714, n5718, n5723_1, n5728,
    n5733_1, n5738_1, n5743_1, n5748, n5753, n5758_1, n5763, n5768, n5772,
    n5776, n5781_1, n5786, n5791, n5796, n5801, n5806, n5811, n5816_1,
    n5821_1, n5825_1, n5828_1, n5833_1, n5838_1, n5842_1, n5846, n5850_1,
    n5855_1, n5859, n5864, n5869, n5874, n5879_1, n5884, n5888_1, n5893_1,
    n5898, n5903_1, n5908_1, n5913_1, n5918_1, n5923_1, n5928_1, n5933_1,
    n5937, n5941_1, n5946_1, n5951_1, n5956, n5961_1, n5966_1, n5971_1,
    n5975_1, n5980_1, n5985_1, n5990, n5994_1, n5998, n6003_1, n6008,
    n6012, n6017, n6022_1, n6027, n6032_1, n6037_1, n6042, n6047_1,
    n6052_1, n6056, n6061, n6066_1, n6071_1, n6076_1, n6081, n6086_1,
    n6091, n6096, n6100_1, n6104, n6109_1, n6114_1, n6119_1, n6123_1,
    n6127, n6132_1, n6137, n6142, n6147, n6152, n6156, n6160, n6165, n6169,
    n6174_1, n6179, n6183, n6188_1, n6192, n6196, n6201_1, n6206, n6211,
    n6216, n6221, n6226, n6230, n6235, n6240, n6245, n6250, n6255, n6260,
    n6265, n6270, n6275, n6279, n6284, n6289, n6293, n6297, n6302, n6306_1,
    n6310, n6315, n6320, n6325_1, n6330, n6335, n6340, n6344_1, n6349,
    n6354, n6359, n6364_1, n6369, n6373, n6376, n6380, n6385, n6390, n6395,
    n6399, n6403, n6408_1, n6413, n6417, n6422, n6427, n6432, n6437, n6442,
    n6447, n6452, n6457, n6462, n6467, n6472, n6477, n6482, n6487, n6492,
    n6497, n6502, n6507, n6512, n6517, n6522, n6526, n6531, n6536, n6541,
    n6546, n6551, n6555, n6560, n6565, n6570, n6575, n6580, n6585, n6590,
    n6595, n6600, n6605, n6610, n6615, n6620, n6624, n6629, n6634, n6638,
    n6642, n6646, n6651, n6656, n6661, n6665, n6670, n6675, n6680;
  assign Pg34972 = ~n8177 | ~Ng22;
  assign n4124_1 = Ng4369 & (Ng4366 | n6090);
  assign Pg34927 = ~n5895 | ~Ng22;
  assign Pg34925 = ~n5912 | ~Ng22;
  assign Pg34923 = ~n4252 | ~Ng22;
  assign Pg34921 = ~n5892 | ~Ng22;
  assign Pg34919 = ~n5869_1 | ~Ng22;
  assign Pg34917 = ~n5669 | ~Ng22;
  assign Pg34915 = ~n5903 | ~Ng22;
  assign Pg34913 = ~n4909 | ~Ng22;
  assign n4133 = Ng890 & (Ng528 | n5931 | ~Ng479);
  assign Pg34597 = 1'b0;
  assign n4135 = ~Pg113 | ~Ng2868;
  assign n4136 = ~Pg113 | ~Ng2873;
  assign Pg34435 = ~n9417;
  assign Pg34425 = ~n5945 | ~n6265_1;
  assign Pg34383 = ~n6264 | n5901 | ~n5930;
  assign Pg34240 = 1'b0;
  assign Pg34239 = 1'b0;
  assign Pg34238 = 1'b0;
  assign Pg34237 = 1'b0;
  assign Pg34236 = 1'b0;
  assign Pg34235 = 1'b0;
  assign Pg34234 = 1'b0;
  assign Pg34233 = 1'b0;
  assign Pg34232 = 1'b0;
  assign Pg34221 = ~n5929 | ~n6265_1;
  assign Pg34201 = ~n6264 | n5938 | ~n6122;
  assign n4151_1 = Ng4646 & (n5875 | n5915);
  assign Pg33950 = 1'b0;
  assign Pg33949 = 1'b0;
  assign Pg33948 = 1'b0;
  assign Pg33947 = 1'b0;
  assign Pg33946 = 1'b0;
  assign Pg33945 = 1'b0;
  assign Pg33935 = ~n5936;
  assign Pg33874 = ~Ng4507 | \[4507]  | n5924;
  assign Pg33659 = ~n9418 | n5947 | ~n6264;
  assign Pg33636 = ~n5950;
  assign n4162 = Pg17291 & (~Ng1171 | n5914);
  assign Pg33435 = (n9185 & (~Ng2729 | n9186)) | (Ng2729 & n9186);
  assign Pg33079 = (n9183 & (~Ng2729 | n9184)) | (Ng2729 & n9184);
  assign Pg32975 = ~n7527;
  assign Pg32454 = 1'b0;
  assign Pg32429 = 1'b0;
  assign Pg32185 = n6847 & n6844 & n6845 & n6846;
  assign Pg31863 = ~n8207;
  assign Pg31862 = ~n8080;
  assign Pg31860 = ~n8192;
  assign Pg31793 = ~n4220;
  assign Pg31521 = ~n9417;
  assign Pg30331 = ~Ng2831;
  assign Pg30330 = ~Ng2834;
  assign Pg30329 = ~\[4426] ;
  assign Pg30327 = ~Ng37;
  assign Pg28042 = n4218 | n4219;
  assign Pg28041 = n4217 | ~n8478;
  assign Pg28030 = n4215 | n4216_1;
  assign Pg26877 = ~n4214;
  assign Pg26876 = ~n4211;
  assign Pg26875 = ~n4208;
  assign Pg26801 = ~n7527;
  assign Pg25590 = 1'b0;
  assign Pg25589 = 1'b0;
  assign Pg25588 = 1'b0;
  assign Pg25587 = 1'b0;
  assign Pg25586 = 1'b0;
  assign Pg25585 = 1'b0;
  assign Pg25584 = 1'b0;
  assign Pg25583 = 1'b0;
  assign Pg25582 = 1'b0;
  assign Pg25259 = ~n8080;
  assign Pg25167 = ~n8207;
  assign Pg25114 = ~n8192;
  assign Pg24151 = 1'b0;
  assign Pg23759 = ~Ng2831;
  assign Pg23652 = ~Ng2834;
  assign Pg23612 = ~\[4426] ;
  assign Pg23190 = ~Ng25 & ~Ng22;
  assign Pg23002 = ~Ng37;
  assign Pg21727 = ~Pg35 & Ng3003;
  assign Pg12833 = ~Pg5;
  assign n4205 = ~Pg35 | n8382;
  assign n4206_1 = Ng1830 | Ng2098 | Ng1696 | Ng1964;
  assign n4207 = n6127_1 & Pg35;
  assign n4208 = n4206_1 & n4207;
  assign n4209 = Ng1710 | Ng1858 | Ng1844 | Ng2126 | Ng1724 | Ng2112 | Ng1992 | Ng1978;
  assign n4210 = n5989 & Pg35;
  assign n4211 = n4209 & n4210;
  assign n4212 = Ng1913 | Ng2047 | Ng1932 | Ng1798 | Ng1664 | Ng1779 | Ng1644 | Ng2066;
  assign n4213 = n5988 & Pg35;
  assign n4214 = n4212 & n4213;
  assign n4215 = n7837 & ~n8125 & (~n5906 | ~n8212);
  assign n4216_1 = ~n5906 & (~n5902 | ~n5905) & n7838;
  assign n4217 = ~Pg35 | n6128;
  assign n4218 = ~Pg35 | Ng962;
  assign n4219 = ~Pg35 | Ng1306;
  assign n4220 = n6888 & (n6889 | n6890 | ~n9117);
  assign n4221 = n6702 & n6703 & (Pg35 | ~Ng5052);
  assign n687 = ~n4221;
  assign n4223 = n6247 & (n6241 | n6246 | n6238);
  assign n692_1 = ~n4223;
  assign n4225 = n6439 & n6440 & (~n6006 | n6441);
  assign n697_1 = ~n4225;
  assign n4227 = n6374 & (Pg35 | ~Ng2380);
  assign n702_1 = ~n4227;
  assign n4229 = n7300 & n7301 & (n4205 | n7302);
  assign n721_1 = ~n4229;
  assign n4231 = n7273 & n7274 & (n4205 | n7275);
  assign n731_1 = ~n4231;
  assign n4233 = n7141 & n7142 & (n4205 | n7143);
  assign n736_1 = ~n4233;
  assign n4235 = n6172 & (Pg35 | ~Ng2984);
  assign n746_1 = ~n4235;
  assign n4237 = n6460 & n6461 & (~n5998_1 | n6462_1);
  assign n751_1 = ~n4237;
  assign n4239 = n7041 & n7042 & (n4205 | n7043);
  assign n756_1 = ~n4239;
  assign n4241 = (n6452_1 | ~Ng1802) & (n6616 | ~Ng1772);
  assign n761_1 = ~n4241;
  assign n4243 = n7229 & n7230 & (n4205 | n6723);
  assign n766_1 = ~n4243;
  assign n4245 = (~Ng6215 | n6667) & (~Ng6219 | n6668);
  assign n771_1 = ~n4245;
  assign n4247 = n6098 & n6099 & (Ng807 | n6093);
  assign n776_1 = ~n4247;
  assign n4249_1 = Ng1061 ^ n8020;
  assign n790_1 = n4249_1 | ~n9152;
  assign n4251 = Ng4172 | Ng4153;
  assign n4252 = n6024 & n6021 & n6022 & n6023;
  assign n795_1 = n4251 & Pg35;
  assign n4254_1 = (n6726 | n6732) & (Pg35 | ~Ng3506);
  assign n805_1 = ~n4254_1;
  assign n4256 = n6874 & n6875 & (Ng749 | n6876);
  assign n810_1 = ~n4256;
  assign n4258 = (~Pg17739 & (~Pg14738 | Pg12350)) | (Pg14738 & Pg12350);
  assign n820_1 = n4258 & ~Pg13068 & ~Pg17607 & Pg35 & ~Pg17646;
  assign n4260 = n6483 & n6484 & (~n6010 | n6485);
  assign n828_1 = ~n4260;
  assign n4262 = n6623 & n6624_1 & (~n8312 | ~Ng1714);
  assign n833_1 = ~n4262;
  assign n841_1 = ~n6738 & ~Ng3155;
  assign n4265 = n7692 & n7693 & (~Ng2165 | ~n8424);
  assign n846_1 = ~n4265;
  assign n4267 = ~Ng3689 | n8508;
  assign n856_1 = Ng3694 & (~Pg35 | n4267);
  assign n4269 = n6463 & n6464 & (~n5998_1 | n6465);
  assign n861_1 = ~n4269;
  assign n4271 = n7364 & (Pg35 | ~Ng1964);
  assign n866_1 = ~n4271;
  assign n4273 = (~Ng4621 | n6202) & (n6201 | ~Ng4639);
  assign n871_1 = ~n4273;
  assign n4275 = n7067 & n7068 & (n4205 | n7069);
  assign n876_1 = ~n4275;
  assign n4277 = n7340 & ~n9252 & (Pg35 | ~Ng2652);
  assign n881_1 = ~n4277;
  assign n4279 = (~Pg17711 & (~Pg14694 | Pg12300)) | (Pg14694 & Pg12300);
  assign n886_1 = n4279 & ~Pg13049 & ~Pg17580 & Pg35 & ~Pg17604;
  assign n4281 = n7755 & n7756 & (Ng490 | ~n8470);
  assign n890_1 = ~n4281;
  assign n4283 = n6293_1 & n6294 & (Ng772 | n6295);
  assign n900_1 = ~n4283;
  assign n4285 = n7081 & n7082 & (n4205 | n7083);
  assign n905_1 = ~n4285;
  assign n4287 = n7437 & ~n9281 & (~Ng6177 | n7438);
  assign n910_1 = ~n4287;
  assign n4289 = (n6738 | n6739) & (Pg35 | ~Ng3161);
  assign n919_1 = ~n4289;
  assign n4291 = n7061 & n7062 & (n4205 | n7063);
  assign n924_1 = ~n4291;
  assign n4293 = ~n5990_1 & n6706 & (~n6860 | ~Ng4543);
  assign n929 = ~n4293;
  assign n4295 = n7625 & (Ng3457 | n7626) & ~n9308;
  assign n934_1 = ~n4295;
  assign n4297 = n6969 & ~n9452 & (n4205 | n6970);
  assign n939_1 = ~n4297;
  assign n4299 = n6352 & n6353 & (~n6000 | n6354_1);
  assign n948_1 = ~n4299;
  assign n4301 = n6326 & (n6327 | n6328 | ~Ng4801);
  assign n953_1 = ~n4301;
  assign n4303 = n6221_1 & n6222 & (Pg35 | ~Ng4584);
  assign n958_1 = ~n4303;
  assign n4305 = ~Pg35 | ~Ng6199;
  assign n963_1 = ~n4305;
  assign n4307 = n6388 & n6389 & (~n6012_1 | n6390_1);
  assign n968_1 = ~n4307;
  assign n4309 = n7962 & n7963 & (Pg35 | ~Ng1379);
  assign n973_1 = ~n4309;
  assign n4311 = n8005 & (Pg35 | ~Ng1579);
  assign n978_1 = ~n4311;
  assign n4313 = (~Ng5176 | n6696) & (~Ng5180 | n6697);
  assign n983_1 = ~n4313;
  assign n4315 = n6179_1 & (Pg35 | ~Ng2890);
  assign n988_1 = ~n4315;
  assign n4317 = n6870 & n6871 & (Pg35 | ~Ng1018);
  assign n993_1 = ~n4317;
  assign n4319 = n7078 & n7079 & (n4205 | n7080);
  assign n998_1 = ~n4319;
  assign n4321 = n7242 & n7243 & (n4205 | n7244);
  assign n1003_1 = ~n4321;
  assign n4323 = (n8033 | ~Ng4258) & (n7997 | ~Ng4264);
  assign n1008_1 = ~n4323;
  assign n4325 = n6486 & n6487_1 & (Ng767 | n6488);
  assign n1013_1 = ~n4325;
  assign n4327 = ~Pg35 | ~Ng5853;
  assign n1018_1 = ~n4327;
  assign n4329 = n6277 & n6278 & (n6279_1 | n6276);
  assign n1031_1 = ~n4329;
  assign n4331 = ~Pg35 | ~Ng5507;
  assign n1041_1 = ~n4331;
  assign n4333 = n6966 & n6967 & (n4205 | n6968);
  assign n1049_1 = ~n4333;
  assign n4335 = n6650 & n6651_1 & (Pg35 | ~Ng291);
  assign n1054_1 = ~n4335;
  assign n4337 = n7057 & ~n9458 & (n4205 | n6682);
  assign n1059_1 = ~n4337;
  assign n4339 = ~n7985 & (Pg35 | ~Ng559);
  assign n1077_1 = ~n4339;
  assign n4341 = n6258 & (Ng608 | n6259) & ~n9441;
  assign n1082 = ~n4341;
  assign n4343 = n7213 & n7214 & (n4205 | n7215);
  assign n1092_1 = ~n4343;
  assign n4345 = n6946 & n6947 & (n4205 | n6948);
  assign n1097_1 = ~n4345;
  assign n4347 = n7003 & ~n9455 & (n4205 | n6673);
  assign n1102 = ~n4347;
  assign n4349 = (~Ng921 | n7975) & (n7974 | ~Ng904);
  assign n1107_1 = ~n4349;
  assign n4351 = ~Pg35 | ~n8251;
  assign n1127 = Ng4871 & n4351;
  assign n4353 = n7114 & n7115 & (n4205 | n7116);
  assign n1132_1 = ~n4353;
  assign n4355 = n7237 & n7238 & (n4205 | n7239);
  assign n1140_1 = ~n4355;
  assign n4357 = n6799 & n6800 & (n6795 | ~Ng1926);
  assign n1145_1 = ~n4357;
  assign n4359 = (n6668 | n6669) & (Pg35 | ~Ng6209);
  assign n1150_1 = ~n4359;
  assign n4361 = n7250 & n7251 & (n4205 | n7252);
  assign n1155_1 = ~n4361;
  assign n4363 = n6840 & n6841 & (Pg35 | ~Ng287);
  assign n1160_1 = ~n4363;
  assign n4365 = ~Pg35 | ~n8253;
  assign n1165_1 = Ng4646 & n4365;
  assign n4367 = n7261 & n7262 & (n4205 | n7263);
  assign n1170_1 = ~n4367;
  assign n4369_1 = n6609 & (n6433 | ~Ng1862);
  assign n1181 = ~n4369_1;
  assign n4371 = n7748 & n7749 & (Pg35 | ~Ng671);
  assign n1186 = ~n4371;
  assign n4373 = Ng843 ^ n8022;
  assign n1191_1 = Ng837 & (~Pg35 | n4373);
  assign n4375 = n6215 & (n6216_1 | ~Ng4322 | ~n8236);
  assign n1196_1 = ~n4375;
  assign n4377 = (Pg35 | ~Ng6395) & (n6503 | ~n9421);
  assign n1209_1 = ~n4377;
  assign n4379 = n6132 & n6133 & (Ng622 | n6134);
  assign n1214 = ~n4379;
  assign n1219_1 = ~n6728 & ~Ng3506;
  assign n4382 = n7333 & (Pg35 | ~Ng2834);
  assign n1237_1 = ~n4382;
  assign n4384 = Ng255 | Ng269 | Ng262 | ~Ng246 | ~Ng239 | ~Ng232 | ~Ng225;
  assign n4385 = Ng255 & Ng262 & Ng269 & ~Ng225 & ~Ng232 & ~Ng246 & ~Ng239;
  assign n1252 = n4384 & Pg35 & (Ng278 | n4385);
  assign n1262 = Ng4836 & n4351;
  assign n4388 = (~Ng1036 | ~n9116) & (n6642_1 | ~Ng1030);
  assign n1267_1 = ~n4388;
  assign n4390 = n7554 & n7763 & (Pg35 | ~Ng5272);
  assign n1272_1 = ~n4390;
  assign n4392 = n7303 & ~n9469 & (n4205 | n7304);
  assign n1282_1 = ~n4392;
  assign n4394 = n7434 & (n4205 | (Ng6195 & n7435));
  assign n1292_1 = ~n4394;
  assign n4396 = n7883 & n7884 & (Ng1135 | ~n8486);
  assign n1297_1 = ~n4396;
  assign n4398 = n6504 & n6505 & (n6506 | ~Ng6395);
  assign n1302 = ~n4398;
  assign n4400 = n6092 & (n6093 | ~Ng807);
  assign n1312_1 = ~n4400;
  assign n4402 = ~Pg35 | ~Ng3853;
  assign n1322_1 = ~n4402;
  assign n4404 = n6759 & n6760 & (n6755 | ~Ng2485);
  assign n1339_1 = ~n4404;
  assign n4406 = n6832 & n6833 & (Ng925 | n6834);
  assign n1344 = ~n4406;
  assign n4408 = n7099 & n7100 & (n4205 | n7101);
  assign n1354_1 = ~n4408;
  assign n4410 = n6807 & n6808 & (~Ng1798 | n6806);
  assign n1362_1 = ~n4410;
  assign n4412 = n6521 & n7806 & (Ng4076 | n7807);
  assign n1367 = ~n4412;
  assign n4414 = n7175 & n7176 & (n4205 | n6713);
  assign n1377_1 = ~n4414;
  assign n4416 = n6645 & n6646_1 & (Ng763 | n6647);
  assign n1382_1 = ~n4416;
  assign n4418 = n6987 & n6988 & (n4205 | n6989);
  assign n1387_1 = ~n4418;
  assign n4420 = n7852 & (Pg35 | ~Ng4427);
  assign n1392_1 = ~n4420;
  assign n1397_1 = Ng4864 & n4351;
  assign n4423 = n6157 & (Pg35 | ~Ng4717);
  assign n1402_1 = ~n4423;
  assign n4425 = n6838 & (Ng590 | n6839) & ~n9448;
  assign n1407_1 = ~n4425;
  assign n4427 = ~n7376 & ~n9274 & (Pg35 | ~Ng1612);
  assign n1415_1 = ~n4427;
  assign n4429 = (~Pg17674 & (~Pg14662 | Pg12238)) | (Pg14662 & Pg12238);
  assign n1420 = n4429 & ~Pg13039 & ~Pg17519 & Pg35 & ~Pg17577;
  assign n4431 = n7463 & (Ng6154 | n7464) & ~n9284;
  assign n1438_1 = ~n4431;
  assign n4433 = n7054 & n7055 & (n4205 | n7056);
  assign n1447 = ~n4433;
  assign n4435 = n6455 & n6456 & (~n5998_1 | ~n8308);
  assign n1452_1 = ~n4435;
  assign n4437_1 = n7395 & n7396 & (Ng744 | n7397);
  assign n1462_1 = ~n4437_1;
  assign n4439 = n6156_1 & (Pg35 | ~Ng4722);
  assign n1467 = ~n4439;
  assign n4441 = n6981 & n6982 & (n4205 | n6983);
  assign n1477 = ~n4441;
  assign n4443 = n6999 & (Pg35 | ~Ng5961);
  assign n1490 = ~n4443;
  assign n4445 = n8018 & n8019 & (~Pg17400 | n8014);
  assign n1500 = ~n4445;
  assign n1504 = Ng4633 & (~Pg35 | (~Ng4639 & ~n6208));
  assign n4448 = n7120 & n7121 & (n4205 | n7122);
  assign n1509 = ~n4448;
  assign n4450 = ~Pg35 | ~Ng5160;
  assign n1522_1 = ~n4450;
  assign n4452_1 = n7026 & n7027 & (n4205 | n7028);
  assign n1527 = ~n4452_1;
  assign n4454 = n6140 & n6141;
  assign n1542_1 = ~n4454;
  assign n4456_1 = ~Pg35 | ~Ng3151;
  assign n1547_1 = ~n4456_1;
  assign n4458 = (Pg35 | ~Ng3522) & (n6725 | n6726);
  assign n1562_1 = ~n4458;
  assign n4460_1 = n6521 & n6522_1 & (Ng4104 | n6523);
  assign n1567 = ~n4460_1;
  assign n4462 = n9378 ^ Pg9251;
  assign n1577_1 = n4462 & Pg35;
  assign n4464 = n6399_1 & n6400 & (~n6008_1 | ~n8287);
  assign n1581 = ~n4464;
  assign n4466 = n6576 & (n6377 | ~Ng2287);
  assign n1601_1 = ~n4466;
  assign n4468 = (~Ng4269 | n8000) & (n7999 | ~Ng4273);
  assign n1606_1 = ~n4468;
  assign n4470_1 = n7880 & ~n9437 & (Pg35 | ~Ng1384);
  assign n1611_1 = ~n4470_1;
  assign n4472 = n7467 & (Pg35 | ~Ng5831);
  assign n1621_1 = ~n4472;
  assign n4474 = n5959 & (~Ng1193 | (~Ng1171 & Ng1183));
  assign n4475_1 = Pg7916 ^ Ng1171;
  assign n1626_1 = Pg35 & (n4474 | n4475_1);
  assign n4477 = (~Ng4264 | n8032) & (n7998 | ~Ng4269);
  assign n1631_1 = ~n4477;
  assign n4479 = (n6311 | n6312) & (Pg35 | ~Ng4818);
  assign n1641_1 = ~n4479;
  assign n4481 = n7064 & n7065 & (n4205 | n7066);
  assign n1646_1 = ~n4481;
  assign n4483 = Ng4864 | Ng4878 | Ng4836 | Ng4871;
  assign n1654 = Pg35 & ~n9298 & (n4483 | ~n8760);
  assign n4485_1 = n7954 & (Pg35 | ~Ng3139);
  assign n1659 = ~n4485_1;
  assign n4487 = n7305 & ~n9470 & (n4205 | n7306);
  assign n1674 = ~n4487;
  assign n4489_1 = ~n5990_1 & ~n5993 & (~n6860 | ~Ng4540);
  assign n1679_1 = ~n4489_1;
  assign n4491 = n7264 & n7265 & (n4205 | n7266);
  assign n1684_1 = ~n4491;
  assign n4493 = n7767 & (~Pg35 | n7766 | n7768);
  assign n1694_1 = ~n4493;
  assign n4495_1 = n6152_1 & (Pg35 | ~Ng4912);
  assign n1699_1 = ~n4495_1;
  assign n4497 = n7354 & (Pg35 | ~Ng2255);
  assign n1704_1 = ~n4497;
  assign n4499_1 = n6227 & (n6228 | n6226_1 | n6229);
  assign n1709_1 = ~n4499_1;
  assign n4501 = n7858 & (~Ng4375 | (Pg35 & ~Ng4382));
  assign n1714 = ~n4501;
  assign n4503 = n6178 & (Pg35 | ~Ng2844);
  assign n1722_1 = ~n4503;
  assign n4505 = (n7758 | ~Ng417) & (n8027 | ~Ng446);
  assign n1727_1 = ~n4505;
  assign n4507 = n7044 & n7045 & (n4205 | n7046);
  assign n1747_1 = ~n4507;
  assign n4509 = n7951 & (Pg35 | ~Ng3490);
  assign n1757_1 = ~n4509;
  assign n1762_1 = ~n6687 & ~Ng5511;
  assign n4512 = (n6728 | n6729) & (Pg35 | ~Ng3512);
  assign n1767_1 = ~n4512;
  assign n4514_1 = n6467_1 & (Pg35 | ~Ng1687);
  assign n1772 = ~n4514_1;
  assign n4516 = n7495 & n7761 & (Pg35 | ~Ng5965);
  assign n1782_1 = ~n4516;
  assign n4518 = n7855 & n7856 & n7857;
  assign n1787_1 = ~n4518;
  assign n4520 = Ng518 & Ng203 & ~Ng513;
  assign n4521 = Ng182 & (Ng168 | Ng174);
  assign n4522 = Ng168 & Ng174;
  assign n1797 = Pg35 & n4520 & (n4521 | n4522);
  assign n4524_1 = n7171 & (Pg35 | ~Ng3961);
  assign n1802 = ~n4524_1;
  assign n4526 = (n7790 | ~n9147) & (n7791 | ~Ng4749);
  assign n1807_1 = ~n4526;
  assign n4528 = n6411 & (Pg35 | ~Ng2089);
  assign n1812_1 = ~n4528;
  assign n4530 = n7198 & n7199 & (n4205 | n7200);
  assign n1821_1 = ~n4530;
  assign n4532 = Ng1052 ^ n7888;
  assign n1836_1 = Pg35 & n4532 & ~Ng979;
  assign n4534_1 = n6562 & n6563 & (n6359_1 | ~Ng2465);
  assign n1849_1 = ~n4534_1;
  assign n4536 = n7050 & n7051 & (n4205 | n7052);
  assign n1854 = ~n4536;
  assign n4538 = ~n5990_1 & n6708 & (~n6860 | ~Ng4480);
  assign n1859_1 = ~n4538;
  assign n1864_1 = ~Ng358 & Pg35 & ~Pg8719;
  assign n4541 = (Pg35 | ~Ng3171) & (n6735 | n6736);
  assign n1873_1 = ~n4541;
  assign n4543 = n6620_1 & (n6452_1 | ~Ng1728);
  assign n1878_1 = ~n4543;
  assign n4545 = n6356 & (Pg35 | ~Ng2514);
  assign n1883_1 = ~n4545;
  assign n4547 = n7569 & (Pg35 | ~Ng3831);
  assign n1888_1 = ~n4547;
  assign n4549_1 = ~Pg35 | ~Ng4917;
  assign n1898_1 = ~n4549_1;
  assign n4551 = (Pg35 | ~Ng1199) & (n4474 | ~n8747);
  assign n1903_1 = ~n4551;
  assign n4553 = (n7903 | n7904) & (Pg35 | ~Ng832);
  assign n1908_1 = ~n4553;
  assign n4555 = n7392 & n7393 & (Ng914 | n7394);
  assign n1916_1 = ~n4555;
  assign n4557 = n6638_1 & ~n9361 & (Ng1008 | n7385);
  assign n4558 = ~n6638_1 | n8083;
  assign n1930_1 = Pg35 & (n4557 | (Ng969 & n4558));
  assign n4560 = n6231 & (n6228 | n6230_1 | n6232);
  assign n1935_1 = ~n4560;
  assign n4562 = n6527 & n6528 & (n6529 | ~Ng4054);
  assign n1940_1 = ~n4562;
  assign n4564 = n7922 & (Pg35 | ~Ng6187);
  assign n1945_1 = ~n4564;
  assign n1950_1 = Ng5073 & (~Pg35 | Ng5069);
  assign n4567 = (n6687 | n6688) & (Pg35 | ~Ng5517);
  assign n1955 = ~n4567;
  assign n4569 = n6910 & n6911 & (n4205 | n6912);
  assign n1964 = ~n4569;
  assign n4571 = n6469 & (n6470 | ~Ng1682);
  assign n1974_1 = ~n4571;
  assign n4573 = n7887 & ~n9473 & (Ng1105 | ~n8488);
  assign n1988 = ~n4573;
  assign n4575 = n6954 & n6955 & (n4205 | n6956);
  assign n1998_1 = ~n4575;
  assign n4577 = n7355 & ~n9261 & (Pg35 | ~Ng2250);
  assign n2012_1 = ~n4577;
  assign n4579 = n6234 & (n6228 | n6233 | n6235_1);
  assign n2017_1 = ~n4579;
  assign n4581 = n7736 & n7737 & (Ng911 | ~n8341);
  assign n2022_1 = ~n4581;
  assign n4583 = n6457_1 & n6458 & (~n5998_1 | n6459);
  assign n2035 = ~n4583;
  assign n4585 = n7058 & n7059 & (n4205 | n7060);
  assign n2040 = ~n4585;
  assign n4587 = n7267 & n7268 & (n4205 | n7269);
  assign n2045 = ~n4587;
  assign n4589 = n7928 & (Pg35 | ~Ng5495);
  assign n2050 = ~n4589;
  assign n4591 = n6167 & (Pg35 | ~Ng2950);
  assign n2055_1 = ~n4591;
  assign n4593 = n7216 & n7217 & (n4205 | n7218);
  assign n2060 = ~n4593;
  assign n4595 = n6949 & n6950 & (n4205 | n6663);
  assign n2070 = ~n4595;
  assign n4597 = n6825 & n6826 & (Pg35 | ~Ng1367);
  assign n2078_1 = ~n4597;
  assign n4599 = n6493 & n6494 & (Pg35 | ~Ng153);
  assign n2087 = ~n4599;
  assign n4601 = n6245_1 & (n6241 | n6244 | n6235_1);
  assign n2092 = ~n4601;
  assign n4603 = n7258 & n7259 & (n4205 | n7260);
  assign n2101_1 = ~n4603;
  assign n4605 = n6592 & (Pg35 | ~Ng2108);
  assign n2106_1 = ~n4605;
  assign n4607_1 = n8029 & (Pg35 | ~Ng437);
  assign n2116 = ~n4607_1;
  assign n4609 = n6835 & n6836 & (Ng758 | n6837);
  assign n2131_1 = ~n4609;
  assign n4611 = n7919 & (Pg35 | ~Ng6533);
  assign n2141_1 = ~n4611;
  assign n4613 = n7105 & n7106 & (n4205 | n7107);
  assign n2146 = ~n4613;
  assign n4615 = n7007 & ~n9456 & (n4205 | n7008);
  assign n2154 = ~n4615;
  assign n4617_1 = n6951 & n6952 & (n4205 | n6953);
  assign n2159_1 = ~n4617_1;
  assign n4619 = n6100 & n6101 & (Ng632 | n6102);
  assign n2164_1 = ~n4619;
  assign n4621 = n7222 & n7223 & (n4205 | n7224);
  assign n2173_1 = ~n4621;
  assign n4623 = n6817 & n6818 & (~Ng1664 | n6816);
  assign n2183_1 = ~n4623;
  assign n4625 = n8014 & (Pg35 | ~\[4421] );
  assign n2188_1 = ~n4625;
  assign n4627_1 = n6915 & n6916 & (n4205 | n6917);
  assign n2193 = ~n4627_1;
  assign n4629 = n7896 & (Pg35 | ~Ng269);
  assign n2198 = ~n4629;
  assign n4631_1 = ~Ng4040 | n8507;
  assign n2203_1 = Ng4045 & (~Pg35 | n4631_1);
  assign n4633 = n7847 & (~Ng4438 | (Pg35 & ~Ng4382));
  assign n2208_1 = ~n4633;
  assign n4635 = ~n6680 & (Pg35 | ~\[4437] );
  assign n2217_1 = ~n4635;
  assign n4637 = Ng4681 | Ng4688 | Ng4674 | Ng4646;
  assign n6680 = Pg35 & ~n9300 & (n4637 | ~n8761);
  assign n4639 = n6521 & n6862 & (~Pg35 | n6863);
  assign n2222 = ~n4639;
  assign n4641 = ~n5990_1 & n6710 & (~n6860 | ~Ng4495);
  assign n2227 = ~n4641;
  assign n4643 = (n6220 | n6223) & (Pg35 | ~Ng4332);
  assign n2252 = ~n4643;
  assign n4645 = n6298 & n6299 & (Pg35 | ~Ng298);
  assign n2257 = ~n4645;
  assign n4647 = n7468 & ~n9285 & (~Ng5831 | n7469);
  assign n2265 = ~n4647;
  assign n4649 = n7898 & (Pg35 | ~Ng262);
  assign n2270_1 = ~n4649;
  assign n4651 = n6830 & n6831 & (Pg35 | ~Ng1024);
  assign n2293_1 = ~n4651;
  assign n4653 = n7307 & n7308 & (n4205 | n7309);
  assign n2301_1 = ~n4653;
  assign n4655 = n6394 & (n6395_1 | ~Ng2241);
  assign n2318_1 = ~n4655;
  assign n4657 = n8003 & n8004 & (Ng1564 | ~n8495);
  assign n2323_1 = ~n4657;
  assign n4659 = n6901 & n6902 & (n4205 | n6903);
  assign n2336_1 = ~n4659;
  assign n4661 = n7902 & (Pg35 | ~Ng872);
  assign n2349_1 = ~n4661;
  assign n4663 = ~n5991 & n6710 & (~n6860 | ~Ng4501);
  assign n2359_1 = ~n4663;
  assign n4665 = (~Ng5869 | n6676) & (~Ng5873 | n6677);
  assign n2364_1 = ~n4665;
  assign n4667 = n6857 & (n6855 | ~Ng5037 | ~n8723);
  assign n2369_1 = ~n4667;
  assign n4669 = n6773 & n6769 & n6774;
  assign n2374_1 = ~n4669;
  assign n4671 = n7153 & n7154 & (n4205 | n7155);
  assign n2388_1 = ~n4671;
  assign n4673 = n7087 & n7088 & (n4205 | n7089);
  assign n2393_1 = ~n4673;
  assign n4675 = (n6677 | n6678) & (Pg35 | ~Ng5863);
  assign n2398_1 = ~n4675;
  assign n4677 = n8005 & (Pg35 | ~Ng1585);
  assign n2403_1 = ~n4677;
  assign n4679 = n6973 & n6974 & (n4205 | n6975);
  assign n2413 = ~n4679;
  assign n4681 = n7038 & n7039 & (n4205 | n7040);
  assign n2418 = ~n4681;
  assign n4683 = n7923 & n7924 & (~n8386 | ~Ng6167);
  assign n2428_1 = ~n4683;
  assign n4685 = n6551_1 & n6552 & (n6340_1 | ~Ng2599);
  assign n2436_1 = ~n4685;
  assign n4687_1 = n7876 & ~n9472 & (Ng1448 | ~n8483);
  assign n2441_1 = ~n4687_1;
  assign n4689 = n7683 & n7684 & (~Ng2299 | ~n8421);
  assign n2449_1 = ~n4689;
  assign n2454_1 = ~n6697 & ~Ng5164;
  assign n4692 = n6652 & n6653 & (Pg35 | ~Ng150);
  assign n2463_1 = ~n4692;
  assign n2468_1 = ~n6658 & ~Ng6549;
  assign n4695 = (n7565 | n7566) & (Pg35 | ~Ng4076);
  assign n2473_1 = ~n4695;
  assign n4697 = n6329 & n6330_1 & (Pg35 | ~Ng4793);
  assign n2478_1 = ~n4697;
  assign n4699 = n7180 & n7181 & (n4205 | n7182);
  assign n2488_1 = ~n4699;
  assign n4701 = n6918 & n6919 & (n4205 | n6920);
  assign n2506 = ~n4701;
  assign n4703 = n7390 & n7391 & (Pg35 | ~Ng1002);
  assign n2516 = ~n4703;
  assign n4705 = Pg35 & ((~n5425 & ~n5965) | ~n8510);
  assign n2521_1 = n4705 & ~Pg17320 & ~Pg17423 & ~Pg17404;
  assign n4707 = n7346 & ~n9256 & (Pg35 | ~Ng2441);
  assign n2535_1 = ~n4707;
  assign n4709 = n6333 & n6743 & (~Pg35 | n6744);
  assign n2540 = ~n4709;
  assign n4711 = (Pg35 | ~Ng6049) & (n6509 | ~n9423);
  assign n2545_1 = ~n4711;
  assign n4713 = n7732 & n7733 & (Ng1256 | ~n8335);
  assign n2550_1 = ~n4713;
  assign n4715 = n6852 & n6853 & (n6851 | ~Ng5016);
  assign n2555_1 = ~n4715;
  assign n4717 = n6451 & (n6452_1 | ~Ng1816);
  assign n2565_1 = ~n4717;
  assign n4719 = ~n1654 & (Pg35 | ~Ng4572);
  assign n2575 = ~n4719;
  assign n2580_1 = Pg35 & (~Ng4462 | ~n6290 | ~Ng10384);
  assign n4722 = n7570 & ~n9301 & (~Ng3831 | n7571);
  assign n2585_1 = ~n4722;
  assign n4724 = (Pg35 | ~Ng3352) & (n6538 | ~n9425);
  assign n2595_1 = ~n4724;
  assign n4726 = n6570_1 & (Pg35 | ~Ng2399);
  assign n2600_1 = ~n4726;
  assign n4728 = n6182 & (Pg35 | ~Ng2138);
  assign n2605_1 = ~n4728;
  assign n4730 = n7374 & (Pg35 | ~Ng1696);
  assign n2610_1 = ~n4730;
  assign n4732 = (n7983 | ~Ng513) & (n7987 | ~Ng504);
  assign n2615_1 = ~n4732;
  assign n4734 = (Pg35 | ~Ng5357) & (n6517_1 | ~n9422);
  assign n2624_1 = ~n4734;
  assign n4736 = n6333 & n6334 & (Ng2763 | n6335_1);
  assign n2629_1 = ~n4736;
  assign n4738 = (n6322 | n6323) & (Pg35 | ~Ng4818);
  assign n2634_1 = ~n4738;
  assign n4740 = n6144 & n6145;
  assign n2639_1 = ~n4740;
  assign n4742 = n6868 & n6869 & (Ng1263 | ~n8336);
  assign n2644_1 = ~n4742;
  assign n4744 = n6432_1 & (n6433 | ~Ng1950);
  assign n2649_1 = ~n4744;
  assign n4746_1 = n7529 & ~n9293 & (~Ng5138 | n7530);
  assign n2654 = ~n4746_1;
  assign n4748 = n6382 & n6383 & (~n6012_1 | n6384);
  assign n2659_1 = ~n4748;
  assign n4750 = (n6197 | n6198) & (Pg35 | ~Ng4659);
  assign n2672_1 = ~n4750;
  assign n4752 = n6777 & n6778 & (~Ng2223 | n6776);
  assign n2677_1 = ~n4752;
  assign n4754 = n7494 & (Ng5808 | n7495) & ~n9288;
  assign n2682_1 = ~n4754;
  assign n4756_1 = n6904 & n6905 & (n4205 | n6906);
  assign n2687_1 = ~n4756_1;
  assign n4758 = n6420 & n6421 & (~n6004 | n6422_1);
  assign n2692_1 = ~n4758;
  assign n4760 = (~Ng3869 | n6717) & (~Ng3873 | n6718);
  assign n2697 = ~n4760;
  assign n4762 = n6378 & ~n9444 & (~n6012_1 | n6379);
  assign n2705_1 = ~n4762;
  assign n4764 = n7864 & (Pg35 | ~Ng2799);
  assign n2710_1 = ~n4764;
  assign n4766_1 = n7009 & n7010 & (n4205 | n7011);
  assign n2715_1 = ~n4766_1;
  assign n4768 = n6589 & ~n9432 & (~Ng2047 | n6588);
  assign n2720_1 = ~n4768;
  assign n4770 = (n6718 | n6719) & (Pg35 | ~Ng3863);
  assign n2725_1 = ~n4770;
  assign n4772 = n7090 & n7091 & (n4205 | n7092);
  assign n2733_1 = ~n4772;
  assign n4774 = n7210 & n7211 & (n4205 | n7212);
  assign n2748_1 = ~n4774;
  assign n4776 = (~Pg35 | ~Ng4411) & (n7854 | ~Ng4401);
  assign n2760_1 = ~n4776;
  assign n4778 = n6976 & ~n9454 & (n4205 | n6977);
  assign n2765_1 = ~n4778;
  assign n4780 = n6945 & (Pg35 | ~Ng6307);
  assign n2770 = ~n4780;
  assign n4782_1 = n7970 & n7971 & (Pg35 | ~Ng1036);
  assign n2778_1 = ~n4782_1;
  assign n4784 = n7341 & ~n9253 & (Pg35 | ~Ng2575);
  assign n2783_1 = ~n4784;
  assign n4786 = n6559 & (Pg35 | ~Ng2533);
  assign n2788_1 = ~n4786;
  assign n4788 = (~Pg35 | ~Ng4443) & (n7845 | ~Ng4434);
  assign n2798_1 = ~n4788;
  assign n4790 = n7464 & n7760 & (Pg35 | ~Ng6311);
  assign n2808_1 = ~n4790;
  assign n4792 = n6993 & n6994 & (n4205 | n6995);
  assign n2813_1 = ~n4792;
  assign n4794 = n7900 & (Pg35 | ~Ng255);
  assign n2818_1 = ~n4794;
  assign n4796 = n7117 & n7118 & (n4205 | n7119);
  assign n2823_1 = ~n4796;
  assign n4798 = ~Pg35 | ~Ng6545;
  assign n2828 = ~n4798;
  assign n4800 = n7347 & ~n9257 & (~Ng2417 | n7348);
  assign n2833_1 = ~n4800;
  assign n4802_1 = n6617 & n6618 & (n6452_1 | ~Ng1772);
  assign n2838_1 = ~n4802_1;
  assign n4804 = n6849 & ~n9233 & (Pg35 | ~Ng5046);
  assign n2843_1 = ~n4804;
  assign n4806 = n6434 & n6435 & (~n6006 | n6436);
  assign n2852_1 = ~n4806;
  assign n4808 = (n6340_1 | ~Ng2629) & (n6550 | ~Ng2599);
  assign n2857_1 = ~n4808;
  assign n4810 = n7829 & n7830 & (Ng572 | n7831);
  assign n2862_1 = ~n4810;
  assign n4812_1 = ~Pg35 | ~Ng2130;
  assign n2867_1 = ~n4812_1;
  assign n4814 = n6521 & n6711 & (Ng4108 | n6712);
  assign n2872_1 = ~n4814;
  assign n4816 = n8028 & (Pg35 | ~Ng424);
  assign n2881_1 = ~n4816;
  assign n4818 = ~n3847_1 & (Pg35 | ~Ng753);
  assign n2895_1 = ~n4818;
  assign n4820 = (Pg35 | ~Ng4054) & (n6526_1 | ~n9419);
  assign n2899_1 = ~n4820;
  assign n4822_1 = (Pg35 | ~Ng5873) & (n6674 | n6675_1);
  assign n2904_1 = ~n4822_1;
  assign n4824 = n7362 & ~n9266 & (~Ng1992 | n7363);
  assign n2909_1 = ~n4824;
  assign n4826 = (~Ng3167 | n6737) & (~Ng3171 | n6738);
  assign n2914_1 = ~n4826;
  assign n4828 = (Pg35 | ~Ng843) & (~Ng837 | ~n8838);
  assign n2919_1 = ~n4828;
  assign n4830 = (~n7739 | ~n9149) & (n7977 | ~Ng817);
  assign n2924_1 = ~n4830;
  assign n4832 = n7004 & n7005 & (n4205 | n7006);
  assign n2929_1 = ~n4832;
  assign n4834 = n7916 & (n7915 | (n7917 & ~Ng26885));
  assign n2951_1 = ~n4834;
  assign n4836 = n7863 & (Pg35 | ~Ng2811);
  assign n2961_1 = ~n4836;
  assign n4838 = n7626 & n7809 & (Pg35 | ~Ng3614);
  assign n2966_1 = ~n4838;
  assign n4840 = (Pg35 | ~Ng3703) & (n6532 | ~n9424);
  assign n2971_1 = ~n4840;
  assign n4842 = n7897 & (Pg35 | ~Ng239);
  assign n2989_1 = ~n4842;
  assign n4844 = n7596 & (Ng3808 | n7597) & ~n9304;
  assign n3013_1 = ~n4844;
  assign n4846 = Ng10384 & Ng4473;
  assign n3018_1 = Ng4462 | ~n6290 | ~Pg35 | n4846;
  assign n4848 = n7183 & n7184 & (n4205 | n7185);
  assign n3023_1 = ~n4848;
  assign n4850 = n7169 & n7170 & (Pg35 | ~Ng4087);
  assign n3028_1 = ~n4850;
  assign n4852 = n6813 & n6809 & n6814;
  assign n3033_1 = ~n4852;
  assign n4854 = (~Pg17760 & (~Pg14779 | Pg12422)) | (Pg14779 & Pg12422);
  assign n3038_1 = n4854 & ~Pg13085 & ~Pg17649 & Pg35 & ~Pg17685;
  assign n4856 = n6301 & n6302_1 & (Pg35 | ~Ng157);
  assign n3042_1 = ~n4856;
  assign n4858 = n7598 & (n4205 | (Ng3498 & n7599));
  assign n3052 = ~n4858;
  assign n4860 = n7752 & n7753 & (Ng586 | n7754);
  assign n3057 = ~n4860;
  assign n4862 = n6749 & n6750 & (n6745 | ~Ng2619);
  assign n3065_1 = ~n4862;
  assign n4864 = n7388 & (Ng1183 | n7389);
  assign n3070 = ~n4864;
  assign n4866 = n6480 & n6481 & (~n6010 | n6482_1);
  assign n3075 = ~n4866;
  assign n4868 = n6611 & ~n9434 & (~Ng1779 | n6610_1);
  assign n3086_1 = ~n4868;
  assign n4870 = ~n7660 & (~Pg35 | n7658 | ~Ng2652);
  assign n3091 = ~n4870;
  assign n4872 = n7356 & ~n9262 & (Pg35 | ~Ng2173);
  assign n3096_1 = ~n4872;
  assign n4874 = n7349 & (Pg35 | ~Ng2389);
  assign n3101_1 = ~n4874;
  assign n4876 = n7772 & (~Pg35 | n7771 | n7773);
  assign n3111 = ~n4876;
  assign n4878 = (Pg35 | ~Ng5527) & (n6684 | n6685);
  assign n3116_1 = ~n4878;
  assign n4880 = n7333 & (Pg35 | ~Ng2803);
  assign n3121 = ~n4880;
  assign n4882_1 = n7380 & n7381 & (Pg35 | ~Ng1345);
  assign n3126 = ~n4882_1;
  assign n4884 = n6996 & n6997 & (n4205 | n6998);
  assign n3131_1 = ~n4884;
  assign n4886 = Ng1146 & (~n4887 | ~Ng1152);
  assign n4887 = ~Ng1183 & Pg13259 & ~Ng1171;
  assign n3136 = Pg35 & (n4886 | (n4887 & ~Ng1099));
  assign n4889 = n6747 & n6748 & (~Ng2625 | n6746);
  assign n3141_1 = ~n4889;
  assign n4891 = n6842 & n6843 & (Pg35 | ~Ng164);
  assign n3146 = ~n4891;
  assign n4893 = n7375 & ~n9273 & (Pg35 | ~Ng1691);
  assign n3151_1 = ~n4893;
  assign n4895 = (n6656_1 | n6662) & (Pg35 | ~Ng6549);
  assign n3156_1 = ~n4895;
  assign n3161 = \[4431]  & Pg35;
  assign n4898 = (Pg35 | ~Ng3873) & (n6715 | n6716);
  assign n3165 = ~n4898;
  assign n4900 = n6921 & n6922 & (n4205 | n6923);
  assign n3170_1 = ~n4900;
  assign n4902 = n7952 & n7953 & (~n8405 | ~Ng3470);
  assign n3175_1 = ~n4902;
  assign n4904_1 = n7177 & n7178 & (n4205 | n7179);
  assign n3180_1 = ~n4904_1;
  assign n4906 = (n7983 | ~Ng518) & (n7987 | ~Ng513);
  assign n3185_1 = ~n4906;
  assign n4908 = Ng538 | Ng209;
  assign n4909 = n6068 & n6065 & n6066 & n6067;
  assign n3190 = n4908 & Pg35;
  assign n4911 = n6545 & ~n9428 & (~Ng2606 | n6544);
  assign n3195 = ~n4911;
  assign n4913 = n7874 & n7875 & (Ng1472 | ~n8482);
  assign n3200 = ~n4913;
  assign n4915 = (n7743 | n8026) & (Pg35 | ~Ng546);
  assign n3205 = ~n4915;
  assign n4917 = (Pg35 | ~Ng5180) & (n6694 | n6695);
  assign n3210_1 = ~n4917;
  assign n4919 = n7150 & n7151 & (n4205 | n7152);
  assign n3228 = ~n4919;
  assign n4921 = n6195 & (n6196_1 | ~Ng4664 | ~n8230);
  assign n3237 = ~n4921;
  assign n4923 = n8014 & (Pg35 | ~Ng1236);
  assign n3242_1 = ~n4923;
  assign n4925 = (Pg35 | ~\[4507] ) & (n7994 | n7995);
  assign n3247_1 = ~n4925;
  assign n4927 = n6177 & (Pg35 | ~Ng2852);
  assign n3252 = ~n4927;
  assign n4929 = n6285 & n6286 & (n6287 | n6284_1);
  assign n3257_1 = ~n4929;
  assign n4931 = n6936 & n6937 & (n4205 | n6938);
  assign n3262_1 = ~n4931;
  assign n4933 = (Pg35 | ~Ng1542) & (n5559 | ~n8744);
  assign n3275_1 = ~n4933;
  assign n4935 = n6907 & n6908 & (n4205 | n6909);
  assign n3286_1 = ~n4935;
  assign n4937 = (n6433 | ~Ng1936) & (n6605_1 | ~Ng1906);
  assign n3291_1 = ~n4937;
  assign n4939_1 = n7988 & (n7986 | n7755);
  assign n3301 = ~n4939_1;
  assign n4941 = n6753 & n6749 & n6754;
  assign n3306_1 = ~n4941;
  assign n4943 = n6710 & n6861 & (Pg35 | ~Ng4477);
  assign n3311 = ~n4943;
  assign n4945 = n6380_1 & n6381 & (~n6012_1 | ~n8279);
  assign n3316_1 = ~n4945;
  assign n4947 = n7240 & ~n9466 & (n4205 | n7241);
  assign n3321 = ~n4947;
  assign n4949 = n7093 & n7094 & (n4205 | n7095);
  assign n3326_1 = ~n4949;
  assign n4951 = n7256 & ~n9468 & (n4205 | n7257);
  assign n3331_1 = ~n4951;
  assign n4953 = n7253 & n7254 & (n4205 | n7255);
  assign n3345 = ~n4953;
  assign n4955 = n6978 & n6979 & (n4205 | n6980);
  assign n3350_1 = ~n4955;
  assign n3355_1 = Ng4681 & n4365;
  assign n4958 = n7159 & n7160 & (n4205 | n7161);
  assign n3365_1 = ~n4958;
  assign n4960 = n7310 & ~n9471 & (n4205 | n7311);
  assign n3370_1 = ~n4960;
  assign n4962 = n6418 & n6419 & (~n6004 | ~n8295);
  assign n3375 = ~n4962;
  assign n4964 = n7403 & (n4205 | (Ng6541 & n7404));
  assign n3386_1 = ~n4964;
  assign n4966 = n7283 & n7284 & (n4205 | n6733);
  assign n3391_1 = ~n4966;
  assign n4968 = n6626 & (Pg35 | ~Ng1636);
  assign n3396_1 = ~n4968;
  assign n4970 = n7788 & (~Pg35 | n7787 | n7789);
  assign n3401_1 = ~n4970;
  assign n4972 = n7899 & (Pg35 | ~Ng232);
  assign n3406_1 = ~n4972;
  assign n4974 = n7989 & (Pg35 | ~Ng168);
  assign n3421_1 = ~n4974;
  assign n4976 = (n6666 | n6672) & (Pg35 | ~Ng6203);
  assign n3426_1 = ~n4976;
  assign n4978_1 = (n7910 | n7911) & (Pg35 | ~Ng355);
  assign n3431_1 = ~n4978_1;
  assign n4980 = ~Pg35 | ~Ng3502;
  assign n3444_1 = ~n4980;
  assign n4982 = n6578 & ~n9431 & (~Ng2204 | n6577);
  assign n3449 = ~n4982;
  assign n4984 = n7125 & n7126 & (n4205 | n7127);
  assign n3454 = ~n4984;
  assign n4986 = n6217 & n6218 & (Pg35 | ~Ng4601);
  assign n3459_1 = ~n4986;
  assign n4988 = n6112 & n6113 & (Ng794 | n6114);
  assign n3464_1 = ~n4988;
  assign n4990 = n8025 & (~Ng703 | n8024);
  assign n3485_1 = ~n4990;
  assign n4992_1 = n7297 & n7298 & (n4205 | n7299);
  assign n3495_1 = ~n4992_1;
  assign n4994 = n6595_1 & n6596 & (n6414 | ~Ng2040);
  assign n3500_1 = ~n4994;
  assign n4996 = n6164 & (Pg35 | ~Ng4176);
  assign n3505 = ~n4996;
  assign n4998 = (~Ng4633 | n6207) & (~Ng4628 | n6209);
  assign n3510_1 = ~n4998;
  assign n5000 = n6159 & (Pg35 | ~Ng4727);
  assign n3519_1 = ~n5000;
  assign n5002_1 = n7470 & ~n9286 & (~n6884 | ~n8444);
  assign n3528_1 = ~n5002_1;
  assign n5004 = n6769 & n6770 & (n6765 | ~Ng2351);
  assign n3533 = ~n5004;
  assign n5006 = ~Ng6727 | ~n8502;
  assign n3543 = Ng6732 & (~Pg35 | n5006);
  assign n5008 = (n6521 | n7943) & (Pg35 | ~Ng4125);
  assign n3553 = ~n5008;
  assign n5010 = n7603 & ~n9306 & (~n8105 | ~n8453);
  assign n3566_1 = ~n5010;
  assign n5012 = n7804 & n7805 & (n7801 | ~n8473);
  assign n3571_1 = ~n5012;
  assign n5014 = n6856 & (n6855 | ~Ng5041 | ~n8379);
  assign n3576 = ~n5014;
  assign n5016_1 = ~Ng4452 & (n7844 | n7846 | ~Ng4430);
  assign n3581_1 = ~n5016_1;
  assign n5018 = n7432 & (Ng6500 | n7433) & ~n9280;
  assign n3591_1 = ~n5018;
  assign n5020 = n7629 & (Pg35 | ~Ng3129);
  assign n3599 = ~n5020;
  assign n5022 = n7810 & (Pg35 | ~Ng3263);
  assign n3604 = ~n5022;
  assign n3613_1 = Ng4674 & n4365;
  assign n5025 = n6491 & n6492_1 & (Pg35 | ~Ng294);
  assign n3618_1 = ~n5025;
  assign n5027 = n6803 & n6799 & n6804;
  assign n3631 = ~n5027;
  assign n5029 = n6165_1 & (Pg35 | ~Ng2994);
  assign n3636_1 = ~n5029;
  assign n5031 = n7276 & n7277 & (n4205 | n7278);
  assign n3641 = ~n5031;
  assign n3646_1 = Ng160 & (~Pg35 | ~n9218);
  assign n5034 = n7823 & n7824 & (Pg35 | ~Ng822);
  assign n3656_1 = ~n5034;
  assign n5036_1 = ~Ng1008 & ~Ng969 & ~n4558;
  assign n3661 = Pg35 & ~n9151 & (n5036_1 | ~n8511);
  assign n5038 = n6554 & (n6340_1 | ~Ng2555);
  assign n3665_1 = ~n5038;
  assign n5040 = n7433 & n7759 & (Pg35 | ~Ng6657);
  assign n3670_1 = ~n5040;
  assign n5042 = n7406 & ~n9277 & (~Ng6523 | n7407);
  assign n3680_1 = ~n5042;
  assign n5044 = n7378 & (Ng1526 | n7379);
  assign n3685_1 = ~n5044;
  assign n5046 = (n6219 | n6220) & (Pg35 | ~Ng4593);
  assign n3690_1 = ~n5046;
  assign n5048 = ~n5049 | Ng854;
  assign n5049 = ~Pg8719 | Ng385 | ~Ng376 | ~Ng370;
  assign n5050 = n6250_1 | ~n9329;
  assign n3695 = n5048 & Pg35 & (n5049 | n5050);
  assign n5052 = n7730 & (n7731 | ~Ng1484);
  assign n3700 = ~n5052;
  assign n5054 = n6155 & (Pg35 | ~Ng4917);
  assign n3705 = ~n5054;
  assign n3710_1 = Ng5077 & (~Pg35 | ~n8914);
  assign n5057 = (n6675_1 | n6681) & (Pg35 | ~Ng5857);
  assign n3715_1 = ~n5057;
  assign n5059 = ~n7669 & (~Pg35 | n7667 | ~Ng2518);
  assign n3725 = ~n5059;
  assign n5061 = n6337 & (Pg35 | ~Ng2648);
  assign n3730 = ~n5061;
  assign n5063 = n7907 & n7908 & (Ng568 | n7909);
  assign n3735 = ~n5063;
  assign n5065 = n7279 & (Pg35 | ~Ng3259);
  assign n3740 = ~n5065;
  assign n5067 = n6927 & n6928 & (n4205 | n6929);
  assign n3745 = ~n5067;
  assign n5069_1 = ~Ng6035 | ~n8504;
  assign n3750_1 = Ng6040 & (~Pg35 | n5069_1);
  assign n3765_1 = ~n6677 & ~Ng5857;
  assign n5072 = n6474 & n6475 & (~n6010 | n6476);
  assign n3770_1 = ~n5072;
  assign n5074 = n7226 & n7227 & (n4205 | n7228);
  assign n3783_1 = ~n5074;
  assign n5076 = n7572 & ~n9302 & (~n6889 | ~n8451);
  assign n3797_1 = ~n5076;
  assign n5078 = ~n5991 & n6708 & (~n6860 | ~Ng4498);
  assign n3807_1 = ~n5078;
  assign n5080 = n7870 & n7871 & (Pg35 | ~Ng2719);
  assign n3817_1 = ~n5080;
  assign n5082 = n7795 & (~Pg35 | n7794 | n7796);
  assign n3822_1 = ~n5082;
  assign n5084 = n7109 & n7110 & (n4205 | n7111);
  assign n3837_1 = ~n5084;
  assign n5086 = n6149 & n6150 & (Ng617 | n6151);
  assign n3842_1 = ~n5086;
  assign n5088 = n7915 & (Pg35 | ~Ng324);
  assign n3851_1 = ~n5088;
  assign n5090 = Ng1270 & ~n6829;
  assign n5091 = ~n5965 | ~Ng1536;
  assign n3856 = Ng1274 & (~Pg35 | (n5090 & n5091));
  assign n5093 = n7920 & n7921 & (~n8381 | ~Ng6513);
  assign n3861_1 = ~n5093;
  assign n5095 = n7913 & n7914 & (n7915 | ~Ng305);
  assign n3866_1 = ~n5095;
  assign n5097 = Ng925 & ~n6834;
  assign n3876_1 = Ng930 & (~Pg35 | (n5097 & ~n6128));
  assign n5099 = n6606 & n6607 & (n6433 | ~Ng1906);
  assign n3881_1 = ~n5099;
  assign n3886 = Pg6745 & Pg35;
  assign n5102 = n7865 & (Pg35 | ~\[4428] );
  assign n3896 = ~n5102;
  assign n5104 = n6153 & (Pg35 | ~Ng4907);
  assign n3907_1 = ~n5104;
  assign n5106 = n6163 & (Pg35 | ~Ng4146);
  assign n3912 = ~n5106;
  assign n5108 = n6557 & n6558 & (~n8269 | ~Ng2541);
  assign n3917 = ~n5108;
  assign n5110 = n6587 & (n6395_1 | ~Ng2153);
  assign n3922 = ~n5110;
  assign n5112 = n7901 & (Pg35 | ~Ng225);
  assign n3932 = ~n5112;
  assign n5114 = n7710 & n7711 & (~Ng1874 | ~n8431);
  assign n3937_1 = ~n5114;
  assign n5116_1 = n7135 & n7136 & (n4205 | n7137);
  assign n3942_1 = ~n5116_1;
  assign n5118 = n7872 & n7873 & (Ng1478 | ~n8481);
  assign n3947 = ~n5118;
  assign n5120 = (n6716 | n6722) & (Pg35 | ~Ng3857);
  assign n3952_1 = ~n5120;
  assign n5122 = ~n7705 & (~Pg35 | n7704 | ~Ng1959);
  assign n3957_1 = ~n5122;
  assign n5124 = n7601 & ~n9305 & (~Ng3480 | n7602);
  assign n3962 = ~n5124;
  assign n5126_1 = n6899 & ~n9450 & (n4205 | n6900);
  assign n3967_1 = ~n5126_1;
  assign n5128 = n7779 & (~Pg35 | n6125 | n7778);
  assign n3980_1 = ~n5128;
  assign n3988 = ~n6718 & ~Ng3857;
  assign n5131_1 = Ng499 & (n7986 | ~Ng513);
  assign n5132 = ~n7986 & (~Ng518 | ~n8468);
  assign n3996_1 = Pg35 & (n5131_1 | n5132);
  assign n5134 = n7818 & (~n6638_1 | Ng1002 | n7819);
  assign n4001 = ~n5134;
  assign n5136 = n6255_1 & n6256 & (Ng776 | n6257);
  assign n4006 = ~n5136;
  assign n4015 = ~n6198 & ~Ng4674 & ~Ng4646 & ~Ng4681;
  assign n5139 = n6819 & n6820 & (n6815 | ~Ng1657);
  assign n4025_1 = ~n5139;
  assign n5141_1 = n6376_1 & (n6377 | ~Ng2375);
  assign n4030 = ~n5141_1;
  assign n5143 = (Pg35 | ~Ng278) & (Ng283 | n7834);
  assign n4052_1 = ~n5143;
  assign n5145 = (n6736 | n6742) & (Pg35 | ~Ng3155);
  assign n4057 = ~n5145;
  assign n5147 = ~n7678 & (~Pg35 | n7677 | ~Ng2384);
  assign n4062 = ~n5147;
  assign n5149 = n6213 & (~n6212 | n6214 | ~Ng4608);
  assign n4070_1 = ~n5149;
  assign n5151 = n6415 & n6416 & (~n6004 | n6417_1);
  assign n4080 = ~n5151;
  assign n5153 = n7866 & (Pg35 | ~Ng2791);
  assign n4089_1 = ~n5153;
  assign n5155 = n6187 & n6188 & (Ng613 | n6189);
  assign n4094_1 = ~n5155;
  assign n5157 = n6614 & (Pg35 | ~Ng1840);
  assign n4104 = ~n5157;
  assign n5159 = n7023 & n7024 & (n4205 | n7025);
  assign n4109 = ~n5159;
  assign n5161 = ~n5991 & ~n5993 & (~n6860 | ~Ng4567);
  assign n4114_1 = ~n5161;
  assign n5163 = n7345 & ~n9255 & (Pg35 | ~Ng2518);
  assign n4119 = ~n5163;
  assign n5165 = (~Pg16718 & (~Pg13895 | Pg11349)) | (Pg13895 & Pg11349);
  assign n4124 = n5165 & ~Pg14421 & ~Pg16603 & Pg35 & ~Pg16624;
  assign n5167 = n6339 & (n6340_1 | ~Ng2643);
  assign n4128 = ~n5167;
  assign n5169 = Ng1489 & (~n5170 | ~Ng1495);
  assign n5170 = ~Ng1514 & Pg13272 & ~Ng1526;
  assign n4133_1 = Pg35 & (n5169 | (n5170 & ~Ng1442));
  assign n5172 = n7342 & ~n9254 & (~Ng2551 | n7343);
  assign n4142_1 = ~n5172;
  assign n5174 = n7526 & (n4205 | (Ng5156 & n7527));
  assign n4147 = ~n5174;
  assign n5176 = n6510 & n6511 & (n6512_1 | ~Ng6049);
  assign n4169_1 = ~n5176;
  assign n5178 = n6579 & n6580_1 & (~n8283 | ~Ng2273);
  assign n4174 = ~n5178;
  assign n5180 = n7783 & (~Pg35 | n7782 | n7784);
  assign n4182_1 = ~n5180;
  assign n5182 = n7627 & (n4205 | (Ng3147 & n7628));
  assign n4192_1 = ~n5182;
  assign n5184 = ~Ng3338 | n8509;
  assign n4197 = Ng3343 & (~Pg35 | n5184);
  assign n5186 = n6581 & (Pg35 | ~Ng2265);
  assign n4202_1 = ~n5186;
  assign n5188 = n6115 & n6116 & (Ng626 | n6117);
  assign n4216 = ~n5188;
  assign n5190 = n6333 & n7811 & (~Pg35 | n7812);
  assign n4221_1 = ~n5190;
  assign n5192 = n6518 & n6519 & (n6520 | ~Ng5357);
  assign n4226_1 = ~n5192;
  assign n5194 = n6318 & n6319 & (Pg35 | ~Ng4983);
  assign n4231_1 = ~n5194;
  assign n5196 = n6325 & (Pg35 | ~Ng4785);
  assign n4239_1 = ~n5196;
  assign n5198 = n7029 & n7030 & (n4205 | n7031);
  assign n4254 = ~n5198;
  assign n5200 = n6154 & (Pg35 | ~Ng4922);
  assign n4259_1 = ~n5200;
  assign n5202 = n7597 & n7808 & (Pg35 | ~Ng3965);
  assign n4267_1 = ~n5202;
  assign n5204 = n6872 & n6873 & (Ng918 | ~n8342);
  assign n4277_1 = ~n5204;
  assign n5206 = n6521 & n7860 & (~Pg35 | n7861);
  assign n4282 = ~n5206;
  assign n5208 = n7361 & ~n9265 & (Pg35 | ~Ng2016);
  assign n4291_1 = ~n5208;
  assign n5210 = n7398 & n7399 & (Ng577 | n7400);
  assign n4296_1 = ~n5210;
  assign n5212 = n6471 & n6472_1 & (~n6010 | n6473);
  assign n4301_1 = ~n5212;
  assign n5214 = n7334 & (Pg35 | ~Ng2771);
  assign n4306 = ~n5214;
  assign n5216 = n6643 & n6644 & (Ng930 | ~n5097);
  assign n4316_1 = ~n5216;
  assign n5218 = n7195 & n7196 & (n4205 | n7197);
  assign n4321_1 = ~n5218;
  assign n5220 = (Pg35 | ~Ng812) & (~n7739 | ~n8961);
  assign n4326_1 = ~n5220;
  assign n5222 = ~n8023 & (~Ng837 | (n7758 & ~n8021));
  assign n4336_1 = ~n5222;
  assign n5224 = n6489 & (Ng599 | n6490) & ~n9446;
  assign n4344_1 = ~n5224;
  assign n5226 = n7929 & n7930 & (~n8394 | ~Ng5475);
  assign n4349_1 = ~n5226;
  assign n5228 = (n7742 | n7743) & (Pg35 | ~Ng736);
  assign n4354_1 = ~n5228;
  assign n5230 = n7015 & n7016 & (n4205 | n7017);
  assign n4359_1 = ~n5230;
  assign n5232 = (Pg35 | ~Ng6741) & (n6497_1 | ~n9420);
  assign n4364_1 = ~n5232;
  assign n5234 = n6174 & (Pg35 | ~Ng2868);
  assign n4374_1 = ~n5234;
  assign n5236 = n7940 & ~n9350 & (n7941 | ~Ng5080);
  assign n4384_1 = ~n5236;
  assign n5238 = n7070 & n7071 & (n4205 | n7072);
  assign n4389_1 = ~n5238;
  assign n5240 = (n6359_1 | ~Ng2495) & (n6561 | ~Ng2465);
  assign n4397_1 = ~n5240;
  assign n5242 = n6367 & n6368 & (~n6002 | n6369_1);
  assign n4402_1 = ~n5242;
  assign n5244 = n7359 & (Pg35 | ~Ng2098);
  assign n4407_1 = ~n5244;
  assign n5246 = n6344 & n6345 & (~n6000 | ~n8265);
  assign n4417_1 = ~n5246;
  assign n5248 = n6314 & (Pg35 | ~Ng4975);
  assign n4427_1 = ~n5248;
  assign n5250 = n6331 & n6332 & (n6323 | ~Ng4785);
  assign n4437 = ~n5250;
  assign n5252 = n7084 & n7085 & (n4205 | n7086);
  assign n4442_1 = ~n5252;
  assign n5254 = n6184 & n6185 & (Ng781 | n6186);
  assign n4447 = ~n5254;
  assign n5256 = n7981 & n7982 & (n7983 | ~Ng686);
  assign n4465_1 = ~n5256;
  assign n5258 = n7815 & n7816 & (Ng1252 | n7817);
  assign n4470 = ~n5258;
  assign n5260 = (n7750 | n7751) & (Pg35 | ~Ng667);
  assign n4475 = ~n5260;
  assign n5262 = n6971 & ~n9453 & (n4205 | n6972);
  assign n4485 = ~n5262;
  assign n5264 = (~Ng5523 | n6686) & (~Ng5527 | n6687);
  assign n4499 = ~n5264;
  assign n5266 = n6827 & n6828 & (Ng1270 | n6829);
  assign n4514 = ~n5266;
  assign n5268 = n6315_1 & (n6316 | n6317 | ~Ng4991);
  assign n4519 = ~n5268;
  assign n5270 = (Pg35 | ~Ng6219) & (n6665_1 | n6666);
  assign n4524 = ~n5270;
  assign n5272 = n7201 & n7202 & (n4205 | n7203);
  assign n4529 = ~n5272;
  assign n5274 = n7496 & (n4205 | (Ng5503 & n7497));
  assign n4534 = ~n5274;
  assign n5276 = n7032 & n7033 & (n4205 | n7034);
  assign n4544_1 = ~n5276;
  assign n5278 = n7147 & n7148 & (n4205 | n7149);
  assign n4559_1 = ~n5278;
  assign n5280 = n6423 & n6424 & (~n6004 | n6425);
  assign n4564_1 = ~n5280;
  assign n4569_1 = ~n6668 & ~Ng6203;
  assign n5283 = n7350 & ~n9258 & (Pg35 | ~Ng2384);
  assign n4582_1 = ~n5283;
  assign n5285 = n6370 & n6371 & (~n6002 | n6372);
  assign n4592 = ~n5285;
  assign n5287 = n6240_1 & (n6241 | n6239 | n6229);
  assign n4597_1 = ~n5287;
  assign n5289 = n6138 & n6139;
  assign n4602 = ~n5289;
  assign n5291 = n6546_1 & n6547 & (~n8262 | ~Ng2675);
  assign n4607 = ~n5291;
  assign n5293 = n7996 & (Pg35 | ~Ng4358);
  assign n4612 = ~n5293;
  assign n4617 = ~n6193 & ~Ng4864 & ~Ng4871 & ~Ng4836;
  assign n5296 = n7102 & n7103 & (n4205 | n7104);
  assign n4631 = ~n5296;
  assign n5298_1 = n6183_1 & (Pg35 | ~Ng2130);
  assign n4636 = ~n5298_1;
  assign n5300 = n6567 & ~n9430 & (~Ng2338 | n6566);
  assign n4644 = ~n5300;
  assign n5302 = n6990 & n6991 & (n4205 | n6992);
  assign n4652_1 = ~n5302;
  assign n5304 = n7867 & (Pg35 | ~Ng2779);
  assign n4657_1 = ~n5304;
  assign n5306 = n7188 & n7189 & (n4205 | n7190);
  assign n4662 = ~n5306;
  assign n5308 = n7018 & n7019 & (n4205 | n7020);
  assign n4672_1 = ~n5308;
  assign n5310 = n7132 & n7133 & (n4205 | n7134);
  assign n4677_1 = ~n5310;
  assign n5312 = n6333 & n6541_1 & (Ng2759 | n6542);
  assign n4682 = ~n5312;
  assign n5314 = n6498 & n6499 & (n6500 | ~Ng6741);
  assign n4687 = ~n5314;
  assign n5316 = n6146 & n6147_1 & (Ng785 | n6148);
  assign n4692_1 = ~n5316;
  assign n5318_1 = n7382 & n7383 & (Ng1259 | n7384);
  assign n4697_1 = ~n5318_1;
  assign n5320 = n7600 & (Pg35 | ~Ng3480);
  assign n4702_1 = ~n5320;
  assign n5322_1 = n6930 & n6931 & (n4205 | n6932);
  assign n4712_1 = ~n5322_1;
  assign n5324 = (n6685 | n6691) & (Pg35 | ~Ng5511);
  assign n4717_1 = ~n5324;
  assign n5326 = n6360 & ~n9443 & (~n6002 | n6361);
  assign n4722_1 = ~n5326;
  assign n5328 = n6346 & n6347 & (~n6000 | n6348);
  assign n4727_1 = ~n5328;
  assign n5330 = n7892 & n7893 & (Pg35 | ~Ng921);
  assign n4741_1 = ~n5330;
  assign n5332 = n7360 & ~n9264 & (Pg35 | ~Ng2093);
  assign n4746 = ~n5332;
  assign n5334 = (~Pg35 | n6290) & (~Ng4473 | n6292);
  assign n4751_1 = ~n5334;
  assign n5336 = n6296 & (Ng604 | n6297_1) & ~n9442;
  assign n4756 = ~n5336;
  assign n5338 = n6896 & n6897 & (n4205 | n6898);
  assign n4761_1 = ~n5338;
  assign n5340 = n6437_1 & n6438 & (~n6006 | ~n8302);
  assign n4766 = ~n5340;
  assign n5342 = n6445 & n6446 & (~n6006 | n6447_1);
  assign n4782 = ~n5342;
  assign n5344 = n6161 & (Pg35 | ~Ng4253);
  assign n4787_1 = ~n5344;
  assign n5346 = ~n7714 & (~Pg35 | n7712 | ~Ng1825);
  assign n4792_1 = ~n5346;
  assign n5348 = ~n7973 & (~Ng969 | (Pg35 & n4558));
  assign n4797 = ~n5348;
  assign n5350 = n7843 & (Pg35 | ~Ng4417);
  assign n4802 = ~n5350;
  assign n5352 = n7231 & n7232 & (n4205 | n7233);
  assign n4807_1 = ~n5352;
  assign n5354 = n7138 & n7139 & (n4205 | n7140);
  assign n4812 = ~n5354;
  assign n5356 = n7371 & ~n9271 & (Pg35 | ~Ng1748);
  assign n4817 = ~n5356;
  assign n5358 = (n6192_1 | n6193) & (Pg35 | ~Ng4849);
  assign n4822 = ~n5358;
  assign n5360 = n7204 & n7205 & (n4205 | n7206);
  assign n4827 = ~n5360;
  assign n5362 = n7408 & ~n9278 & (~n8213 | ~n8440);
  assign n4832_1 = ~n5362;
  assign n4837_1 = Pg35 & ~n8535;
  assign n5365 = n7674 & n7675 & (~Ng2433 | ~n8418);
  assign n4842_1 = ~n5365;
  assign n5367 = n6783 & n6779 & n6784;
  assign n4859_1 = ~n5367;
  assign n4864_1 = ~n6175;
  assign n5370 = (n6414 | ~Ng2070) & (n6594 | ~Ng2040);
  assign n4873_1 = ~n5370;
  assign n5372 = (~Pg16775 & (~Pg13966 | Pg11418)) | (Pg13966 & Pg11418);
  assign n4887_1 = n5372 & ~Pg14518 & ~Pg16659 & Pg35 & ~Pg16693;
  assign n5374 = n7436 & (Pg35 | ~Ng6177);
  assign n4899 = ~n5374;
  assign n5376 = n7096 & n7097 & (n4205 | n7098);
  assign n4914_1 = ~n5376;
  assign n5378 = Ng1395 ^ n7877;
  assign n4919_1 = Pg35 & n5378 & ~Ng1322;
  assign n5380 = n6600_1 & ~n9433 & (~Ng1913 | n6599);
  assign n4924_1 = ~n5380;
  assign n5382 = n6573 & n6574 & (n6377 | ~Ng2331);
  assign n4929_1 = ~n5382;
  assign n5384 = n6984 & n6985 & (n4205 | n6986);
  assign n4934_1 = ~n5384;
  assign n5386 = n7191 & ~n9464 & (n4205 | n7192);
  assign n4944 = ~n5386;
  assign n5388 = (~Ng1266 | n7967) & (n7966 | ~Ng1249);
  assign n4958_1 = ~n5388;
  assign n5390 = n7498 & (Pg35 | ~Ng5485);
  assign n4963_1 = ~n5390;
  assign n5392 = n7746 & n7747 & (Pg35 | ~Ng676);
  assign n4968_1 = ~n5392;
  assign n5394 = n6864 & n6865 & (Pg35 | ~Ng2741);
  assign n4973 = ~n5394;
  assign n5396 = n7501 & ~n9290 & (~n8100 | ~n8446);
  assign n4978 = ~n5396;
  assign n5398 = n6706 & n6861 & (Pg35 | ~Ng4423);
  assign n4983_1 = ~n5398;
  assign n5400 = n6892 & n6893 & (n4205 | n6894);
  assign n4992 = ~n5400;
  assign n5402 = n6362 & n6363 & (~n6002 | ~n8272);
  assign n4997 = ~n5402;
  assign n5404 = n6401 & n6402 & (~n6008_1 | n6403_1);
  assign n5002 = ~n5404;
  assign n5406 = n6757 & n6758 & (~Ng2491 | n6756);
  assign n5011_1 = ~n5406;
  assign n5408 = n6194 & ~n9439 & (Pg35 | ~Ng4843);
  assign n5016 = ~n5408;
  assign n5410 = n6404 & n6405 & (~n6008_1 | n6406);
  assign n5021 = ~n5410;
  assign n5412 = n7352 & ~n9260 & (~Ng2283 | n7353);
  assign n5026 = ~n5412;
  assign n5414 = n6939 & n6940 & (n4205 | n6941);
  assign n5031_1 = ~n5414;
  assign n5416_1 = n7334 & (Pg35 | ~Ng2831);
  assign n5036 = ~n5416_1;
  assign n5418 = n6568 & n6569 & (~n8276 | ~Ng2407);
  assign n5041 = ~n5418;
  assign n5420 = n6173 & (Pg35 | ~Ng2988);
  assign n5046_1 = ~n5420;
  assign n5422 = n7869 & (Pg35 | ~Ng2763);
  assign n5051_1 = ~n5422;
  assign n5424 = n6631 & ~n9356 & (n5964 | Ng1351);
  assign n5425 = ~n6631 | n8082;
  assign n5064 = Pg35 & (n5424 | (Ng1312 & n5425));
  assign n5427 = n7112 & n7113 & (n4205 | n6692);
  assign n5069 = ~n5427;
  assign n5429 = n6160_1 & (Pg35 | ~Ng4249);
  assign n5074_1 = ~n5429;
  assign n5431 = (n7826 | ~Ng446) & (~Ng645 | ~n8475);
  assign n5079_1 = ~n5431;
  assign n5433 = n7906 & ~n8132 & (Pg35 | ~Ng728);
  assign n5088_1 = ~n5433;
  assign n5435 = n7990 & (Pg35 | ~Ng405);
  assign n5093_1 = ~n5435;
  assign n5437 = n7885 & n7886 & (Ng1129 | ~n8487);
  assign n5098 = ~n5437;
  assign n5439 = (n6395_1 | ~Ng2227) & (n6583 | ~Ng2197);
  assign n5103 = ~n5439;
  assign n5441 = n7370 & ~n9270 & (Pg35 | ~Ng1825);
  assign n5116 = ~n5441;
  assign n5443 = n7248 & ~n9467 & (n4205 | n7249);
  assign n5121 = ~n5443;
  assign n5445 = n8030 & n8031 & (Pg35 | ~Ng401);
  assign n5126 = ~n5445;
  assign n5447 = n6630 & (n6470 | ~Ng1592);
  assign n5131 = ~n5447;
  assign n5449 = n8012 & n8013 & (Ng1221 | ~n8497);
  assign n5141 = ~n5449;
  assign n5451 = n7035 & n7036 & (n4205 | n7037);
  assign n5146 = ~n5451;
  assign n5453 = (n7401 | n7402) & (Pg35 | ~Ng142);
  assign n5156 = ~n5453;
  assign n5455 = n6797 & n6798 & (~Ng1932 | n6796);
  assign n5165_1 = ~n5455;
  assign n5457 = n6823 & n6819 & n6824;
  assign n5170_1 = ~n5457;
  assign n5459 = n7525 & ~n9292 & (Pg35 | ~Ng5467);
  assign n5180_1 = ~n5459;
  assign n5461_1 = ~Pg35 | ~Ng2689;
  assign n5185_1 = ~n5461_1;
  assign n5463 = (Pg35 | ~Ng6565) & (n6655 | n6656_1);
  assign n5190_1 = ~n5463;
  assign n5465 = n7728 & n7729 & (~Ng1604 | ~n8437);
  assign n5195_1 = ~n5465;
  assign n5467 = n6793 & n6794 & (Pg35 | ~Ng2036);
  assign n5200_1 = ~n5467;
  assign n5469 = n6548 & (Pg35 | ~Ng2667);
  assign n5205_1 = ~n5469;
  assign n5471 = n8009 & n8010 & (~Pg17423 | n8005);
  assign n5210_1 = ~n5471;
  assign n5473 = n7856 & n7859 & (Pg35 | ~Ng4411);
  assign n5214_1 = ~n5473;
  assign n5475 = n6612 & n6613 & (~n8305 | ~Ng1848);
  assign n5218_1 = ~n5475;
  assign n5477 = n7935 & ~n9474 & (\[4434]  | n7936);
  assign n5223_1 = ~n5477;
  assign n5479 = n7499 & ~n9289 & (~Ng5485 | n7500);
  assign n5228_1 = ~n5479;
  assign n5481 = (n7335 | n7336) & (Pg35 | ~Ng2735);
  assign n5233_1 = ~n5481;
  assign n5483 = n7665 & n7666 & (~Ng2567 | ~n8414);
  assign n5241_1 = ~n5483;
  assign n5485 = n7798 & n7799 & (n7800 | n7801);
  assign n5246_1 = ~n5485;
  assign n5487 = n6224 & n6225 & (Pg35 | ~Ng4311);
  assign n5251 = ~n5487;
  assign n5489 = n7021 & ~n9457 & (n4205 | n7022);
  assign n5256_1 = ~n5489;
  assign n5491 = n6622 & ~n9435 & (~Ng1644 | n6621);
  assign n5273 = ~n5491;
  assign n5493 = n6648 & (Ng595 | n6649) & ~n9447;
  assign n5278_1 = ~n5493;
  assign n5495 = n6779 & n6780 & (n6775 | ~Ng2217);
  assign n5283_1 = ~n5495;
  assign n5497 = Ng1404 ^ n8011;
  assign n5288_1 = n5497 | ~n9150;
  assign n5499 = n6787 & n6788 & (~Ng2066 | n6786);
  assign n5293_1 = ~n5499;
  assign n5501 = n7128 & ~n9461 & (n4205 | n7129);
  assign n5303_1 = ~n5501;
  assign n5503 = n6392 & (Pg35 | ~Ng2246);
  assign n5308_1 = ~n5503;
  assign n5505 = n6349_1 & n6350 & (~n6000 | n6351);
  assign n5313_1 = ~n5505;
  assign n5507 = (n6697 | n6698) & (Pg35 | ~Ng5170);
  assign n5318 = ~n5507;
  assign n5509 = n7862 & (Pg35 | ~Ng2823);
  assign n5331_1 = ~n5509;
  assign n5511 = n6190 & (n6191 | ~Ng4854 | ~n8228);
  assign n5339_1 = ~n5511;
  assign n5513 = n6636 & n6637 & (Ng1274 | ~n5090);
  assign n5349 = ~n5513;
  assign n5515 = n6237 & (n6228 | n6236 | n6238);
  assign n5361_1 = ~n5515;
  assign n5517 = n6358 & (n6359_1 | ~Ng2509);
  assign n5371_1 = ~n5517;
  assign n5519 = n7881 & n7882 & (Pg35 | ~Ng1266);
  assign n5381_1 = ~n5519;
  assign n5521 = n6913 & ~n9451 & (n4205 | n6914);
  assign n5393_1 = ~n5521;
  assign n5523 = n7531 & ~n9294 & (~n6885 | ~n8449);
  assign n5398_1 = ~n5523;
  assign n5525 = n6957 & n6958 & (n4205 | n6959);
  assign n5406_1 = ~n5525;
  assign n5527 = n6137_1 & (Pg35 | ~Ng2999);
  assign n5416 = ~n5527;
  assign n5529 = n7827 & (Pg35 | ~Ng699);
  assign n5421_1 = ~n5529;
  assign n5531 = n6627 & n6628 & (n6470 | ~Ng1636);
  assign n5426_1 = ~n5531;
  assign n5533 = n7207 & n7208 & (n4205 | n7209);
  assign n5431_1 = ~n5533;
  assign n5535 = ~n7696 & (~Pg35 | n7695 | ~Ng2093);
  assign n5436 = ~n5535;
  assign n5537 = (Pg35 | ~Ng1052) & (n7889 | ~n9148);
  assign n5451_1 = ~n5537;
  assign n5539 = n6396 & n6397 & (~n6008_1 | n6398);
  assign n5461 = ~n5539;
  assign n5541 = n7968 & n7969 & (Ng956 | ~n8498);
  assign n5466_1 = ~n5541;
  assign n5543 = n6453 & ~n9445 & (~n5998_1 | n6454);
  assign n5471_1 = ~n5543;
  assign n5545 = n7465 & (n4205 | (Ng5849 & n7466));
  assign n5476_1 = ~n5545;
  assign n5547 = n7337 & ~n9251 & (~Ng2685 | n7338);
  assign n5486_1 = ~n5547;
  assign n5549 = n6584 & n6585_1 & (n6395_1 | ~Ng2197);
  assign n5491_1 = ~n5549;
  assign n5551 = n6565_1 & (n6359_1 | ~Ng2421);
  assign n5496_1 = ~n5551;
  assign n5553 = n7891 & ~n9438 & (Pg35 | ~Ng1041);
  assign n5501_1 = ~n5553;
  assign n5555 = n7755 & n7832 & (~Pg35 | n7833);
  assign n5506_1 = ~n5555;
  assign n5557 = ~Ng4405 & (n7846 | ~Ng4388 | n7853);
  assign n5511_1 = ~n5557;
  assign n5559 = n5958 & (~Ng1536 | (Ng1526 & ~Ng1514));
  assign n5560 = Pg7946 ^ Ng1514;
  assign n5516_1 = Pg35 & (n5559 | n5560);
  assign n5562 = (~Ng6561 | n6657) & (~Ng6565 | n6658);
  assign n5526_1 = ~n5562;
  assign n5564 = n6168 & (Pg35 | ~Ng2936);
  assign n5531_1 = ~n5564;
  assign n5566 = n7813 & (~n6631 | Ng1345 | n7814);
  assign n5536_1 = ~n5566;
  assign n5568 = ~Pg35 | ~Ng4727;
  assign n5549_1 = ~n5568;
  assign n5570 = (~Pg17778 & (~Pg14828 | Pg12470)) | (Pg14828 & Pg12470);
  assign n5554_1 = n5570 & ~Pg13099 & ~Pg17688 & Pg35 & ~Pg17722;
  assign n5572 = n7193 & ~n9465 & (n4205 | n7194);
  assign n5563_1 = ~n5572;
  assign n5574 = n7367 & ~n9269 & (~Ng1858 | n7368);
  assign n5578_1 = ~n5574;
  assign n5576 = n7895 & (Pg35 | ~Ng246);
  assign n5583_1 = ~n5576;
  assign n5578 = n7315 & n7316 & (n4205 | n7317);
  assign n5588_1 = ~n5578;
  assign n5580 = n7719 & n7720 & (~Ng1740 | ~n8434);
  assign n5593_1 = ~n5580;
  assign n5582 = n6933 & n6934 & (n4205 | n6935);
  assign n5598 = ~n5582;
  assign n5584 = n6364 & n6365 & (~n6002 | n6366);
  assign n5603_1 = ~n5584;
  assign n5586 = n6430 & (Pg35 | ~Ng1955);
  assign n5608_1 = ~n5586;
  assign n5588 = n6942 & n6943 & (n4205 | n6944);
  assign n5618_1 = ~n5588;
  assign n5590 = n6895 & ~n9449 & (n4205 | n6654);
  assign n5623_1 = ~n5590;
  assign n5592 = n7234 & n7235 & (n4205 | n7236);
  assign n5628 = ~n5592;
  assign n5594 = n6603 & (Pg35 | ~Ng1974);
  assign n5638 = ~n5594;
  assign n5596 = n6477_1 & n6478 & (~n6010 | n6479);
  assign n5643_1 = ~n5596;
  assign n5598_1 = n6601 & n6602 & (~n8298 | ~Ng1982);
  assign n5658_1 = ~n5598_1;
  assign n5600 = n7144 & n7145 & (n4205 | n7146);
  assign n5666_1 = ~n5600;
  assign n5602 = n7802 & n7803 & (n7801 | ~n8472);
  assign n5671 = ~n5602;
  assign n5604 = ~Ng6381 | n8503;
  assign n5676_1 = Ng6386 & (~Pg35 | n5604);
  assign n5606 = n6848 & ~n9232 & (Pg35 | ~Ng5029);
  assign n5695 = ~n5606;
  assign n5608 = n6158 & (Pg35 | ~Ng4732);
  assign n5700_1 = ~n5608;
  assign n5610 = n7567 & (n4205 | (Ng3849 & n7568));
  assign n5710_1 = ~n5610;
  assign n5612 = n7324 & n7325 & (n4205 | n7326);
  assign n5718 = ~n5612;
  assign n5614 = n7925 & (Pg35 | ~Ng5841);
  assign n5723_1 = ~n5614;
  assign n5616 = n6320_1 & n6321 & (n6312 | ~Ng4975);
  assign n5728 = ~n5616;
  assign n5618 = n6129 & n6130 & (Ng790 | n6131);
  assign n5733_1 = ~n5618;
  assign n5620 = n7000 & n7001 & (n4205 | n7002);
  assign n5738_1 = ~n5620;
  assign n5622 = n7366 & ~n9268 & (Pg35 | ~Ng1882);
  assign n5743_1 = ~n5622;
  assign n5624 = n7439 & ~n9282 & (~n6886 | ~n8442);
  assign n5748 = ~n5624;
  assign n5626 = n7762 & (Pg35 | ~Ng5619);
  assign n5758_1 = ~n5626;
  assign n5628_1 = (n7774 | ~n9144) & (n7775 | ~Ng4939);
  assign n5763 = ~n5628_1;
  assign n5630 = n7321 & n7322 & (n4205 | n7323);
  assign n5772 = ~n5630;
  assign n5632 = n7288 & n7289 & (n4205 | n7290);
  assign n5781_1 = ~n5632;
  assign n5634 = n7528 & (Pg35 | ~Ng5138);
  assign n5786 = ~n5634;
  assign n5636 = n7130 & ~n9462 & (n4205 | n7131);
  assign n5791 = ~n5636;
  assign n5638_1 = n7357 & ~n9263 & (~Ng2126 | n7358);
  assign n5796 = ~n5638_1;
  assign n5640 = n7365 & ~n9267 & (Pg35 | ~Ng1959);
  assign n5811 = ~n5640;
  assign n5642 = n7937 & n7938 & (Ng5097 | ~n8494);
  assign n5816_1 = ~n5642;
  assign n5644 = n7318 & n7319 & (n4205 | n7320);
  assign n5821_1 = ~n5644;
  assign n5646 = ~n7851 & ((Pg35 & Ng4388) | ~Ng4430);
  assign n5833_1 = ~n5646;
  assign n5648 = n7868 & (Pg35 | ~Ng2767);
  assign n5838_1 = ~n5648;
  assign n5650 = n7848 & n7849 & (n7844 | n7846);
  assign n5846 = ~n5650;
  assign n5652 = n6866 & n6867 & (Pg35 | ~Ng1361);
  assign n5855_1 = ~n5652;
  assign n5654 = n6407 & n6408 & (~n6008_1 | n6409);
  assign n5869 = ~n5654;
  assign n5656 = (n6377 | ~Ng2361) & (n6572 | ~Ng2331);
  assign n5879_1 = ~n5656;
  assign n5658 = n6877 & n6878 & (Ng582 | n6879);
  assign n5888_1 = ~n5658;
  assign n5660 = n7351 & ~n9259 & (Pg35 | ~Ng2307);
  assign n5903_1 = ~n5660;
  assign n5662_1 = n7820 & n7821 & (Ng907 | n7822);
  assign n5908_1 = ~n5662_1;
  assign n5664 = n7369 & (Pg35 | ~Ng1830);
  assign n5918_1 = ~n5664;
  assign n5666 = n7245 & n7246 & (n4205 | n7247);
  assign n5923_1 = ~n5666;
  assign n5668 = Ng2932 | Ng2999;
  assign n5669 = n6085 & n6082 & n6083 & n6084;
  assign n5928_1 = n5668 & Pg35;
  assign n5671_1 = n6385_1 & n6386 & (~n6012_1 | n6387);
  assign n5933_1 = ~n5671_1;
  assign n5673 = n7825 & n7826 & (Pg35 | ~Ng681);
  assign n5941_1 = ~n5673;
  assign n5675 = n7740 & n7741 & (Pg35 | ~Ng827);
  assign n5946_1 = ~n5675;
  assign n5677 = n6513 & n6514 & (Pg35 | ~Ng5698);
  assign n5951_1 = ~n5677;
  assign n5679 = n6556 & ~n9429 & (~Ng2472 | n6555_1);
  assign n5961_1 = ~n5679;
  assign n5681 = n7012 & n7013 & (n4205 | n7014);
  assign n5966_1 = ~n5681;
  assign n5683 = n6449 & (Pg35 | ~Ng1821);
  assign n5975_1 = ~n5683;
  assign n5685 = n7270 & n7271 & (n4205 | n7272);
  assign n5980_1 = ~n5685;
  assign n5687 = n7948 & (Pg35 | ~Ng3841);
  assign n5985_1 = ~n5687;
  assign n5689 = n6590_1 & n6591 & (~n8291 | ~Ng2116);
  assign n5990 = ~n5689;
  assign n5691 = n7285 & n7286 & (n4205 | n7287);
  assign n5998 = ~n5691;
  assign n5693 = n7172 & n7173 & (n4205 | n7174);
  assign n6003_1 = ~n5693;
  assign n5695_1 = n6181 & (Pg35 | ~Ng2689);
  assign n6032_1 = ~n5695_1;
  assign n5697 = ~n8329 & (Pg35 | ~Ng4382);
  assign n6037_1 = ~n5697;
  assign n5699 = (n6658 | n6659) & (Pg35 | ~Ng6555);
  assign n6042 = ~n5699;
  assign n5701 = n7734 & (n7735 | ~Ng1141);
  assign n6047_1 = ~n5701;
  assign n5703 = n6625 & (Pg35 | ~Ng1706);
  assign n6061 = ~n5703;
  assign n5705 = n7405 & (Pg35 | ~Ng6523);
  assign n6066_1 = ~n5705;
  assign n5707 = n7291 & n7292 & (n4205 | n7293);
  assign n6071_1 = ~n5707;
  assign n5709 = ~n7723 & (~Pg35 | n7721 | ~Ng1691);
  assign n6076_1 = ~n5709;
  assign n5711 = n6169_1 & (Pg35 | ~Ng2922);
  assign n6081 = ~n5711;
  assign n5713 = n7931 & (Pg35 | ~Ng5148);
  assign n6091 = ~n5713;
  assign n5715 = ~\[4415]  | n8506;
  assign n6096 = Ng5348 & (~Pg35 | n5715);
  assign n5717 = n6243 & (n6241 | n6242 | n6232);
  assign n6104 = ~n5717;
  assign n5719 = n6170 & (Pg35 | ~Ng2912);
  assign n6109_1 = ~n5719;
  assign n5721 = n7047 & n7048 & (n4205 | n7049);
  assign n6119_1 = ~n5721;
  assign n5723 = n6924 & n6925 & (n4205 | n6926);
  assign n6127 = ~n5723;
  assign n5725 = n6789 & n6790 & (n6785 | ~Ng2060);
  assign n6132_1 = ~n5725;
  assign n5727 = n7073 & n7074 & (n4205 | n7075);
  assign n6142 = ~n5727;
  assign n5729 = Pg135 | n6097;
  assign n5730 = ~Ng4349 | ~Ng4358;
  assign n5731 = ~Ng4633 | n8232;
  assign n6152 = Pg35 & (n5729 | n5730 | n5731);
  assign n5733 = n7630 & ~n9309 & (n7631 | ~Ng3129);
  assign n6165 = ~n5733;
  assign n5735 = (n6695 | n6701) & (Pg35 | ~Ng5164);
  assign n6174_1 = ~n5735;
  assign n5737 = n7926 & n7927 & (~n8390 | ~Ng5821);
  assign n6183 = ~n5737;
  assign n5739 = n6960 & n6961 & (n4205 | n6962);
  assign n6188_1 = ~n5739;
  assign n5741 = n7701 & n7702 & (~Ng2008 | ~n8428);
  assign n6196 = ~n5741;
  assign n5743 = n6533 & n6534 & (n6535 | ~Ng3703);
  assign n6206 = ~n5743;
  assign n5745 = n6142_1 & n6143;
  assign n6216 = ~n5745;
  assign n5747 = n7757 & ~n9330 & (n7758 | ~Ng411);
  assign n6221 = ~n5747;
  assign n5749 = n7186 & ~n9463 & (n4205 | n7187);
  assign n6230 = ~n5749;
  assign n5751 = n6180 & (Pg35 | ~Ng2697);
  assign n6235 = ~n5751;
  assign n5753_1 = n7960 & n7961 & (Ng1300 | ~n8496);
  assign n6245 = ~n5753_1;
  assign n5755 = n7156 & n7157 & (n4205 | n7158);
  assign n6255 = ~n5755;
  assign n5757 = n6854 & (n6855 | ~Ng5046 | ~n8722);
  assign n6265 = ~n5757;
  assign n5759 = ~n7687 & (~Pg35 | n7686 | ~Ng2250);
  assign n6270 = ~n5759;
  assign n5761 = ~n5991 & n6706 & (~n6860 | ~Ng4546);
  assign n6279 = ~n5761;
  assign n5763_1 = n6763 & n6764 & (Pg35 | ~Ng2461);
  assign n6284 = ~n5763_1;
  assign n5765 = n6171 & (Pg35 | ~Ng2907);
  assign n6297 = ~n5765;
  assign n5767 = n6767 & n6768 & (~Ng2357 | n6766);
  assign n6302 = ~n5767;
  assign n5769 = n6880 & n6881 & (Pg35 | ~Ng146);
  assign n6310 = ~n5769;
  assign n5771 = n6162 & (Pg35 | ~Ng4300);
  assign n6315 = ~n5771;
  assign n5773 = n6858 & (n6855 | Ng5016 | ~n8380);
  assign n6320 = ~n5773;
  assign n5775 = n7955 & n7956 & (~n8409 | ~Ng3119);
  assign n6325_1 = ~n5775;
  assign n5777 = ~n7965 & (~Ng1312 | (Pg35 & n5425));
  assign n6330 = ~n5777;
  assign n5779 = n7553 & (Ng5115 | n7554) & ~n9296;
  assign n6344_1 = ~n5779;
  assign n5781 = n6539 & n6540 & (Pg35 | ~Ng3347);
  assign n6349 = ~n5781;
  assign n5783 = n6891 & (Pg35 | ~Ng6653);
  assign n6354 = ~n5783;
  assign n5785 = n7219 & n7220 & (n4205 | n7221);
  assign n6364_1 = ~n5785;
  assign n5787 = n7280 & n7281 & (n4205 | n7282);
  assign n6369 = ~n5787;
  assign n5789 = n7076 & ~n9459 & (n4205 | n7077);
  assign n6380 = ~n5789;
  assign n5791_1 = n7225 & (Pg35 | ~Ng3610);
  assign n6385 = ~n5791_1;
  assign n5793 = n6176 & (Pg35 | ~Ng2860);
  assign n6390 = ~n5793;
  assign n5795 = n7949 & n7950 & (~n8401 | ~Ng3821);
  assign n6403 = ~n5795;
  assign n5797 = n7944 & n7945 & (Pg35 | ~Ng4057);
  assign n6408_1 = ~n5797;
  assign n5799 = n7108 & (Pg35 | ~Ng5268);
  assign n6417 = ~n5799;
  assign n5801_1 = n6333 & n7656 & (Ng2735 | n7657);
  assign n6422 = ~n5801_1;
  assign n5803 = n6963 & n6964 & (n4205 | n6965);
  assign n6432 = ~n5803;
  assign n5805 = n7339 & (Pg35 | ~Ng2657);
  assign n6437 = ~n5805;
  assign n5807 = n7932 & n7933 & (n7934 | ~Ng5128);
  assign n6447 = ~n5807;
  assign n5809 = n7655 & ~n9312 & (Pg35 | ~Ng3111);
  assign n6457 = ~n5809;
  assign n5811_1 = n6199 & ~n9440 & (Pg35 | ~Ng4653);
  assign n6462 = ~n5811_1;
  assign n5813 = (Pg35 | ~Ng4349) & (n5968 | ~n8636);
  assign n6467 = ~n5813;
  assign n5815 = n6809 & n6810 & (n6805 | ~Ng1792);
  assign n6472 = ~n5815;
  assign n5817 = n6413_1 & (n6414 | ~Ng2084);
  assign n6477 = ~n5817;
  assign n5819 = n7330 & n7331 & (n4205 | n7332);
  assign n6482 = ~n5819;
  assign n5821 = n8233 ^ Ng4311;
  assign n6487 = n5821 & ~n8235;
  assign n5823 = n6341 & n6342 & (~n6000 | n6343);
  assign n6492 = ~n5823;
  assign n5825 = n7327 & n7328 & (n4205 | n7329);
  assign n6517 = ~n5825;
  assign n5827 = n7991 & n7992 & (Ng385 | n7993);
  assign n6541 = ~n5827;
  assign n5829 = n6426 & n6427_1 & (~n6004 | n6428);
  assign n6546 = ~n5829;
  assign n5831 = n7344 & (Pg35 | ~Ng2523);
  assign n6551 = ~n5831;
  assign n5833 = n7312 & n7313 & (n4205 | n7314);
  assign n6580 = ~n5833;
  assign n5835 = n6166 & (Pg35 | ~Ng2960);
  assign n6585 = ~n5835;
  assign n5837 = ~Ng5689 | ~n8505;
  assign n6590 = Ng5694 & (~Pg35 | n5837);
  assign n5839 = n7123 & ~n9460 & (n4205 | n7124);
  assign n6595 = ~n5839;
  assign n5841 = (~Ng3518 | n6727) & (~Ng3522 | n6728);
  assign n6605 = ~n5841;
  assign n5843 = n7632 & ~n9310 & (~n6890 | ~n8456);
  assign n6610 = ~n5843;
  assign n5845 = n7294 & n7295 & (n4205 | n7296);
  assign n6615 = ~n5845;
  assign n5847 = n7843 & (Pg35 | ~Ng4455);
  assign n6620 = ~n5847;
  assign n5849 = n6210 & n6211_1 & (n6206_1 | ~Ng4628);
  assign n6624 = ~n5849;
  assign n5851 = n6598 & (n6414 | ~Ng1996);
  assign n6629 = ~n5851;
  assign n5853 = n7841 & ~n8127 & (Pg35 | ~Ng4527);
  assign n6638 = ~n5853;
  assign n5855 = n7372 & ~n9272 & (~Ng1724 | n7373);
  assign n6651 = ~n5855;
  assign n5857 = (~Ng1379 | ~n9115) & (n6635 | ~Ng1373);
  assign n6656 = ~n5857;
  assign n5859_1 = (~Pg16744 & (~Pg13926 | Pg11388)) | (Pg13926 & Pg11388);
  assign n6661 = n5859_1 & ~Pg14451 & ~Pg16627 & Pg35 & ~Pg16656;
  assign n5861 = n6442_1 & n6443 & (~n6006 | n6444);
  assign n6665 = ~n5861;
  assign n5863 = n7053 & (Pg35 | ~Ng5615);
  assign n6670 = ~n5863;
  assign n5865 = Pg35 & (Ng5845 | Ng5831);
  assign n5866 = Ng2724 | Ng2729;
  assign n5867 = n8206 & Ng2735;
  assign n5868 = ~n8373 & (n5866 | (n5867 & ~Ng2771));
  assign n5869_1 = n6058 & n6059 & n6060;
  assign n3891_1 = ~n5869_1;
  assign n5871 = n8259 | ~Ng1514;
  assign n5872 = Pg17423 & (n5871 | ~Ng1526);
  assign n5873 = Pg17320 & (Ng1526 | n5871);
  assign n5874_1 = Ng4709 | ~Ng4785;
  assign n5875 = n8208 | n8316;
  assign n5876 = Ng4674 & (n5874_1 | n5875 | ~Ng4743);
  assign n5877 = ~Ng3129 & ~Ng3143;
  assign n5878 = ~n8373 & (n5866 | (n5867 & ~Ng2803));
  assign n2738_1 = ~n5669;
  assign n5880 = Ng4420 | Ng4427;
  assign n5881 = Pg35 & (Ng6537 | Ng6523);
  assign n5882 = n8210 | n8317;
  assign n5883 = ~Ng4888 | Ng4899 | Ng4975;
  assign n5884_1 = Ng4836 & (n5882 | n5883);
  assign n5885 = Pg35 & (Ng6191 | Ng6177);
  assign n5886 = ~Ng1183 | n8288;
  assign n5887 = Pg17400 & (n5886 | ~Ng1171);
  assign n5888 = ~Ng4899 | Ng4975;
  assign n5889 = Ng4871 & (n5882 | n5888 | ~Ng4944);
  assign n2237_1 = ~n4252;
  assign n2890_1 = ~n4909;
  assign n5892 = n6075 & n6076 & n6077;
  assign n1349_1 = ~n5892;
  assign n5894 = Pg17316 & (Ng1171 | n5886);
  assign n5895 = n6033 & n6034 & n6035;
  assign n2511_1 = ~n5895;
  assign n5897 = n5970 | ~Ng4180;
  assign n5898_1 = ~n5997 & (n5897 | (Ng1105 & ~Ng947));
  assign n5899 = ~n8370 & (n5866 | (n5867 & ~Ng2783));
  assign n5648_1 = ~n5930;
  assign n5901 = n6273 & n6272 & n6271 & n6269 & n6266 & n6267 & n6268 & n6270_1;
  assign n5902 = Pg35 & (Ng3480 | Ng3494);
  assign n5903 = n6042_1 & n6039 & n6040 & n6041;
  assign n1586 = ~n5903;
  assign n5905 = Pg35 & (Ng5152 | Ng5138);
  assign n5906 = Pg35 & (Ng3845 | Ng3831);
  assign n5907 = Ng4899 | ~Ng4975;
  assign n5908 = Ng4864 & (n5882 | n5907 | ~Ng4933);
  assign n5909 = Ng1514 | n8259;
  assign n5910 = Pg17404 & (~Ng1526 | n5909);
  assign n5911 = Ng1430 & (Ng1526 | n5909);
  assign n5912 = n6050 & n6047 & n6048 & n6049;
  assign n4939 = ~n5912;
  assign n5914 = Ng1183 | n8288;
  assign n5915 = ~Ng4698 | Ng4709 | Ng4785;
  assign n5916 = ~n8255 & (n5866 | (n5867 & ~Ng2787));
  assign n4035_1 = ~n5929;
  assign n5918 = Pg35 & (Ng5499 | Ng5485);
  assign n5919 = ~n8370 & (n5866 | (n5867 & ~Ng2815));
  assign n5920 = ~n8255 & (n5866 | (n5867 & ~Ng2819));
  assign n5921 = Ng1087 & (Ng1171 | n5914);
  assign n5922 = n5971 | ~Ng4180;
  assign n5923 = ~n5999 & (n5922 | (Ng1300 & ~Ng1291));
  assign n5924 = ~Pg134 & (~Pg99 | ~Ng37);
  assign n5925 = ~n7957 & (n5866 | (n5867 & ~Ng2807));
  assign n5926 = ~Ng4899 | ~Ng4975;
  assign n5927 = Ng4878 & (n5882 | n5926 | ~Ng4955);
  assign n3802_1 = ~n5945;
  assign n5929 = n6123 & (n6124 | n6125 | n6126);
  assign n5930 = n6108 & n6106 & n6103 & n6104_1 & n6105 & n6107;
  assign n5931 = n8184 | n8185;
  assign n6497 = ~Pg35 & Ng2975;
  assign n5933 = Ng482 & ~Ng528 & Ng490;
  assign n5934 = ~n8469 & (Ng528 | n5933);
  assign n5935 = n5883 & n6136 & (n5907 | ~Ng4933);
  assign n5936 = n5935 & \[4651]  & \[4658]  & ~n5924;
  assign n2341_1 = ~n6122;
  assign n5938 = n6310_1 & n6309 & n6308 & n6306 & n6303 & n6304 & n6305 & n6307;
  assign n5939 = ~Ng4709 | Ng4785;
  assign n5940 = Ng4681 & (n5875 | n5939 | ~Ng4754);
  assign n5941 = ~n7957 & (n5866 | (n5867 & ~Ng2775));
  assign n5942 = ~n6001 & (n5922 | (Ng1472 & ~Ng1291));
  assign n3296_1 = ~n8177;
  assign n5944 = ~n6003 & (n5897 | (Ng956 & ~Ng947));
  assign n5945 = ~n6109 & (n6090 | (n6110 & n6111));
  assign n2027_1 = ~n9418;
  assign n5947 = n8226 | n8227;
  assign n5948 = ~n6005 & (n5897 | (Ng1129 & ~Ng947));
  assign n5949 = n5915 & n6135 & (n5939 | ~Ng4754);
  assign n5950 = n5949 & \[4651]  & \[4658]  & ~n5924;
  assign n5951 = ~Ng4709 | ~Ng4785;
  assign n5952 = Ng4688 & (n5875 | n5951 | ~Ng4765);
  assign n5953 = ~n6007 & (n5922 | (Ng1478 & ~Ng1291));
  assign n5954 = ~n6009 & (n5897 | (Ng1135 & ~Ng947));
  assign n6179 = ~Pg35 & Ng4392;
  assign n5956_1 = ~n6011 & (n5922 | (Ng1448 & ~Ng1291));
  assign n5957 = \[4436]  & (~Pg12368 | Pg9048);
  assign n5958 = n5963 & Pg7946 & (n5964 | n5965);
  assign n5959 = n7386 & Pg7916 & n8439;
  assign n5960 = ~Ng518 & ~Ng482 & ~n8181 & ~Ng499 & ~Ng528 & ~Ng490;
  assign n5961 = n9154 & (~Ng718 | ~Ng655 | ~Ng753);
  assign n5962 = n5960 & n5961 & (~Ng807 | ~Ng554);
  assign n5963 = Ng1339 & Ng1521 & ~Ng1532;
  assign n5964 = n8082 & Ng1367 & Ng1345 & Ng1379;
  assign n5965 = Ng1351 | Ng1312;
  assign n5966 = ~Pg113 & ~n5924;
  assign n5967 = Pg72 | Pg73;
  assign n5968 = Ng65 & (n5966 | n5967);
  assign n5969 = ~Ng691 | Ng209;
  assign n5970 = ~Pg134 & (n5969 | ~n6128);
  assign n5971 = ~Pg134 & (n5091 | n5969);
  assign n5972 = ~n4252 ^ n5912;
  assign n5973 = ~n5895 ^ n5903;
  assign n5974 = n4252 ^ n5912;
  assign n5975 = n5895 ^ n5903;
  assign n5976 = (n5972 | n5973) & (n5974 | n5975);
  assign n5977 = ~n4909 ^ n5669;
  assign n5978 = ~n5869_1 ^ n5892;
  assign n5979 = n4909 ^ n5669;
  assign n5980 = n5869_1 ^ n5892;
  assign n5981 = (n5977 | n5978) & (n5979 | n5980);
  assign n5982 = n7978 & n7979;
  assign n5983 = Ng225 | n8137;
  assign n5984 = ~n8137 | ~Ng225;
  assign n5985 = ~n9436 & (n5982 | (n5983 & n5984));
  assign n2498_1 = ~n5949;
  assign n6675 = ~n5935;
  assign n5988 = Ng2357 | Ng2491 | Ng2223 | Ng2472 | Ng2204 | Ng2625 | Ng2338 | Ng2606;
  assign n5989 = Ng2283 | Ng2685 | Ng2417 | Ng2537 | Ng2671 | Ng2551 | Ng2403 | Ng2269;
  assign n5990_1 = ~n6860 & (~Pg73 | Pg72);
  assign n5991 = ~n6860 & (Pg73 | ~Pg72);
  assign n5992 = ~Pg35 & (~n6015 | ~n8158);
  assign n5993 = Ng4578 & ~n6860;
  assign n5994 = ~Ng2756 | ~Ng2748 | ~Ng2735 | ~Ng2741;
  assign n5995 = n8198 & Pg35;
  assign n5996 = n5994 & n5995 & (Ng2756 | Ng2748);
  assign n5997 = ~n5970 & n6448 & (~Ng1105 | Ng947);
  assign n5998_1 = Pg35 & (n5898_1 | (~\[4421]  & n5997));
  assign n5999 = ~n5971 & n6336 & (~Ng1300 | Ng1291);
  assign n6000 = Pg35 & (n5923 | (n5999 & ~Ng1585));
  assign n6001 = ~n5971 & n6355 & (~Ng1472 | Ng1291);
  assign n6002 = Pg35 & (n5942 | (Ng1585 & n6001));
  assign n6003 = ~n5970 & n6410 & (~Ng956 | Ng947);
  assign n6004 = Pg35 & (n5944 | (~\[4421]  & n6003));
  assign n6005 = ~n5970 & n6429 & (~Ng1129 | Ng947);
  assign n6006 = Pg35 & (n5948 | (\[4421]  & n6005));
  assign n6007 = ~n5971 & n6391 & (~Ng1478 | Ng1291);
  assign n6008_1 = Pg35 & (n5953 | (n6007 & Ng1585));
  assign n6009 = ~n5970 & n6466 & (~Ng1135 | Ng947);
  assign n6010 = Pg35 & (n5954 | (n6009 & \[4421] ));
  assign n6011 = ~n5971 & n6373_1 & (~Ng1448 | Ng1291);
  assign n6012_1 = Pg35 & (n5956_1 | (~Ng1585 & n6011));
  assign n6013 = (n6027_1 | ~Ng758) & (~Ng586 | n8157);
  assign n6014 = ~n5992 & n9071 & (n6063 | ~Ng613);
  assign n6015 = n8147 | n8150;
  assign n6016 = n6013 & n6014 & (n6015 | ~Ng794);
  assign n6017_1 = (n6031 | ~Ng2950) & (n6056_1 | ~Ng2955);
  assign n6018 = n6036 & n9070 & (~Ng2868 | n8149);
  assign n6019 = n8151 | ~Ng51 | n8148;
  assign n6020 = n6017_1 & n6018 & (~Ng37 | n6019);
  assign n6021 = (Ng4927 | n8168) & (Ng4737 | n8169);
  assign n6022 = (~Ng947 | n8163) & (~Ng4300 | n8166);
  assign n6023 = (~Ng1291 | n8161) & (n6016 | n8142);
  assign n6024 = n9072 & (~Ng4172 | n8155);
  assign n6025 = (n6015 | ~Ng785) & (~Ng568 | n8157);
  assign n6026 = ~n5992 & n9079 & (~\[4426]  | n8159);
  assign n6027_1 = n8151 | ~Ng51 | n8150;
  assign n6028 = n6025 & n6026 & (n6027_1 | ~Ng744);
  assign n6029 = (~Pg92 | n6019) & (~Pg127 | n8149);
  assign n6030 = n9078 & (~Ng2975 | n6056_1);
  assign n6031 = ~n8144 | ~Ng51 | n8150;
  assign n6032 = n6029 & n6030 & (n6031 | ~Ng2970);
  assign n6033 = (n8155 | ~Ng4146) & (n8166 | ~Ng4249);
  assign n6034 = (n8173 | ~Ng2697) & (n6028 | n8142);
  assign n6035 = n9080 & n9081 & (n8163 | ~Ng939);
  assign n6036 = ~Ng51 | n8143 | ~n8144;
  assign n6037 = (n8149 | ~Ng2890) & (n8174 | ~Ng2984);
  assign n6038 = n6036 & n6037 & (~Pg100 | n6019);
  assign n6039 = (n8161 | ~Ng1287) & (n8163 | ~Ng943);
  assign n6040 = (n8166 | ~Ng4245) & (n8171 | ~Ng2145);
  assign n6041 = (n8155 | ~Ng4157) & (n8173 | ~Ng2704);
  assign n6042_1 = n9086 & (n8142 | (n9085 & n9083));
  assign n6043 = (n6031 | ~Ng2960) & (n6056_1 | ~Ng2965);
  assign n6044 = (n8149 | ~Ng2873) & (~\[4433]  | n6019);
  assign n6045 = n8150 | ~Ng48 | n8146;
  assign n6046 = n6043 & n6044 & (n6045 | ~Ng2878);
  assign n6047 = (~Ng2689 | n8173) & (n8163 | Ng952);
  assign n6048 = (n8155 | ~Ng4176) & (~Ng2130 | n8171);
  assign n6049 = (n8161 | Ng1296) & (n8166 | ~Ng4253);
  assign n6050 = n9077 & (n8142 | (n9076 & n9074));
  assign n6051 = (n8159 | ~Ng546) & (~Ng582 | n8157);
  assign n6052 = ~n5992 & n9093 & (n6063 | ~Ng622);
  assign n6053 = n6051 & n6052 & (n6027_1 | ~Ng767);
  assign n6054 = (n6045 | ~Ng2864) & (n6080 | ~Ng2860);
  assign n6055 = (n6031 | ~Ng2922) & (n8149 | Ng2994);
  assign n6056_1 = n8150 | ~n8144 | Ng51;
  assign n6057 = n6054 & n6055 & (n6056_1 | ~Ng2927);
  assign n6058 = (n8168 | ~Ng4907) & (n8173 | ~Ng3151);
  assign n6059 = (n8169 | ~Ng4717) & (n6053 | n8142);
  assign n6060 = n9094 & n9095 & (n6057 | n8142);
  assign n6061_1 = (~Ng595 | n8157) & (Pg35 | n8158);
  assign n6062 = (n8159 | ~Ng538) & (n6027_1 | ~Ng776);
  assign n6063 = n8143 | n8156;
  assign n6064 = n6061_1 & n6062 & (n6063 | ~Ng632);
  assign n6065 = (n8169 | ~Ng4727) & (n8171 | ~Ng6199);
  assign n6066 = (n8168 | ~Ng4917) & (n8173 | ~Ng3853);
  assign n6067 = (n8153 | ~Ng45) & (n6064 | n8142);
  assign n6068 = n9089 & (n8142 | (n9088 & n9087));
  assign n6069 = (n6015 | ~Ng807) & (~Ng577 | n8157);
  assign n6070 = ~n5992 & n9097 & (n8159 | ~Ng542);
  assign n6071 = n6069 & n6070 & (n6027_1 | ~Ng763);
  assign n6072 = (n6031 | ~Ng2936) & (n6080 | ~Ng2894);
  assign n6073 = n6036 & n9096 & (n8149 | ~Ng2988);
  assign n6074 = n6072 & n6073 & (n6056_1 | ~Ng2941);
  assign n6075 = (n8169 | ~Ng4722) & (n6071 | n8142);
  assign n6076 = (n8171 | ~Ng5160) & (n8173 | ~Ng6545);
  assign n6077 = n9098 & n9099 & (n6074 | n8142);
  assign n6078 = (n6045 | ~Ng2856) & (n6056_1 | ~Ng2917);
  assign n6079 = (n6031 | ~Ng2912) & (n8149 | ~Ng2999);
  assign n6080 = n8154 | ~Ng48 | n8150;
  assign n6081_1 = n6078 & n6079 & (n6080 | ~Ng2852);
  assign n6082 = (n8168 | ~Ng4922) & (n8173 | ~Ng3502);
  assign n6083 = (n8169 | ~Ng4732) & (n8171 | ~Ng5853);
  assign n6084 = (n8153 | ~Ng46) & (n6081_1 | n8142);
  assign n6085 = n9092 & (n8142 | (n9091 & n9090));
  assign n6086 = n5981 ^ n5976;
  assign n6087 = n6086 & (~Ng55 | (~Pg56 & Pg54));
  assign n6088 = ~n6086 & Ng55 & (Pg56 | ~Pg54);
  assign n6089 = ~n8177 & ~Pg53 & ~Pg56 & ~Pg54;
  assign n6090 = n8179 | Ng4311 | n8178;
  assign n6091_1 = n5962 & (~Pg12184 | Pg11678);
  assign n6092 = (n7743 | ~Ng554) & (Pg35 | ~Ng807);
  assign n6093 = ~Ng794 | n6114;
  assign n6094 = n9158 & (Ng4584 | ~Ng4608 | Ng4593);
  assign n6095 = Ng4584 ^ Ng4608;
  assign n6096_1 = Ng4601 ^ Ng4593;
  assign n6097 = n6094 & (Ng4616 | n6095 | n6096_1);
  assign n6098 = ~n6093 | ~Ng807 | n7743;
  assign n6099 = Pg35 | ~Ng794;
  assign n6100 = ~Ng632 | ~n6102 | n8183;
  assign n6101 = Pg35 | ~Ng626;
  assign n6102 = ~Ng626 | n6117;
  assign n6103 = n8068 | n6269;
  assign n6104_1 = ~Ng2070 | n6267 | Ng2040;
  assign n6105 = ~Ng1936 | n6272 | Ng1906;
  assign n6106 = ~Ng2227 | n6271 | Ng2197;
  assign n6107 = (n8078 | n6266) & (n8080 | n6268);
  assign n6108 = (n8070 | n6270_1) & (n8066 | n6273);
  assign n6109 = ~n6124 & (~n9100 | ~n9101);
  assign n6110 = (n5730 | n7445) & (n8191 | n8192);
  assign n6111 = (n8188 | n7507) & (n8190 | n7476);
  assign n6112 = ~Ng794 | ~n6114 | n7743;
  assign n6113 = Pg35 | ~Ng790;
  assign n6114 = ~Ng790 | n6131;
  assign n6115 = ~Ng626 | ~n6117 | n8183;
  assign n6116 = Pg35 | ~Ng622;
  assign n6117 = ~Ng622 | n6134;
  assign n6118 = (n8205 | n6306) & (n8207 | n6310_1);
  assign n6119 = (n8203 | n6303) & (n8204 | n6305);
  assign n6120 = (n8201 | n6309) & (n8202 | n6308);
  assign n6121 = (n8197 | n6307) & (n8199 | n6304);
  assign n6122 = n6121 & n6118 & n6119 & n6120;
  assign n6123 = n8065 | n6090 | n7796;
  assign n6124 = n8179 | ~Ng4311 | n8178;
  assign n6125 = n5926 | n8211;
  assign n6126 = ~Ng4878 | n8210;
  assign n6127_1 = Ng2389 | Ng2657 | Ng2523 | Ng2255;
  assign n6128 = Ng1193 & (Ng969 | Ng1008);
  assign n6129 = ~Ng790 | ~n6131 | n7743;
  assign n6130 = Pg35 | ~Ng785;
  assign n6131 = ~Ng785 | n6148;
  assign n6132 = ~Ng622 | ~n6134 | n8183;
  assign n6133 = Pg35 | ~Ng617;
  assign n6134 = ~Ng617 | n6151;
  assign n6135 = (n5874_1 | ~Ng4743) & (n5951 | ~Ng4765);
  assign n6136 = (n5888 | ~Ng4944) & (n5926 | ~Ng4955);
  assign n6137_1 = ~Pg35 | ~Ng2994;
  assign n6138 = (~Pg35 | ~Ng1287) & ~n8478;
  assign n6139 = Pg35 | ~Ng1283;
  assign n6140 = n4219 & (~Pg35 | ~Ng1296);
  assign n6141 = Pg35 | ~Ng1291;
  assign n6142_1 = n4217 & (~Pg35 | ~Ng943);
  assign n6143 = Pg35 | ~Ng939;
  assign n6144 = n4218 & (~Pg35 | ~Ng952);
  assign n6145 = Pg35 | ~Ng947;
  assign n6146 = ~Ng785 | ~n6148 | n7743;
  assign n6147_1 = Pg35 | ~Ng781;
  assign n6148 = ~Ng781 | n6186;
  assign n6149 = ~Ng617 | ~n6151 | n8183;
  assign n6150 = Pg35 | ~Ng613;
  assign n6151 = ~Ng613 | n6189;
  assign n6152_1 = ~Pg35 | ~Ng4927;
  assign n6153 = ~Pg35 | ~Ng4912;
  assign n6154 = ~Pg35 | ~Ng4907;
  assign n6155 = ~Pg35 | ~Ng4922;
  assign n6156_1 = ~Pg35 | ~Ng4737;
  assign n6157 = ~Pg35 | ~Ng4722;
  assign n6158 = ~Pg35 | ~Ng4717;
  assign n6159 = ~Pg35 | ~Ng4732;
  assign n6160_1 = ~Pg35 | ~Ng4245;
  assign n6161 = ~Pg35 | ~Ng4249;
  assign n6162 = ~Pg35 | ~Ng4253;
  assign n6163 = ~Pg35 | ~Ng4157;
  assign n6164 = ~Pg35 | ~Ng4146;
  assign n6165_1 = ~Pg35 | ~Ng2988;
  assign n6166 = ~Pg35 | ~Ng2970;
  assign n6167 = ~Pg35 | ~Ng2960;
  assign n6168 = ~Pg35 | ~Ng2950;
  assign n6169_1 = ~Pg35 | ~Ng2936;
  assign n6170 = ~Pg35 | ~Ng2922;
  assign n6171 = ~Pg35 | ~Ng2912;
  assign n6172 = ~Pg35 | ~Ng2907;
  assign n6173 = ~Pg35 | ~Ng2868;
  assign n6174 = ~Pg35 | ~Ng2873;
  assign n6175 = (~Pg35 | ~Ng37) & n9187;
  assign n6176 = ~Pg35 | ~Ng2894;
  assign n6177 = ~Pg35 | ~Ng2860;
  assign n6178 = ~Pg35 | ~Ng2852;
  assign n6179_1 = ~Pg35 | ~Ng2844;
  assign n6180 = ~Pg35 | ~Ng2704;
  assign n6181 = ~Pg35 | ~Ng2697;
  assign n6182 = ~Pg35 | ~Ng2145;
  assign n6183_1 = ~Pg35 | ~Ng2138;
  assign n6184 = ~Ng781 | ~n6186 | n7743;
  assign n6185 = Pg35 | ~Ng776;
  assign n6186 = ~Ng776 | n6257;
  assign n6187 = ~Ng613 | ~n6189 | n8183;
  assign n6188 = Pg35 | ~Ng608;
  assign n6189 = ~Ng608 | n6259;
  assign n6190 = (Pg35 | ~Ng4854) & (n6193 | ~Ng4859);
  assign n6191 = ~Ng4849 | n8229;
  assign n6192_1 = n6191 ^ Ng4854;
  assign n6193 = ~Pg35 | ~n8228;
  assign n6194 = n8229 | Ng4849 | ~n8228;
  assign n6195 = (Pg35 | ~Ng4664) & (n6198 | ~Ng4669);
  assign n6196_1 = ~Ng4659 | n8231;
  assign n6197 = n6196_1 ^ Ng4664;
  assign n6198 = ~Pg35 | ~n8230;
  assign n6199 = n8231 | Ng4659 | ~n8230;
  assign n6200 = n5968 | Ng4643;
  assign n6201 = Pg35 & (Ng4621 | n6200);
  assign n6202 = Ng4639 | n6205;
  assign n6203 = ~n5968 & (~Ng4621 | Ng4639 | ~Ng4628);
  assign n6204 = ~n5968 & Ng4340;
  assign n6205 = ~Pg35 | n6200;
  assign n6206_1 = n6202 & (Ng4621 | n6205);
  assign n6207 = n6206_1 & (Ng4628 | n6205);
  assign n6208 = ~Ng4621 | n6200;
  assign n6209 = Pg35 & (Ng4633 | ~Ng4639 | n6208);
  assign n6210 = n6208 | ~Ng4639 | Ng4628;
  assign n6211_1 = Pg35 | ~Ng4621;
  assign n6212 = ~n5968 & (~Ng4616 | ~n8234);
  assign n6213 = (~Ng4616 | n6220) & (Pg35 | ~Ng4608);
  assign n6214 = ~Ng4601 | n8061;
  assign n6215 = (Pg35 | ~Ng4322) & (~Ng4332 | n8235);
  assign n6216_1 = n5968 | n8062;
  assign n6217 = ~Ng4608 | ~n6214 | n6220;
  assign n6218 = Ng4608 | ~n6212 | n6214;
  assign n6219 = Ng4601 ^ n8061;
  assign n6220 = ~Pg35 | ~n6212;
  assign n6221_1 = n8234 | n6220 | ~Ng4593;
  assign n6222 = ~n8234 | ~n6212 | Ng4593;
  assign n6223 = ~n8062 ^ Ng4584;
  assign n6224 = n8236 | ~Ng4322 | n8235;
  assign n6225 = ~n8236 | n6216_1 | Ng4322;
  assign n6226_1 = ~n8329 & (~Pg35 | Ng2827);
  assign n6227 = n9193 & (~Pg35 | ~n6229 | ~Ng2819);
  assign n6228 = n5966 & Ng111;
  assign n6229 = ~Ng2729 | n5994 | ~Ng2724;
  assign n6230_1 = ~n8329 & (~Pg35 | Ng2811);
  assign n6231 = n9194 & (~Pg35 | ~n6232 | ~Ng2807);
  assign n6232 = Ng2729 | n5994 | ~Ng2724;
  assign n6233 = ~n8329 & (~Pg35 | Ng2823);
  assign n6234 = n9195 & (~Pg35 | ~n6235_1 | ~Ng2815);
  assign n6235_1 = ~Ng2729 | n5994 | Ng2724;
  assign n6236 = ~n8329 & (~Pg35 | Ng2799);
  assign n6237 = n9196 & (~Pg35 | ~n6238 | ~Ng2803);
  assign n6238 = n5994 | n5866;
  assign n6239 = ~n8329 & (~Pg35 | Ng2795);
  assign n6240_1 = n9197 & (~Pg35 | ~n6229 | ~Ng2787);
  assign n6241 = n5966 & Ng85;
  assign n6242 = ~n8329 & (~Pg35 | Ng2779);
  assign n6243 = n9198 & (~Pg35 | ~n6232 | ~Ng2775);
  assign n6244 = ~n8329 & (~Pg35 | Ng2791);
  assign n6245_1 = n9199 & (~Pg35 | ~n6235_1 | ~Ng2783);
  assign n6246 = ~n8329 & (~Pg35 | Ng2767);
  assign n6247 = n9200 & (~Pg35 | ~n6238 | ~Ng2771);
  assign n6248 = ~Ng182 ^ n9201;
  assign n6249 = (Ng392 & ~Ng441) | (~Ng411 & (~Ng392 | ~Ng441));
  assign n6250_1 = ~Ng417 & n6248 & n6249 & ~Ng691;
  assign n6251 = ~Ng703 & ~n5049 & n5050;
  assign n6252 = Ng376 & Ng385 & Pg8719;
  assign n6253 = Ng896 & (n6252 | n6251);
  assign n6254 = (~Ng890 | ~Ng896) & (n6253 | ~Ng862);
  assign n6255_1 = ~Ng776 | ~n6257 | n7743;
  assign n6256 = Pg35 | ~Ng772;
  assign n6257 = ~Ng772 | n6295;
  assign n6258 = Pg35 | ~Ng604;
  assign n6259 = ~Ng604 | n6297_1;
  assign n6260_1 = ~Ng4141 & ~Ng4082;
  assign n6261 = Ng4093 | Ng4098;
  assign n6262 = ~Ng4076 | ~Ng4112;
  assign n6263 = n6260_1 & (Ng4087 | n6261 | n6262);
  assign n6264 = Pg113 & ~n5924;
  assign n6265_1 = (~n6090 | ~n6124) & n6264;
  assign n6266 = ~Ng504 | Ng528 | n8186;
  assign n6267 = n8187 | Ng504 | Ng528;
  assign n6268 = n8186 | Ng504 | Ng528;
  assign n6269 = ~Ng528 | ~Ng504 | n8187;
  assign n6270_1 = ~Ng504 | ~Ng528 | n8186;
  assign n6271 = Ng504 | ~Ng528 | n8186;
  assign n6272 = n8187 | Ng528 | ~Ng504;
  assign n6273 = n8187 | ~Ng528 | Ng504;
  assign n6274 = (~Ng4961 | ~n8237) & ~n8238;
  assign n6275_1 = (~n8237 | ~Ng4950) & ~n8238;
  assign n6276 = (~Pg35 | ~n8238) & (~n8237 | ~Ng4939);
  assign n6277 = Pg35 | ~Ng4939;
  assign n6278 = ~Pg35 | ~n6279_1 | ~Ng4933;
  assign n6279_1 = n7774 & n8237;
  assign n6280 = ~n8238 & (~n8237 | ~Ng4894);
  assign n6281 = n8239 | ~Ng101;
  assign n6282 = n6281 & (~Ng4771 | ~n8239);
  assign n6283 = n6281 & (~n8239 | ~Ng4760);
  assign n6284_1 = (~Pg35 | n6281) & (~n8239 | ~Ng4749);
  assign n6285 = Pg35 | ~Ng4749;
  assign n6286 = ~Pg35 | ~n6287 | ~Ng4743;
  assign n6287 = n7790 & n8239;
  assign n6288 = n6281 & (~n8239 | ~Ng4704);
  assign n6289_1 = ~n5967 & (n5924 | Ng4507);
  assign n6290 = ~Ng26960 | n6289_1 | Ng4477;
  assign n6291 = n6290 & ~Ng4459 & (Ng4462 | ~Ng4473);
  assign n6292 = Ng4643 & Pg35 & Ng4462 & ~Ng10384;
  assign n6293_1 = ~Ng772 | ~n6295 | n7743;
  assign n6294 = Pg35 | ~Ng767;
  assign n6295 = ~Ng767 | n6488;
  assign n6296 = Pg35 | ~Ng599;
  assign n6297_1 = ~Ng599 | n6490;
  assign n6298 = Ng142 | n8245;
  assign n6299 = ~Ng142 | n7834 | ~n8245;
  assign n6300 = n4520 & (Ng182 | Ng174 | Ng168);
  assign n6301 = Ng160 | n9218;
  assign n6302_1 = ~n9218 | ~Ng160 | n7402;
  assign n6303 = n8200 | ~Ng2756 | Ng2741;
  assign n6304 = n8195 | n8198;
  assign n6305 = ~Ng2741 | n8196;
  assign n6306 = ~Ng2756 | ~Ng2741 | n8200;
  assign n6307 = Ng2741 | n8196;
  assign n6308 = n8200 | Ng2741 | Ng2756;
  assign n6309 = n8200 | Ng2756 | ~Ng2741;
  assign n6310_1 = n8195 | ~n8206;
  assign n6311 = n6126 ^ Ng4983;
  assign n6312 = ~Pg35 | n6317;
  assign n6313 = (n5907 | ~n8252) & (~Pg35 | n5888);
  assign n6314 = (n6312 | ~Ng4899) & (n6313 | n8251);
  assign n6315_1 = (Pg35 | ~Ng4991) & (n6312 | ~Ng4966);
  assign n6316 = n6126 | ~Ng4983;
  assign n6317 = n8251 | n8252;
  assign n6318 = n6316 | Ng4991 | n6317;
  assign n6319 = ~Ng4991 | n6312 | ~n6316;
  assign n6320_1 = ~n8252 | Ng4975 | n8251;
  assign n6321 = Pg35 | ~Ng4966;
  assign n6322 = n8065 ^ Ng4793;
  assign n6323 = ~Pg35 | n6328;
  assign n6324 = (~Pg35 | n5939) & (n5874_1 | ~n8254);
  assign n6325 = (n6323 | ~Ng4709) & (n6324 | n8253);
  assign n6326 = (Pg35 | ~Ng4801) & (n6323 | ~Ng4776);
  assign n6327 = n8065 | ~Ng4793;
  assign n6328 = n8253 | n8254;
  assign n6329 = n6327 | Ng4801 | n6328;
  assign n6330_1 = ~Ng4801 | n6323 | ~n6327;
  assign n6331 = ~n8254 | Ng4785 | n8253;
  assign n6332 = Pg35 | ~Ng4776;
  assign n6333 = ~Pg35 | Ng2841;
  assign n6334 = n9223 & (~Pg35 | ~Ng2763 | ~n6335_1);
  assign n6335_1 = ~Ng2759 | n6542;
  assign n6336 = ~Ng2689 | ~Ng2697 | ~Ng2704;
  assign n6337 = (~n6000 | n8261) & (~n8262 | ~Ng2567);
  assign n6338 = ~n5923 & (~n5999 | Ng1589);
  assign n6339 = (Pg35 & ~n8648) | (~Ng2629 & (~Pg35 | ~n8648));
  assign n6340_1 = ~Pg35 | n8263;
  assign n6341 = Pg35 | ~Ng2571;
  assign n6342 = ~Pg35 | ~n6343 | ~Ng2583;
  assign n6343 = n8066 | ~n8263;
  assign n6344 = Pg35 | ~Ng2583;
  assign n6345 = ~Pg35 | ~Ng2579 | n8265;
  assign n6346 = Pg35 | ~Ng2579;
  assign n6347 = ~Pg35 | ~n6348 | ~Ng2575;
  assign n6348 = ~Ng2629 | n8266;
  assign n6349_1 = Pg35 | ~Ng2563;
  assign n6350 = ~Pg35 | ~n6351 | ~Ng2571;
  assign n6351 = ~n8263 | ~Ng2599 | Ng2629;
  assign n6352 = Pg35 | ~Ng2567;
  assign n6353 = ~Pg35 | ~n6354_1 | ~Ng2563;
  assign n6354_1 = Ng2599 | n8266;
  assign n6355 = ~Ng2689 | ~Ng2697 | Ng2704;
  assign n6356 = (~n6002 | n8268) & (~n8269 | ~Ng2433);
  assign n6357 = ~n5942 & (~n6001 | ~Ng1589);
  assign n6358 = (Pg35 & ~n8650) | (~Ng2495 & (~Pg35 | ~n8650));
  assign n6359_1 = ~Pg35 | n8270;
  assign n6360 = Pg35 | ~Ng2437;
  assign n6361 = n8068 | ~n8270;
  assign n6362 = Pg35 | ~Ng2449;
  assign n6363 = ~Pg35 | ~Ng2445 | n8272;
  assign n6364 = Pg35 | ~Ng2445;
  assign n6365 = ~Pg35 | ~n6366 | ~Ng2441;
  assign n6366 = ~Ng2495 | n8273;
  assign n6367 = Pg35 | ~Ng2429;
  assign n6368 = ~Pg35 | ~n6369_1 | ~Ng2437;
  assign n6369_1 = ~n8270 | ~Ng2465 | Ng2495;
  assign n6370 = Pg35 | ~Ng2433;
  assign n6371 = ~Pg35 | ~n6372 | ~Ng2429;
  assign n6372 = Ng2465 | n8273;
  assign n6373_1 = ~Ng2704 | ~Ng2689 | Ng2697;
  assign n6374 = (~n6012_1 | n8275) & (~n8276 | ~Ng2299);
  assign n6375 = ~n5956_1 & (~n6011 | Ng1589);
  assign n6376_1 = (Pg35 & ~n8652) | (~Ng2361 & (~Pg35 | ~n8652));
  assign n6377 = ~Pg35 | n8277;
  assign n6378 = Pg35 | ~Ng2303;
  assign n6379 = n8070 | ~n8277;
  assign n6380_1 = Pg35 | ~Ng2315;
  assign n6381 = ~Pg35 | ~Ng2311 | n8279;
  assign n6382 = Pg35 | ~Ng2311;
  assign n6383 = ~Pg35 | ~n6384 | ~Ng2307;
  assign n6384 = ~Ng2361 | n8280;
  assign n6385_1 = Pg35 | ~Ng2295;
  assign n6386 = ~Pg35 | ~n6387 | ~Ng2303;
  assign n6387 = ~n8277 | ~Ng2331 | Ng2361;
  assign n6388 = Pg35 | ~Ng2299;
  assign n6389 = ~Pg35 | ~n6390_1 | ~Ng2295;
  assign n6390_1 = Ng2331 | n8280;
  assign n6391 = Ng2704 | ~Ng2689 | Ng2697;
  assign n6392 = (~n6008_1 | n8282) & (~n8283 | ~Ng2165);
  assign n6393 = ~n5953 & (~n6007 | ~Ng1589);
  assign n6394 = (Pg35 & ~n8654) | (~Ng2227 & (~Pg35 | ~n8654));
  assign n6395_1 = ~Pg35 | n8284;
  assign n6396 = Pg35 | ~Ng2169;
  assign n6397 = ~Pg35 | ~n6398 | ~Ng2181;
  assign n6398 = Ng2197 | n8285;
  assign n6399_1 = Pg35 | ~Ng2181;
  assign n6400 = ~Pg35 | ~Ng2177 | n8287;
  assign n6401 = Pg35 | ~Ng2177;
  assign n6402 = ~Pg35 | ~n6403_1 | ~Ng2173;
  assign n6403_1 = n8285 | ~Ng2153;
  assign n6404 = Pg35 | ~Ng2161;
  assign n6405 = ~Pg35 | ~n6406 | ~Ng2169;
  assign n6406 = ~n8284 | ~Ng2197 | Ng2227;
  assign n6407 = Pg35 | ~Ng2165;
  assign n6408 = ~Pg35 | ~n6409 | ~Ng2161;
  assign n6409 = ~Ng2153 | Ng2197 | ~n8284;
  assign n6410 = ~Ng2130 | ~Ng2138 | ~Ng2145;
  assign n6411 = (~n6004 | n8290) & (~n8291 | ~Ng2008);
  assign n6412 = ~n5944 & (~n6003 | Ng1246);
  assign n6413_1 = (Pg35 & ~n8656) | (~Ng2070 & (~Pg35 | ~n8656));
  assign n6414 = ~Pg35 | n8292;
  assign n6415 = Pg35 | ~Ng2012;
  assign n6416 = ~Pg35 | ~n6417_1 | ~Ng2024;
  assign n6417_1 = Ng2040 | n8293;
  assign n6418 = Pg35 | ~Ng2024;
  assign n6419 = ~Pg35 | ~Ng2020 | n8295;
  assign n6420 = Pg35 | ~Ng2020;
  assign n6421 = ~Pg35 | ~n6422_1 | ~Ng2016;
  assign n6422_1 = n8293 | ~Ng1996;
  assign n6423 = Pg35 | ~Ng2004;
  assign n6424 = ~Pg35 | ~n6425 | ~Ng2012;
  assign n6425 = ~n8292 | ~Ng2040 | Ng2070;
  assign n6426 = Pg35 | ~Ng2008;
  assign n6427_1 = ~Pg35 | ~n6428 | ~Ng2004;
  assign n6428 = ~Ng1996 | Ng2040 | ~n8292;
  assign n6429 = ~Ng2130 | ~Ng2138 | Ng2145;
  assign n6430 = (~n6006 | n8297) & (~n8298 | ~Ng1874);
  assign n6431 = ~n5948 & (~n6005 | ~Ng1246);
  assign n6432_1 = (Pg35 & ~n8658) | (~Ng1936 & (~Pg35 | ~n8658));
  assign n6433 = ~Pg35 | n8299;
  assign n6434 = Pg35 | ~Ng1878;
  assign n6435 = ~Pg35 | ~n6436 | ~Ng1890;
  assign n6436 = Ng1906 | n8300;
  assign n6437_1 = Pg35 | ~Ng1890;
  assign n6438 = ~Pg35 | ~Ng1886 | n8302;
  assign n6439 = Pg35 | ~Ng1886;
  assign n6440 = ~Pg35 | ~n6441 | ~Ng1882;
  assign n6441 = n8300 | ~Ng1862;
  assign n6442_1 = Pg35 | ~Ng1870;
  assign n6443 = ~Pg35 | ~n6444 | ~Ng1878;
  assign n6444 = ~n8299 | ~Ng1906 | Ng1936;
  assign n6445 = Pg35 | ~Ng1874;
  assign n6446 = ~Pg35 | ~n6447_1 | ~Ng1870;
  assign n6447_1 = ~Ng1862 | Ng1906 | ~n8299;
  assign n6448 = ~Ng2145 | ~Ng2130 | Ng2138;
  assign n6449 = (~n5998_1 | n8304) & (~n8305 | ~Ng1740);
  assign n6450 = ~n5898_1 & (~n5997 | Ng1246);
  assign n6451 = (Pg35 & ~n8660) | (~Ng1802 & (~Pg35 | ~n8660));
  assign n6452_1 = ~Pg35 | n8306;
  assign n6453 = Pg35 | ~Ng1744;
  assign n6454 = n8078 | ~n8306;
  assign n6455 = Pg35 | ~Ng1756;
  assign n6456 = ~Pg35 | ~Ng1752 | n8308;
  assign n6457_1 = Pg35 | ~Ng1752;
  assign n6458 = ~Pg35 | ~n6459 | ~Ng1748;
  assign n6459 = ~Ng1802 | n8309;
  assign n6460 = Pg35 | ~Ng1736;
  assign n6461 = ~Pg35 | ~n6462_1 | ~Ng1744;
  assign n6462_1 = ~n8306 | ~Ng1772 | Ng1802;
  assign n6463 = Pg35 | ~Ng1740;
  assign n6464 = ~Pg35 | ~n6465 | ~Ng1736;
  assign n6465 = Ng1772 | n8309;
  assign n6466 = Ng2145 | ~Ng2130 | Ng2138;
  assign n6467_1 = (~n6010 | n8311) & (~n8312 | ~Ng1604);
  assign n6468 = ~n5954 & (~n6009 | ~Ng1246);
  assign n6469 = (Pg35 & ~n8662) | (~Ng1668 & (~Pg35 | ~n8662));
  assign n6470 = ~Pg35 | n8313;
  assign n6471 = Pg35 | ~Ng1608;
  assign n6472_1 = ~Pg35 | ~n6473 | ~Ng1620;
  assign n6473 = n8080 | ~n8313;
  assign n6474 = Pg35 | ~Ng1620;
  assign n6475 = ~Pg35 | ~n6476 | ~Ng1616;
  assign n6476 = Ng1592 | n8314;
  assign n6477_1 = Pg35 | ~Ng1616;
  assign n6478 = ~Pg35 | ~n6479 | ~Ng1612;
  assign n6479 = ~Ng1668 | n8315;
  assign n6480 = Pg35 | ~Ng1600;
  assign n6481 = ~Pg35 | ~n6482_1 | ~Ng1608;
  assign n6482_1 = Ng1668 | n8314;
  assign n6483 = Pg35 | ~Ng1604;
  assign n6484 = ~Pg35 | ~n6485 | ~Ng1600;
  assign n6485 = Ng1636 | n8315;
  assign n6486 = ~Ng767 | ~n6488 | n7743;
  assign n6487_1 = Pg35 | ~Ng763;
  assign n6488 = ~Ng763 | n6647;
  assign n6489 = Pg35 | ~Ng595;
  assign n6490 = ~Ng595 | n6649;
  assign n6491 = Ng298 | n8244;
  assign n6492_1 = ~n8244 | n7834 | ~Ng298;
  assign n6493 = Ng157 | n8250;
  assign n6494 = ~n8250 | n7402 | ~Ng157;
  assign n6495 = (~Pg35 | n7426) & (n6500 | ~Ng6682);
  assign n6496 = ~Ng6741 | Ng6682;
  assign n6497_1 = n6495 & (~n5884_1 | n6496);
  assign n6498 = Pg35 | ~Ng6736;
  assign n6499 = ~Pg35 | ~n5884_1 | Ng6741 | ~n9420;
  assign n6500 = ~Pg35 | n5884_1;
  assign n6501 = (~Pg35 | n7454) & (n6506 | ~Ng6336);
  assign n6502_1 = ~Ng6395 | Ng6336;
  assign n6503 = n6501 & (~n5952 | n6502_1);
  assign n6504 = Pg35 | ~Ng6390;
  assign n6505 = ~Pg35 | ~n5952 | Ng6395 | ~n9421;
  assign n6506 = ~Pg35 | n5952;
  assign n6507_1 = (~Pg35 | n7488) & (n6512_1 | ~Ng5990);
  assign n6508 = ~Ng6049 | Ng5990;
  assign n6509 = n6507_1 & (~n5940 | n6508);
  assign n6510 = Pg35 | ~Ng6044;
  assign n6511 = ~Pg35 | ~n5940 | Ng6049 | ~n9423;
  assign n6512_1 = ~Pg35 | n5940;
  assign n6513 = n7791 | ~Ng5703;
  assign n6514 = ~n9224 | Ng5703 | n8322;
  assign n6515 = (~Pg35 | n7548) & (n6520 | ~Ng5297);
  assign n6516 = ~Ng5357 | Ng5297;
  assign n6517_1 = n6515 & (~n4151_1 | n6516);
  assign n6518 = Pg35 | ~Ng5352;
  assign n6519 = ~Pg35 | ~n4151_1 | Ng5357 | ~n9422;
  assign n6520 = ~Pg35 | n4151_1;
  assign n6521 = ~Pg35 | Ng2841;
  assign n6522_1 = n9226 & (~Pg35 | ~Ng4104 | ~n6523);
  assign n6523 = ~Ng4108 | n6712;
  assign n6524 = (~Pg35 | n7590) & (n6529 | ~Ng3990);
  assign n6525 = ~Ng4054 | Ng3990;
  assign n6526_1 = n6524 & (~n5927 | n6525);
  assign n6527 = Pg35 | ~Ng4049;
  assign n6528 = ~Pg35 | ~n5927 | Ng4054 | ~n9419;
  assign n6529 = ~Pg35 | n5927;
  assign n6530 = (~Pg35 | n8327) & (n6535 | ~Ng3639);
  assign n6531_1 = ~Ng3703 | Ng3639;
  assign n6532 = n6530 & (~n5889 | n6531_1);
  assign n6533 = Pg35 | ~Ng3698;
  assign n6534 = ~Pg35 | ~n5889 | Ng3703 | ~n9424;
  assign n6535 = ~Pg35 | n5889;
  assign n6536_1 = (n7775 | ~Ng3288) & (~Pg35 | n7638);
  assign n6537 = ~Ng3352 | Ng3288;
  assign n6538 = n6536_1 & (~n5908 | n6537);
  assign n6539 = n7775 | ~Ng3352;
  assign n6540 = ~n9425 | Ng3352 | n8328;
  assign n6541_1 = n9227 & (~Pg35 | ~Ng2759 | ~n6542);
  assign n6542 = ~Ng2756 | n8258;
  assign n6543 = ~Pg35 | n5966;
  assign n6544 = n6543 & (~Pg35 | (n5911 & ~n6273));
  assign n6545 = Pg35 | ~Ng2555;
  assign n6546_1 = Pg35 | ~Ng2671;
  assign n6547 = Ng2675 | ~Pg35 | n8261;
  assign n6548 = (~Ng2671 | ~n8262) & (n8261 | ~n8680);
  assign n6549 = ~n6273 & n8330;
  assign n6550 = Pg35 & (n6549 | ~n8263);
  assign n6551_1 = n8266 | ~Pg35 | n6549;
  assign n6552 = Pg35 | ~Ng2606;
  assign n6553 = ~Ng2555 & (Ng2599 | ~n8263);
  assign n6554 = ~Pg35 | n6549 | n6553 | Ng2629;
  assign n6555_1 = n6543 & (~Pg35 | (n5872 & ~n6269));
  assign n6556 = Pg35 | ~Ng2421;
  assign n6557 = Pg35 | ~Ng2537;
  assign n6558 = Ng2541 | ~Pg35 | n8268;
  assign n6559 = (~Ng2537 | ~n8269) & (n8268 | ~n8685);
  assign n6560_1 = ~n6269 & n8330;
  assign n6561 = Pg35 & (n6560_1 | ~n8270);
  assign n6562 = n8273 | ~Pg35 | n6560_1;
  assign n6563 = Pg35 | ~Ng2472;
  assign n6564 = ~Ng2421 & (Ng2465 | ~n8270);
  assign n6565_1 = ~Pg35 | n6560_1 | n6564 | Ng2495;
  assign n6566 = n6543 & (~Pg35 | (n5910 & ~n6270_1));
  assign n6567 = Pg35 | ~Ng2287;
  assign n6568 = Pg35 | ~Ng2403;
  assign n6569 = Ng2407 | ~Pg35 | n8275;
  assign n6570_1 = (~Ng2403 | ~n8276) & (n8275 | ~n8690);
  assign n6571 = ~n6270_1 & n8330;
  assign n6572 = Pg35 & (n6571 | ~n8277);
  assign n6573 = n8280 | ~Pg35 | n6571;
  assign n6574 = Pg35 | ~Ng2338;
  assign n6575_1 = ~Ng2287 & (Ng2331 | ~n8277);
  assign n6576 = ~Pg35 | n6571 | n6575_1 | Ng2361;
  assign n6577 = n6543 & (~Pg35 | (n5873 & ~n6271));
  assign n6578 = Pg35 | ~Ng2153;
  assign n6579 = Pg35 | ~Ng2269;
  assign n6580_1 = Ng2273 | ~Pg35 | n8282;
  assign n6581 = (~Ng2269 | ~n8283) & (n8282 | ~n8695);
  assign n6582 = ~n6271 & n8330;
  assign n6583 = Pg35 & (n6582 | ~n8284);
  assign n6584 = ~Pg35 | n6582 | ~n8284 | ~Ng2153;
  assign n6585_1 = Pg35 | ~Ng2204;
  assign n6586 = ~Ng2153 & (Ng2197 | ~n8284);
  assign n6587 = ~Pg35 | n6582 | n6586 | Ng2227;
  assign n6588 = n6543 & (~Pg35 | (n5921 & ~n6267));
  assign n6589 = Pg35 | ~Ng1996;
  assign n6590_1 = Pg35 | ~Ng2112;
  assign n6591 = Ng2116 | ~Pg35 | n8290;
  assign n6592 = (~Ng2112 | ~n8291) & (n8290 | ~n8700);
  assign n6593 = ~n6267 & n8330;
  assign n6594 = Pg35 & (n6593 | ~n8292);
  assign n6595_1 = ~Pg35 | n6593 | ~n8292 | ~Ng1996;
  assign n6596 = Pg35 | ~Ng2047;
  assign n6597 = ~Ng1996 & (Ng2040 | ~n8292);
  assign n6598 = ~Pg35 | n6593 | n6597 | Ng2070;
  assign n6599 = n6543 & (~Pg35 | (n5887 & ~n6272));
  assign n6600_1 = Pg35 | ~Ng1862;
  assign n6601 = Pg35 | ~Ng1978;
  assign n6602 = Ng1982 | ~Pg35 | n8297;
  assign n6603 = (~Ng1978 | ~n8298) & (n8297 | ~n8705);
  assign n6604 = ~n6272 & n8330;
  assign n6605_1 = Pg35 & (n6604 | ~n8299);
  assign n6606 = ~Pg35 | n6604 | ~n8299 | ~Ng1862;
  assign n6607 = Pg35 | ~Ng1913;
  assign n6608 = ~Ng1862 & (Ng1906 | ~n8299);
  assign n6609 = ~Pg35 | n6604 | n6608 | Ng1936;
  assign n6610_1 = n6543 & (~Pg35 | (n5894 & ~n6266));
  assign n6611 = Pg35 | ~Ng1728;
  assign n6612 = Pg35 | ~Ng1844;
  assign n6613 = Ng1848 | ~Pg35 | n8304;
  assign n6614 = (~Ng1844 | ~n8305) & (n8304 | ~n8710);
  assign n6615_1 = ~n6266 & n8330;
  assign n6616 = Pg35 & (n6615_1 | ~n8306);
  assign n6617 = n8309 | ~Pg35 | n6615_1;
  assign n6618 = Pg35 | ~Ng1779;
  assign n6619 = ~Ng1728 & (Ng1772 | ~n8306);
  assign n6620_1 = ~Pg35 | n6615_1 | n6619 | Ng1802;
  assign n6621 = n6543 & (~Pg35 | (n4162 & ~n6268));
  assign n6622 = Pg35 | ~Ng1592;
  assign n6623 = Pg35 | ~Ng1710;
  assign n6624_1 = Ng1714 | ~Pg35 | n8311;
  assign n6625 = (~Ng1710 | ~n8312) & (n8311 | ~n8715);
  assign n6626 = (n6470 | ~Ng1668) & (n8314 | n9114);
  assign n6627 = n9114 | ~Pg35 | n8315;
  assign n6628 = Pg35 | ~Ng1644;
  assign n6629_1 = ~Ng1592 & (Ng1636 | ~n8313);
  assign n6630 = ~Pg35 | n6629_1 | Ng1668 | n9114;
  assign n6631 = Ng1333 | Ng1322;
  assign n6632 = n6631 & (Ng1345 | ~n8333);
  assign n6633 = n6632 & (Ng1361 | ~n8333);
  assign n6634_1 = n6633 & (Ng1367 | ~n8333);
  assign n6635 = Pg35 & (~n6634_1 | Ng1379 | ~n8333);
  assign n6636 = n8005 | ~Ng1274 | n5090;
  assign n6637 = Pg35 | ~Ng1270;
  assign n6638_1 = Ng990 | Ng979;
  assign n6639 = n6638_1 & (Ng1002 | ~n8339);
  assign n6640 = n6639 & (Ng1018 | ~n8339);
  assign n6641 = n6640 & (Ng1024 | ~n8339);
  assign n6642_1 = Pg35 & (~n6641 | Ng1036 | ~n8339);
  assign n6643 = n8014 | ~Ng930 | n5097;
  assign n6644 = Pg35 | ~Ng925;
  assign n6645 = ~Ng763 | ~n6647 | n7743;
  assign n6646_1 = Pg35 | ~Ng758;
  assign n6647 = ~Ng758 | n6837;
  assign n6648 = Pg35 | ~Ng590;
  assign n6649 = ~Ng590 | n6839;
  assign n6650 = Ng294 | n8243;
  assign n6651_1 = ~n8243 | n7834 | ~Ng294;
  assign n6652 = Ng153 | n8249;
  assign n6653 = ~n8249 | n7402 | ~Ng153;
  assign n6654 = ~Ng6561 | n8346;
  assign n6655 = n6654 & (~n4287_1 | (Ng6561 & Ng6565));
  assign n6656_1 = n7942 & n8344;
  assign n6657 = Pg35 & (Ng6565 | n6656_1);
  assign n6658 = n6656_1 | ~Pg35 | Ng6561;
  assign n6659 = ~Ng6555 | ~Ng6549;
  assign n6660 = Ng6555 | ~Ng6549;
  assign n6661_1 = ~Ng6555 | Ng6549;
  assign n6662 = n6660 & (~Pg35 | n6661_1);
  assign n6663 = ~Ng6215 | n8348;
  assign n6664 = ~Pg35 | ~Ng6227;
  assign n6665_1 = n6663 & (n6664 | (Ng6215 & Ng6219));
  assign n6666 = n8218 & n8347;
  assign n6667 = Pg35 & (Ng6219 | n6666);
  assign n6668 = n6666 | ~Pg35 | Ng6215;
  assign n6669 = ~Ng6203 | ~Ng6209;
  assign n6670_1 = ~Ng6203 | Ng6209;
  assign n6671 = Ng6203 | ~Ng6209;
  assign n6672 = n6670_1 & (~Pg35 | n6671);
  assign n6673 = ~Ng5869 | n8350;
  assign n6674 = n6673 & (~n1064_1 | (Ng5869 & Ng5873));
  assign n6675_1 = n8218 & n8344;
  assign n6676 = Pg35 & (Ng5873 | n6675_1);
  assign n6677 = n6675_1 | ~Pg35 | Ng5869;
  assign n6678 = ~Ng5863 | ~Ng5857;
  assign n6679 = Ng5863 | ~Ng5857;
  assign n6680_1 = ~Ng5863 | Ng5857;
  assign n6681 = n6679 & (~Pg35 | n6680_1);
  assign n6682 = ~Ng5523 | n8351;
  assign n6683 = ~Pg35 | ~Ng5535;
  assign n6684 = n6682 & (n6683 | (Ng5523 & Ng5527));
  assign n6685 = ~n6261 & n8347;
  assign n6686 = Pg35 & (Ng5527 | n6685);
  assign n6687 = n6685 | ~Pg35 | Ng5523;
  assign n6688 = ~Ng5517 | ~Ng5511;
  assign n6689 = Ng5517 | ~Ng5511;
  assign n6690 = ~Ng5517 | Ng5511;
  assign n6691 = n6689 & (~Pg35 | n6690);
  assign n6692 = ~Ng5176 | n8352;
  assign n6693 = ~Pg35 | ~Ng5188;
  assign n6694 = n6692 & (n6693 | (Ng5176 & Ng5180));
  assign n6695 = ~n6261 & n8344;
  assign n6696 = Pg35 & (Ng5180 | n6695);
  assign n6697 = n6695 | ~Pg35 | Ng5176;
  assign n6698 = ~Ng5170 | ~Ng5164;
  assign n6699 = Ng5170 | ~Ng5164;
  assign n6700 = ~Ng5170 | Ng5164;
  assign n6701 = n6699 & (~Pg35 | n6700);
  assign n6702 = n9230 | ~Pg35 | Ng5057;
  assign n6703 = ~n9230 | n6855 | ~Ng5057;
  assign n6704 = (n6860 & ~Ng4549) | (~n5967 & (~n6860 | ~Ng4549));
  assign n6705 = ~n5993 & n6704;
  assign n6706 = n6860 | ~Ng4575;
  assign n6707 = (n6860 & ~Ng4504) | (~n5967 & (~n6860 | ~Ng4504));
  assign n6708 = n6860 | ~Ng4572;
  assign n6709 = n6707 & n6708;
  assign n6710 = ~\[4437]  | n6860;
  assign n6711 = n9231 & (~Pg35 | ~Ng4108 | ~n6712);
  assign n6712 = ~Ng4098 | n8326;
  assign n6713 = ~Ng3869 | n8365;
  assign n6714 = ~Pg35 | ~Ng3881;
  assign n6715 = n6713 & (n6714 | (Ng3869 & Ng3873));
  assign n6716 = n8220 & n8347;
  assign n6717 = Pg35 & (Ng3873 | n6716);
  assign n6718 = n6716 | ~Pg35 | Ng3869;
  assign n6719 = ~Ng3857 | ~Ng3863;
  assign n6720 = ~Ng3857 | Ng3863;
  assign n6721 = Ng3857 | ~Ng3863;
  assign n6722 = n6720 & (~Pg35 | n6721);
  assign n6723 = ~Ng3518 | n8366;
  assign n6724 = ~Pg35 | ~Ng3530;
  assign n6725 = n6723 & (n6724 | (Ng3518 & Ng3522));
  assign n6726 = n8220 & n8344;
  assign n6727 = Pg35 & (Ng3522 | n6726);
  assign n6728 = n6726 | ~Pg35 | Ng3518;
  assign n6729 = ~Ng3512 | ~Ng3506;
  assign n6730 = Ng3512 | ~Ng3506;
  assign n6731 = ~Ng3512 | Ng3506;
  assign n6732 = n6730 & (~Pg35 | n6731);
  assign n6733 = ~Ng3167 | n8367;
  assign n6734 = ~Pg35 | ~Ng3179;
  assign n6735 = n6733 & (n6734 | (Ng3167 & Ng3171));
  assign n6736 = n7942 & n8347;
  assign n6737 = Pg35 & (Ng3171 | n6736);
  assign n6738 = n6736 | ~Pg35 | Ng3167;
  assign n6739 = ~Ng3161 | ~Ng3155;
  assign n6740 = Ng3161 | ~Ng3155;
  assign n6741 = ~Ng3161 | Ng3155;
  assign n6742 = n6740 & (~Pg35 | n6741);
  assign n6743 = Pg35 | ~Ng2748;
  assign n6744 = n8258 ^ Ng2756;
  assign n6745 = ~Pg35 | n5920;
  assign n6746 = n6543 & (~Pg35 | ~n6306) & n6745;
  assign n6747 = n8085 | ~n8329 | ~n5920 | n6306;
  assign n6748 = Pg35 | ~Ng2610;
  assign n6749 = n8369 | n6306 | ~n8368;
  assign n6750 = (Pg35 | ~Ng2625) & (~Ng2610 | n8369);
  assign n6751 = (n6745 & ~Ng2587) | (~Ng2610 & (~n6745 | ~Ng2587));
  assign n6752 = n6751 & n6749;
  assign n6753 = ~n8415 | Ng2619 | n8369;
  assign n6754 = (Pg35 | ~Ng2595) & (n6745 | ~Ng2587);
  assign n6755 = ~Pg35 | n5919;
  assign n6756 = n6543 & (~Pg35 | ~n6303) & n6755;
  assign n6757 = n8087 | ~n8329 | ~n5919 | n6303;
  assign n6758 = Pg35 | ~Ng2476;
  assign n6759 = n8371 | n6303 | ~n8368;
  assign n6760 = (Pg35 | ~Ng2491) & (~Ng2476 | n8371);
  assign n6761 = (n6755 & ~Ng2453) | (~Ng2476 & (~n6755 | ~Ng2453));
  assign n6762 = n6761 & n6759;
  assign n6763 = ~Pg35 | ~Ng2453 | n8416;
  assign n6764 = n6759 & (Ng2485 | Ng2476 | n8371);
  assign n6765 = ~Pg35 | n5925;
  assign n6766 = n6543 & (~Pg35 | ~n6305) & n6765;
  assign n6767 = n8089 | ~n8329 | ~n5925 | n6305;
  assign n6768 = Pg35 | ~Ng2342;
  assign n6769 = n8372 | n6305 | ~n8368;
  assign n6770 = (Pg35 | ~Ng2357) & (~Ng2342 | n8372);
  assign n6771 = (n6765 & ~Ng2319) | (~Ng2342 & (~n6765 | ~Ng2319));
  assign n6772 = n6771 & n6769;
  assign n6773 = ~n8422 | Ng2351 | n8372;
  assign n6774 = (Pg35 | ~Ng2327) & (n6765 | ~Ng2319);
  assign n6775 = ~Pg35 | n5878;
  assign n6776 = n6543 & (~Pg35 | ~n6307) & n6775;
  assign n6777 = n8091 | ~n8329 | ~n5878 | n6307;
  assign n6778 = Pg35 | ~Ng2208;
  assign n6779 = n8374 | n6307 | ~n8368;
  assign n6780 = (Pg35 | ~Ng2223) & (~Ng2208 | n8374);
  assign n6781 = (n6775 & ~Ng2185) | (~Ng2208 & (~n6775 | ~Ng2185));
  assign n6782 = n6781 & n6779;
  assign n6783 = ~n8425 | Ng2217 | n8374;
  assign n6784 = (Pg35 | ~Ng2193) & (n6775 | ~Ng2185);
  assign n6785 = ~Pg35 | n5916;
  assign n6786 = n6543 & (~Pg35 | ~n6309) & n6785;
  assign n6787 = n8093 | ~n8329 | ~n5916 | n6309;
  assign n6788 = Pg35 | ~Ng2051;
  assign n6789 = n8375 | n6309 | ~n8368;
  assign n6790 = (Pg35 | ~Ng2066) & (~Ng2051 | n8375);
  assign n6791 = (n6785 & ~Ng2028) | (~Ng2051 & (~n6785 | ~Ng2028));
  assign n6792 = n6791 & n6789;
  assign n6793 = ~Pg35 | ~Ng2028 | n8426;
  assign n6794 = n6789 & (Ng2051 | Ng2060 | n8375);
  assign n6795 = ~Pg35 | n5899;
  assign n6796 = n6543 & (~Pg35 | ~n6308) & n6795;
  assign n6797 = n8095 | ~n8329 | ~n5899 | n6308;
  assign n6798 = Pg35 | ~Ng1917;
  assign n6799 = n8376 | n6308 | ~n8368;
  assign n6800 = (Pg35 | ~Ng1932) & (~Ng1917 | n8376);
  assign n6801 = (n6795 & ~Ng1894) | (~Ng1917 & (~n6795 | ~Ng1894));
  assign n6802 = n6801 & n6799;
  assign n6803 = ~n8432 | Ng1926 | n8376;
  assign n6804 = (Pg35 | ~Ng1902) & (n6795 | ~Ng1894);
  assign n6805 = ~Pg35 | n5941;
  assign n6806 = n6543 & (~Pg35 | ~n6304) & n6805;
  assign n6807 = n8097 | ~n8329 | ~n5941 | n6304;
  assign n6808 = Pg35 | ~Ng1783;
  assign n6809 = n8377 | n6304 | ~n8368;
  assign n6810 = (Pg35 | ~Ng1798) & (~Ng1783 | n8377);
  assign n6811 = (n6805 & ~Ng1760) | (~Ng1783 & (~n6805 | ~Ng1760));
  assign n6812 = n6811 & n6809;
  assign n6813 = ~n8435 | Ng1792 | n8377;
  assign n6814 = (Pg35 | ~Ng1768) & (n6805 | ~Ng1760);
  assign n6815 = ~Pg35 | n5868;
  assign n6816 = n6543 & (~Pg35 | ~n6310_1) & n6815;
  assign n6817 = n8099 | ~n8329 | ~n5868 | n6310_1;
  assign n6818 = Pg35 | ~Ng1648;
  assign n6819 = n8378 | n6310_1 | ~n8368;
  assign n6820 = (Pg35 | ~Ng1664) & (~Ng1648 | n8378);
  assign n6821 = (n6815 & ~Ng1624) | (~Ng1648 & (~n6815 | ~Ng1624));
  assign n6822 = n6821 & n6819;
  assign n6823 = ~n8438 | Ng1657 | n8378;
  assign n6824 = (Pg35 | ~Ng1632) & (n6815 | ~Ng1624);
  assign n6825 = ~Ng1373 | ~Pg35 | n6634_1;
  assign n6826 = Ng1373 | ~n6634_1 | n7814;
  assign n6827 = ~Ng1270 | ~n6829 | n8005;
  assign n6828 = Pg35 | ~Ng1263;
  assign n6829 = ~Ng1263 | ~n8336;
  assign n6830 = ~Ng1030 | ~Pg35 | n6641;
  assign n6831 = Ng1030 | ~n6641 | n7819;
  assign n6832 = ~Ng925 | ~n6834 | n8014;
  assign n6833 = Pg35 | ~Ng918;
  assign n6834 = ~Ng918 | ~n8342;
  assign n6835 = ~Ng758 | ~n6837 | n7743;
  assign n6836 = Pg35 | ~Ng749;
  assign n6837 = ~Ng749 | n6876;
  assign n6838 = Pg35 | ~Ng582;
  assign n6839 = ~Ng582 | n6879;
  assign n6840 = ~n8242 | Ng291;
  assign n6841 = ~Ng291 | n7834 | n8242;
  assign n6842 = ~n8248 | Ng150;
  assign n6843 = ~Ng150 | n7402 | n8248;
  assign n6844 = (~Ng2950 | ~Ng2955) & (~Ng2927 | ~Ng2922);
  assign n6845 = ~Ng2936 | ~Ng2941;
  assign n6846 = (~Ng2975 | ~Ng2970) & (~Ng2902 | ~Ng2907);
  assign n6847 = (~Ng2965 | ~Ng2960) & (~Ng2917 | ~Ng2912);
  assign n6848 = n6855 | ~n8353 | ~Ng5033 | ~n8355;
  assign n6849 = n6855 | ~Ng5052 | ~n8357 | ~n9229;
  assign n6850 = n8364 | ~Ng5029 | Ng5062;
  assign n6851 = Pg35 & n6850 & (Ng5029 | ~Ng5062);
  assign n6852 = ~Ng5029 | n6855 | Ng5016 | Ng5022;
  assign n6853 = ~Pg35 | n8355;
  assign n6854 = n9234 & (~Pg35 | Ng5046 | n8722);
  assign n6855 = ~Pg35 | n8364;
  assign n6856 = n9235 & (~Pg35 | Ng5041 | n8379);
  assign n6857 = n9236 & (~Pg35 | Ng5037 | n8723);
  assign n6858 = n9237 & (~Pg35 | ~Ng5016 | n8380);
  assign n6859 = ~Ng4372 | ~Pg35 | Ng4581;
  assign n6860 = ~Pg35 | ~Ng4581;
  assign n6861 = n6859 & (n6860 | (Pg72 & Pg73));
  assign n6862 = Pg35 | ~Ng4093;
  assign n6863 = n8326 ^ Ng4098;
  assign n6864 = ~n8257 | ~Ng2748 | n7336;
  assign n6865 = ~Ng2841 | Ng2748 | n8257;
  assign n6866 = ~Ng1367 | ~Pg35 | n6633;
  assign n6867 = n7814 | ~n6633 | Ng1367;
  assign n6868 = n8336 | ~Ng1263 | n8005;
  assign n6869 = Pg35 | ~Ng1259;
  assign n6870 = ~Ng1024 | ~Pg35 | n6640;
  assign n6871 = n7819 | ~n6640 | Ng1024;
  assign n6872 = n8342 | ~Ng918 | n8014;
  assign n6873 = Pg35 | ~Ng914;
  assign n6874 = ~Ng749 | ~n6876 | n7743;
  assign n6875 = Pg35 | ~Ng744;
  assign n6876 = ~Ng744 | n7397;
  assign n6877 = ~Ng582 | ~n6879 | n8183;
  assign n6878 = Pg35 | ~Ng577;
  assign n6879 = ~Ng577 | n7400;
  assign n6880 = Ng164 | ~n8247;
  assign n6881 = n8247 | n7402 | ~Ng164;
  assign n6882 = (~n5880 | ~n8105) & ~n8213;
  assign n6883 = n6885 | n6886;
  assign n6884 = Pg35 & Ng5817;
  assign n6885 = Pg35 & Ng5124;
  assign n6886 = Pg35 & Ng6163;
  assign n6887 = n6883 & (n6884 | (n6885 & n6886));
  assign n6888 = n8104 | n8101 | n8103 | n5880 | n8213 | n8105;
  assign n6889 = Pg35 & Ng3817;
  assign n6890 = Pg35 & Ng3115;
  assign n6891 = (n4205 | n7404) & (~n8381 | ~Ng6657);
  assign n6892 = Pg35 | ~Ng6649;
  assign n6893 = ~Pg35 | ~n6894 | ~Ng6605;
  assign n6894 = ~Ng6561 | n8383;
  assign n6895 = Pg35 | ~Ng6645;
  assign n6896 = Pg35 | ~Ng6641;
  assign n6897 = ~Pg35 | ~n6898 | ~Ng6589;
  assign n6898 = ~Ng6561 | n8384;
  assign n6899 = Pg35 | ~Ng6637;
  assign n6900 = n8222 | n6659;
  assign n6901 = Pg35 | ~Ng6633;
  assign n6902 = ~Pg35 | ~n6903 | ~Ng6649;
  assign n6903 = n6659 | n8383;
  assign n6904 = Pg35 | ~Ng6629;
  assign n6905 = ~Pg35 | ~n6906 | ~Ng6645;
  assign n6906 = n8346 | n6659;
  assign n6907 = Pg35 | ~Ng6625;
  assign n6908 = ~Pg35 | ~n6909 | ~Ng6641;
  assign n6909 = n6659 | n8384;
  assign n6910 = Pg35 | ~Ng6621;
  assign n6911 = ~Pg35 | ~n6912 | ~Ng6637;
  assign n6912 = n8222 | n6661_1;
  assign n6913 = Pg35 | ~Ng6617;
  assign n6914 = n6661_1 | n8383;
  assign n6915 = Pg35 | ~Ng6613;
  assign n6916 = ~Pg35 | ~n6917 | ~Ng6629;
  assign n6917 = n8346 | n6661_1;
  assign n6918 = Pg35 | ~Ng6609;
  assign n6919 = ~Pg35 | ~n6920 | ~Ng6625;
  assign n6920 = n6661_1 | n8384;
  assign n6921 = Pg35 | ~Ng6601;
  assign n6922 = ~Pg35 | ~n6923 | ~Ng6621;
  assign n6923 = n8222 | n6660;
  assign n6924 = Pg35 | ~Ng6593;
  assign n6925 = ~Pg35 | ~n6926 | ~Ng6617;
  assign n6926 = n8383 | n6660;
  assign n6927 = Pg35 | ~Ng6585;
  assign n6928 = ~Pg35 | ~n6929 | ~Ng6613;
  assign n6929 = n8346 | n6660;
  assign n6930 = Pg35 | ~Ng6581;
  assign n6931 = ~Pg35 | ~n6932 | ~Ng6609;
  assign n6932 = n8384 | n6660;
  assign n6933 = Pg35 | ~Ng6605;
  assign n6934 = ~Pg35 | ~n6935 | ~Ng6601;
  assign n6935 = n8222 | n8385;
  assign n6936 = Pg35 | ~Ng6597;
  assign n6937 = ~Pg35 | ~n6938 | ~Ng6593;
  assign n6938 = n8383 | n8385;
  assign n6939 = Pg35 | ~Ng6589;
  assign n6940 = ~Pg35 | ~n6941 | ~Ng6585;
  assign n6941 = n8346 | n8385;
  assign n6942 = Pg35 | ~Ng6573;
  assign n6943 = ~Pg35 | ~n6944 | ~Ng6581;
  assign n6944 = n8384 | n8385;
  assign n6945 = (n4205 | n7435) & (~n8386 | ~Ng6311);
  assign n6946 = Pg35 | ~Ng6303;
  assign n6947 = ~Pg35 | ~n6948 | ~Ng6259;
  assign n6948 = ~Ng6215 | n8387;
  assign n6949 = Pg35 | ~Ng6299;
  assign n6950 = ~Pg35 | ~n6663 | ~Ng6251;
  assign n6951 = Pg35 | ~Ng6295;
  assign n6952 = ~Pg35 | ~n6953 | ~Ng6243;
  assign n6953 = ~Ng6215 | n8388;
  assign n6954 = Pg35 | ~Ng6291;
  assign n6955 = ~Pg35 | ~n6956 | ~Ng6307;
  assign n6956 = n8217 | n6669;
  assign n6957 = Pg35 | ~Ng6287;
  assign n6958 = ~Pg35 | ~n6959 | ~Ng6303;
  assign n6959 = n6669 | n8387;
  assign n6960 = Pg35 | ~Ng6283;
  assign n6961 = ~Pg35 | ~n6962 | ~Ng6299;
  assign n6962 = n8348 | n6669;
  assign n6963 = Pg35 | ~Ng6279;
  assign n6964 = ~Pg35 | ~n6965 | ~Ng6295;
  assign n6965 = n6669 | n8388;
  assign n6966 = Pg35 | ~Ng6275;
  assign n6967 = ~Pg35 | ~n6968 | ~Ng6291;
  assign n6968 = n8217 | n6671;
  assign n6969 = Pg35 | ~Ng6271;
  assign n6970 = n6671 | n8387;
  assign n6971 = Pg35 | ~Ng6267;
  assign n6972 = n8348 | n6671;
  assign n6973 = Pg35 | ~Ng6263;
  assign n6974 = ~Pg35 | ~n6975 | ~Ng6279;
  assign n6975 = n6671 | n8388;
  assign n6976 = Pg35 | ~Ng6255;
  assign n6977 = n8217 | n6670_1;
  assign n6978 = Pg35 | ~Ng6247;
  assign n6979 = ~Pg35 | ~n6980 | ~Ng6271;
  assign n6980 = n8387 | n6670_1;
  assign n6981 = Pg35 | ~Ng6239;
  assign n6982 = ~Pg35 | ~n6983 | ~Ng6267;
  assign n6983 = n8348 | n6670_1;
  assign n6984 = Pg35 | ~Ng6235;
  assign n6985 = ~Pg35 | ~n6986 | ~Ng6263;
  assign n6986 = n8388 | n6670_1;
  assign n6987 = Pg35 | ~Ng6259;
  assign n6988 = ~Pg35 | ~n6989 | ~Ng6255;
  assign n6989 = n8217 | n8389;
  assign n6990 = Pg35 | ~Ng6251;
  assign n6991 = ~Pg35 | ~n6992 | ~Ng6247;
  assign n6992 = n8387 | n8389;
  assign n6993 = Pg35 | ~Ng6243;
  assign n6994 = ~Pg35 | ~n6995 | ~Ng6239;
  assign n6995 = n8348 | n8389;
  assign n6996 = Pg35 | ~Ng6227;
  assign n6997 = ~Pg35 | ~n6998 | ~Ng6235;
  assign n6998 = n8388 | n8389;
  assign n6999 = (n4205 | n7466) & (~n8390 | ~Ng5965);
  assign n7000 = Pg35 | ~Ng5957;
  assign n7001 = ~Pg35 | ~n7002 | ~Ng5913;
  assign n7002 = ~Ng5869 | n8391;
  assign n7003 = Pg35 | ~Ng5953;
  assign n7004 = Pg35 | ~Ng5949;
  assign n7005 = ~Pg35 | ~n7006 | ~Ng5897;
  assign n7006 = ~Ng5869 | n8392;
  assign n7007 = Pg35 | ~Ng5945;
  assign n7008 = n8223 | n6678;
  assign n7009 = Pg35 | ~Ng5941;
  assign n7010 = ~Pg35 | ~n7011 | ~Ng5957;
  assign n7011 = n6678 | n8391;
  assign n7012 = Pg35 | ~Ng5937;
  assign n7013 = ~Pg35 | ~n7014 | ~Ng5953;
  assign n7014 = n8350 | n6678;
  assign n7015 = Pg35 | ~Ng5933;
  assign n7016 = ~Pg35 | ~n7017 | ~Ng5949;
  assign n7017 = n6678 | n8392;
  assign n7018 = Pg35 | ~Ng5929;
  assign n7019 = ~Pg35 | ~n7020 | ~Ng5945;
  assign n7020 = n8223 | n6680_1;
  assign n7021 = Pg35 | ~Ng5925;
  assign n7022 = n6680_1 | n8391;
  assign n7023 = Pg35 | ~Ng5921;
  assign n7024 = ~Pg35 | ~n7025 | ~Ng5937;
  assign n7025 = n8350 | n6680_1;
  assign n7026 = Pg35 | ~Ng5917;
  assign n7027 = ~Pg35 | ~n7028 | ~Ng5933;
  assign n7028 = n6680_1 | n8392;
  assign n7029 = Pg35 | ~Ng5909;
  assign n7030 = ~Pg35 | ~n7031 | ~Ng5929;
  assign n7031 = n8223 | n6679;
  assign n7032 = Pg35 | ~Ng5901;
  assign n7033 = ~Pg35 | ~n7034 | ~Ng5925;
  assign n7034 = n8391 | n6679;
  assign n7035 = Pg35 | ~Ng5893;
  assign n7036 = ~Pg35 | ~n7037 | ~Ng5921;
  assign n7037 = n8350 | n6679;
  assign n7038 = Pg35 | ~Ng5889;
  assign n7039 = ~Pg35 | ~n7040 | ~Ng5917;
  assign n7040 = n8392 | n6679;
  assign n7041 = Pg35 | ~Ng5913;
  assign n7042 = ~Pg35 | ~n7043 | ~Ng5909;
  assign n7043 = n8223 | n8393;
  assign n7044 = Pg35 | ~Ng5905;
  assign n7045 = ~Pg35 | ~n7046 | ~Ng5901;
  assign n7046 = n8391 | n8393;
  assign n7047 = Pg35 | ~Ng5897;
  assign n7048 = ~Pg35 | ~n7049 | ~Ng5893;
  assign n7049 = n8350 | n8393;
  assign n7050 = Pg35 | ~Ng5881;
  assign n7051 = ~Pg35 | ~n7052 | ~Ng5889;
  assign n7052 = n8392 | n8393;
  assign n7053 = (n4205 | n7497) & (~n8394 | ~Ng5619);
  assign n7054 = Pg35 | ~Ng5611;
  assign n7055 = ~Pg35 | ~n7056 | ~Ng5567;
  assign n7056 = ~Ng5523 | n8395;
  assign n7057 = Pg35 | ~Ng5607;
  assign n7058 = Pg35 | ~Ng5603;
  assign n7059 = ~Pg35 | ~n7060 | ~Ng5551;
  assign n7060 = ~Ng5523 | n8396;
  assign n7061 = Pg35 | ~Ng5599;
  assign n7062 = ~Pg35 | ~n7063 | ~Ng5615;
  assign n7063 = n8221 | n6688;
  assign n7064 = Pg35 | ~Ng5595;
  assign n7065 = ~Pg35 | ~n7066 | ~Ng5611;
  assign n7066 = n6688 | n8395;
  assign n7067 = Pg35 | ~Ng5591;
  assign n7068 = ~Pg35 | ~n7069 | ~Ng5607;
  assign n7069 = n8351 | n6688;
  assign n7070 = Pg35 | ~Ng5587;
  assign n7071 = ~Pg35 | ~n7072 | ~Ng5603;
  assign n7072 = n6688 | n8396;
  assign n7073 = Pg35 | ~Ng5583;
  assign n7074 = ~Pg35 | ~n7075 | ~Ng5599;
  assign n7075 = n8221 | n6690;
  assign n7076 = Pg35 | ~Ng5579;
  assign n7077 = n6690 | n8395;
  assign n7078 = Pg35 | ~Ng5575;
  assign n7079 = ~Pg35 | ~n7080 | ~Ng5591;
  assign n7080 = n8351 | n6690;
  assign n7081 = Pg35 | ~Ng5571;
  assign n7082 = ~Pg35 | ~n7083 | ~Ng5587;
  assign n7083 = n6690 | n8396;
  assign n7084 = Pg35 | ~Ng5563;
  assign n7085 = ~Pg35 | ~n7086 | ~Ng5583;
  assign n7086 = n8221 | n6689;
  assign n7087 = Pg35 | ~Ng5555;
  assign n7088 = ~Pg35 | ~n7089 | ~Ng5579;
  assign n7089 = n8395 | n6689;
  assign n7090 = Pg35 | ~Ng5547;
  assign n7091 = ~Pg35 | ~n7092 | ~Ng5575;
  assign n7092 = n8351 | n6689;
  assign n7093 = Pg35 | ~Ng5543;
  assign n7094 = ~Pg35 | ~n7095 | ~Ng5571;
  assign n7095 = n8396 | n6689;
  assign n7096 = Pg35 | ~Ng5567;
  assign n7097 = ~Pg35 | ~n7098 | ~Ng5563;
  assign n7098 = n8221 | n8397;
  assign n7099 = Pg35 | ~Ng5559;
  assign n7100 = ~Pg35 | ~n7101 | ~Ng5555;
  assign n7101 = n8395 | n8397;
  assign n7102 = Pg35 | ~Ng5551;
  assign n7103 = ~Pg35 | ~n7104 | ~Ng5547;
  assign n7104 = n8351 | n8397;
  assign n7105 = Pg35 | ~Ng5535;
  assign n7106 = ~Pg35 | ~n7107 | ~Ng5543;
  assign n7107 = n8396 | n8397;
  assign n7108 = (n7934 | ~Ng5272) & (n4205 | n7527);
  assign n7109 = Pg35 | ~Ng5264;
  assign n7110 = ~Pg35 | ~n7111 | ~Ng5220;
  assign n7111 = ~Ng5176 | n8398;
  assign n7112 = Pg35 | ~Ng5260;
  assign n7113 = ~Pg35 | ~n6692 | ~Ng5212;
  assign n7114 = Pg35 | ~Ng5256;
  assign n7115 = ~Pg35 | ~n7116 | ~Ng5204;
  assign n7116 = ~Ng5176 | n8399;
  assign n7117 = Pg35 | ~Ng5252;
  assign n7118 = ~Pg35 | ~n7119 | ~Ng5268;
  assign n7119 = n8225 | n6698;
  assign n7120 = Pg35 | ~Ng5248;
  assign n7121 = ~Pg35 | ~n7122 | ~Ng5264;
  assign n7122 = n6698 | n8398;
  assign n7123 = Pg35 | ~Ng5244;
  assign n7124 = n8352 | n6698;
  assign n7125 = Pg35 | ~Ng5240;
  assign n7126 = ~Pg35 | ~n7127 | ~Ng5256;
  assign n7127 = n6698 | n8399;
  assign n7128 = Pg35 | ~Ng5236;
  assign n7129 = n8225 | n6700;
  assign n7130 = Pg35 | ~Ng5232;
  assign n7131 = n6700 | n8398;
  assign n7132 = Pg35 | ~Ng5228;
  assign n7133 = ~Pg35 | ~n7134 | ~Ng5244;
  assign n7134 = n8352 | n6700;
  assign n7135 = Pg35 | ~Ng5224;
  assign n7136 = ~Pg35 | ~n7137 | ~Ng5240;
  assign n7137 = n6700 | n8399;
  assign n7138 = Pg35 | ~Ng5216;
  assign n7139 = ~Pg35 | ~n7140 | ~Ng5236;
  assign n7140 = n8225 | n6699;
  assign n7141 = Pg35 | ~Ng5208;
  assign n7142 = ~Pg35 | ~n7143 | ~Ng5232;
  assign n7143 = n8398 | n6699;
  assign n7144 = Pg35 | ~Ng5200;
  assign n7145 = ~Pg35 | ~n7146 | ~Ng5228;
  assign n7146 = n8352 | n6699;
  assign n7147 = Pg35 | ~Ng5196;
  assign n7148 = ~Pg35 | ~n7149 | ~Ng5224;
  assign n7149 = n8399 | n6699;
  assign n7150 = Pg35 | ~Ng5220;
  assign n7151 = ~Pg35 | ~n7152 | ~Ng5216;
  assign n7152 = n8225 | n8400;
  assign n7153 = Pg35 | ~Ng5212;
  assign n7154 = ~Pg35 | ~n7155 | ~Ng5208;
  assign n7155 = n8398 | n8400;
  assign n7156 = Pg35 | ~Ng5204;
  assign n7157 = ~Pg35 | ~n7158 | ~Ng5200;
  assign n7158 = n8352 | n8400;
  assign n7159 = Pg35 | ~Ng5188;
  assign n7160 = ~Pg35 | ~n7161 | ~Ng5196;
  assign n7161 = n8399 | n8400;
  assign n7162 = (~Ng4507 & n9239) | (~Pg113 & (~Ng4507 | ~n9239));
  assign n7163 = n7162 & Pg35;
  assign n7164 = n9241 | ~Pg115 | Ng4157;
  assign n7165 = ~n9241 | Pg115 | Ng4157;
  assign n7166 = n9240 | ~Pg126 | Ng4146;
  assign n7167 = ~n9240 | Pg126 | Ng4146;
  assign n7168 = n7167 & n7164 & n7165 & n7166;
  assign n7169 = ~n8325 | n7566 | ~Ng4093;
  assign n7170 = ~Ng2841 | Ng4093 | n8325;
  assign n7171 = (n4205 | n7568) & (~n8401 | ~Ng3965);
  assign n7172 = Pg35 | ~Ng3957;
  assign n7173 = ~Pg35 | ~n7174 | ~Ng3913;
  assign n7174 = ~Ng3869 | n8402;
  assign n7175 = Pg35 | ~Ng3953;
  assign n7176 = ~Pg35 | ~n6713 | ~Ng3905;
  assign n7177 = Pg35 | ~Ng3949;
  assign n7178 = ~Pg35 | ~n7179 | ~Ng3897;
  assign n7179 = ~Ng3869 | n8403;
  assign n7180 = Pg35 | ~Ng3945;
  assign n7181 = ~Pg35 | ~n7182 | ~Ng3961;
  assign n7182 = n8219 | n6719;
  assign n7183 = Pg35 | ~Ng3941;
  assign n7184 = ~Pg35 | ~n7185 | ~Ng3957;
  assign n7185 = n6719 | n8402;
  assign n7186 = Pg35 | ~Ng3937;
  assign n7187 = n8365 | n6719;
  assign n7188 = Pg35 | ~Ng3933;
  assign n7189 = ~Pg35 | ~n7190 | ~Ng3949;
  assign n7190 = n6719 | n8403;
  assign n7191 = Pg35 | ~Ng3929;
  assign n7192 = n8219 | n6721;
  assign n7193 = Pg35 | ~Ng3925;
  assign n7194 = n6721 | n8402;
  assign n7195 = Pg35 | ~Ng3921;
  assign n7196 = ~Pg35 | ~n7197 | ~Ng3937;
  assign n7197 = n8365 | n6721;
  assign n7198 = Pg35 | ~Ng3917;
  assign n7199 = ~Pg35 | ~n7200 | ~Ng3933;
  assign n7200 = n6721 | n8403;
  assign n7201 = Pg35 | ~Ng3909;
  assign n7202 = ~Pg35 | ~n7203 | ~Ng3929;
  assign n7203 = n8219 | n6720;
  assign n7204 = Pg35 | ~Ng3901;
  assign n7205 = ~Pg35 | ~n7206 | ~Ng3925;
  assign n7206 = n8402 | n6720;
  assign n7207 = Pg35 | ~Ng3893;
  assign n7208 = ~Pg35 | ~n7209 | ~Ng3921;
  assign n7209 = n8365 | n6720;
  assign n7210 = Pg35 | ~Ng3889;
  assign n7211 = ~Pg35 | ~n7212 | ~Ng3917;
  assign n7212 = n8403 | n6720;
  assign n7213 = Pg35 | ~Ng3913;
  assign n7214 = ~Pg35 | ~n7215 | ~Ng3909;
  assign n7215 = n8219 | n8404;
  assign n7216 = Pg35 | ~Ng3905;
  assign n7217 = ~Pg35 | ~n7218 | ~Ng3901;
  assign n7218 = n8402 | n8404;
  assign n7219 = Pg35 | ~Ng3897;
  assign n7220 = ~Pg35 | ~n7221 | ~Ng3893;
  assign n7221 = n8365 | n8404;
  assign n7222 = Pg35 | ~Ng3881;
  assign n7223 = ~Pg35 | ~n7224 | ~Ng3889;
  assign n7224 = n8403 | n8404;
  assign n7225 = (n4205 | n7599) & (~n8405 | ~Ng3614);
  assign n7226 = Pg35 | ~Ng3606;
  assign n7227 = ~Pg35 | ~n7228 | ~Ng3562;
  assign n7228 = ~Ng3518 | n8406;
  assign n7229 = Pg35 | ~Ng3602;
  assign n7230 = ~Pg35 | ~n6723 | ~Ng3554;
  assign n7231 = Pg35 | ~Ng3598;
  assign n7232 = ~Pg35 | ~n7233 | ~Ng3546;
  assign n7233 = ~Ng3518 | n8407;
  assign n7234 = Pg35 | ~Ng3594;
  assign n7235 = ~Pg35 | ~n7236 | ~Ng3610;
  assign n7236 = n8224 | n6729;
  assign n7237 = Pg35 | ~Ng3590;
  assign n7238 = ~Pg35 | ~n7239 | ~Ng3606;
  assign n7239 = n6729 | n8406;
  assign n7240 = Pg35 | ~Ng3586;
  assign n7241 = n8366 | n6729;
  assign n7242 = Pg35 | ~Ng3582;
  assign n7243 = ~Pg35 | ~n7244 | ~Ng3598;
  assign n7244 = n6729 | n8407;
  assign n7245 = Pg35 | ~Ng3578;
  assign n7246 = ~Pg35 | ~n7247 | ~Ng3594;
  assign n7247 = n8224 | n6731;
  assign n7248 = Pg35 | ~Ng3574;
  assign n7249 = n6731 | n8406;
  assign n7250 = Pg35 | ~Ng3570;
  assign n7251 = ~Pg35 | ~n7252 | ~Ng3586;
  assign n7252 = n8366 | n6731;
  assign n7253 = Pg35 | ~Ng3566;
  assign n7254 = ~Pg35 | ~n7255 | ~Ng3582;
  assign n7255 = n6731 | n8407;
  assign n7256 = Pg35 | ~Ng3558;
  assign n7257 = n8224 | n6730;
  assign n7258 = Pg35 | ~Ng3550;
  assign n7259 = ~Pg35 | ~n7260 | ~Ng3574;
  assign n7260 = n8406 | n6730;
  assign n7261 = Pg35 | ~Ng3542;
  assign n7262 = ~Pg35 | ~n7263 | ~Ng3570;
  assign n7263 = n8366 | n6730;
  assign n7264 = Pg35 | ~Ng3538;
  assign n7265 = ~Pg35 | ~n7266 | ~Ng3566;
  assign n7266 = n8407 | n6730;
  assign n7267 = Pg35 | ~Ng3562;
  assign n7268 = ~Pg35 | ~n7269 | ~Ng3558;
  assign n7269 = n8224 | n8408;
  assign n7270 = Pg35 | ~Ng3554;
  assign n7271 = ~Pg35 | ~n7272 | ~Ng3550;
  assign n7272 = n8406 | n8408;
  assign n7273 = Pg35 | ~Ng3546;
  assign n7274 = ~Pg35 | ~n7275 | ~Ng3542;
  assign n7275 = n8366 | n8408;
  assign n7276 = Pg35 | ~Ng3530;
  assign n7277 = ~Pg35 | ~n7278 | ~Ng3538;
  assign n7278 = n8407 | n8408;
  assign n7279 = (n4205 | n7628) & (~n8409 | ~Ng3263);
  assign n7280 = Pg35 | ~Ng3255;
  assign n7281 = ~Pg35 | ~n7282 | ~Ng3211;
  assign n7282 = ~Ng3167 | n8410;
  assign n7283 = Pg35 | ~Ng3251;
  assign n7284 = ~Pg35 | ~n6733 | ~Ng3203;
  assign n7285 = Pg35 | ~Ng3247;
  assign n7286 = ~Pg35 | ~n7287 | ~Ng3195;
  assign n7287 = ~Ng3167 | n8411;
  assign n7288 = Pg35 | ~Ng3243;
  assign n7289 = ~Pg35 | ~n7290 | ~Ng3259;
  assign n7290 = n8216 | n6739;
  assign n7291 = Pg35 | ~Ng3239;
  assign n7292 = ~Pg35 | ~n7293 | ~Ng3255;
  assign n7293 = n6739 | n8410;
  assign n7294 = Pg35 | ~Ng3235;
  assign n7295 = ~Pg35 | ~n7296 | ~Ng3251;
  assign n7296 = n8367 | n6739;
  assign n7297 = Pg35 | ~Ng3231;
  assign n7298 = ~Pg35 | ~n7299 | ~Ng3247;
  assign n7299 = n6739 | n8411;
  assign n7300 = Pg35 | ~Ng3227;
  assign n7301 = ~Pg35 | ~n7302 | ~Ng3243;
  assign n7302 = n8216 | n6741;
  assign n7303 = Pg35 | ~Ng3223;
  assign n7304 = n6741 | n8410;
  assign n7305 = Pg35 | ~Ng3219;
  assign n7306 = n8367 | n6741;
  assign n7307 = Pg35 | ~Ng3215;
  assign n7308 = ~Pg35 | ~n7309 | ~Ng3231;
  assign n7309 = n6741 | n8411;
  assign n7310 = Pg35 | ~Ng3207;
  assign n7311 = n8216 | n6740;
  assign n7312 = Pg35 | ~Ng3199;
  assign n7313 = ~Pg35 | ~n7314 | ~Ng3223;
  assign n7314 = n8410 | n6740;
  assign n7315 = Pg35 | ~Ng3191;
  assign n7316 = ~Pg35 | ~n7317 | ~Ng3219;
  assign n7317 = n8367 | n6740;
  assign n7318 = Pg35 | ~Ng3187;
  assign n7319 = ~Pg35 | ~n7320 | ~Ng3215;
  assign n7320 = n8411 | n6740;
  assign n7321 = Pg35 | ~Ng3211;
  assign n7322 = ~Pg35 | ~n7323 | ~Ng3207;
  assign n7323 = n8216 | n8412;
  assign n7324 = Pg35 | ~Ng3203;
  assign n7325 = ~Pg35 | ~n7326 | ~Ng3199;
  assign n7326 = n8410 | n8412;
  assign n7327 = Pg35 | ~Ng3195;
  assign n7328 = ~Pg35 | ~n7329 | ~Ng3191;
  assign n7329 = n8367 | n8412;
  assign n7330 = Pg35 | ~Ng3179;
  assign n7331 = ~Pg35 | ~n7332 | ~Ng3187;
  assign n7332 = n8411 | n8412;
  assign n7333 = n9246 | ~Pg35 | n9245;
  assign n7334 = n9250 | ~Pg35 | n9249;
  assign n7335 = n8106 ^ Ng2741;
  assign n7336 = ~Pg35 | ~Ng2841;
  assign n7337 = Ng2681 | Ng2675 | ~n8414;
  assign n7338 = ~Pg35 | n8413;
  assign n7339 = (~n8414 & ~Ng2661) | (n7338 & (~n8414 | Ng2661));
  assign n7340 = n8415 | n8107 | n8369;
  assign n7341 = n8369 | n8264 | n8205;
  assign n7342 = Ng2547 | Ng2541 | ~n8418;
  assign n7343 = ~Pg35 | n8417;
  assign n7344 = (~Ng2527 & ~n8418) | (n7343 & (Ng2527 | ~n8418));
  assign n7345 = n8419 | n8108 | n8371;
  assign n7346 = n8371 | n8271 | n8203;
  assign n7347 = Ng2413 | Ng2407 | ~n8421;
  assign n7348 = ~Pg35 | n8420;
  assign n7349 = (~n8421 & ~Ng2393) | (n7348 & (~n8421 | Ng2393));
  assign n7350 = n8422 | n8109 | n8372;
  assign n7351 = n8372 | n8278 | n8204;
  assign n7352 = Ng2279 | Ng2273 | ~n8424;
  assign n7353 = ~Pg35 | n8423;
  assign n7354 = (~n8424 & ~Ng2259) | (n7353 & (~n8424 | Ng2259));
  assign n7355 = n8425 | n8110 | n8374;
  assign n7356 = n8374 | n8286 | n8197;
  assign n7357 = Ng2122 | Ng2116 | ~n8428;
  assign n7358 = ~Pg35 | n8427;
  assign n7359 = (~Ng2102 & ~n8428) | (n7358 & (Ng2102 | ~n8428));
  assign n7360 = n8429 | n8111 | n8375;
  assign n7361 = n8375 | n8294 | n8201;
  assign n7362 = Ng1988 | Ng1982 | ~n8431;
  assign n7363 = ~Pg35 | n8430;
  assign n7364 = (~Ng1968 & ~n8431) | (n7363 & (Ng1968 | ~n8431));
  assign n7365 = n8432 | n8112 | n8376;
  assign n7366 = n8376 | n8301 | n8202;
  assign n7367 = Ng1854 | Ng1848 | ~n8434;
  assign n7368 = ~Pg35 | n8433;
  assign n7369 = (~n8434 & ~Ng1834) | (n7368 & (~n8434 | Ng1834));
  assign n7370 = n8435 | n8113 | n8377;
  assign n7371 = n8377 | n8307 | n8199;
  assign n7372 = Ng1720 | Ng1714 | ~n8437;
  assign n7373 = ~Pg35 | n8436;
  assign n7374 = (~n8437 & ~Ng1700) | (n7373 & (~n8437 | Ng1700));
  assign n7375 = n8438 | n8114 | n8378;
  assign n7376 = ~n8207 & ~n8378 & (~Ng1636 | Ng1592);
  assign n7377 = ~n5559 & (~Ng1526 | ~n7379);
  assign n7378 = (n7377 & (Pg35 | ~Ng1514)) | (~Pg35 & ~Ng1514);
  assign n7379 = ~Pg7946 | ~Ng1514;
  assign n7380 = ~Ng1361 | ~Pg35 | n6632;
  assign n7381 = n7814 | ~n6632 | Ng1361;
  assign n7382 = ~Ng1259 | ~n7384 | n8005;
  assign n7383 = Pg35 | ~Ng1256;
  assign n7384 = ~Ng1256 | ~n8335;
  assign n7385 = n8083 & Ng1024 & Ng1002 & Ng1036;
  assign n7386 = n7385 | Ng1008 | Ng969;
  assign n7387 = ~n4474 & (~Ng1183 | ~n7389);
  assign n7388 = (Pg35 & n7387) | (~Ng1171 & (~Pg35 | n7387));
  assign n7389 = ~Pg7916 | ~Ng1171;
  assign n7390 = ~Ng1018 | ~Pg35 | n6639;
  assign n7391 = n7819 | ~n6639 | Ng1018;
  assign n7392 = ~Ng914 | ~n7394 | n8014;
  assign n7393 = Pg35 | ~Ng911;
  assign n7394 = ~Ng911 | ~n8341;
  assign n7395 = ~Ng744 | ~n7397 | n7743;
  assign n7396 = Pg35 | ~Ng739;
  assign n7397 = ~n6091_1 | ~Ng739 | n8180;
  assign n7398 = ~Ng577 | ~n7400 | n8183;
  assign n7399 = Pg35 | ~Ng586;
  assign n7400 = ~Ng586 | n7754;
  assign n7401 = ~n4520 ^ Ng146;
  assign n7402 = ~Pg35 | n8246;
  assign n7403 = ~Ng6541 | ~n8381 | ~n8382;
  assign n7404 = ~Ng6561 | n8222;
  assign n7405 = (n7407 & (n8441 | Ng6527)) | (n8441 & ~Ng6527);
  assign n7406 = Ng6519 | Ng6513 | n8441;
  assign n7407 = ~Pg35 | ~n8440;
  assign n7408 = ~Ng6505 | Ng6500 | n8441;
  assign n7409 = (~Pg13099 | ~Ng6593) & (~Ng6605 | ~Ng6723);
  assign n7410 = (~Pg17764 | ~Ng6649) & (~Pg17722 | ~Ng6597);
  assign n7411 = (~Pg17871 | ~Ng6617) & (~Pg12470 | ~Ng6601);
  assign n7412 = ~Ng6633 | ~Pg14749 | n7423;
  assign n7413 = (n7410 | n6496) & (n7409 | n7426);
  assign n7414 = ~Ng6741 | ~Ng6682;
  assign n7415 = n7412 & n7413 & (n7411 | n7414);
  assign n7416 = (~Pg13099 | ~Ng6581) & (~Ng6589 | ~Ng6723);
  assign n7417 = (~Pg17871 | ~Ng6609) & (~Pg12470 | ~Ng6585);
  assign n7418 = ~Ng6641 | ~Pg17764 | n7414;
  assign n7419 = ~Ng6625 | ~Pg14749 | n7426;
  assign n7420 = (n7417 | n6496) & (n7416 | n7423);
  assign n7421 = n7418 & n7419 & n7420;
  assign n7422 = n9123 & (~Pg17778 | n6496 | ~Ng6637);
  assign n7423 = Ng6682 | Ng6741;
  assign n7424 = n7422 & (~Pg14828 | n7423 | ~Ng6621);
  assign n7425 = n9122 & (~Pg17778 | n7414 | ~Ng6629);
  assign n7426 = Ng6741 | ~Ng6682;
  assign n7427 = n7425 & (~Pg14828 | n7426 | ~Ng6613);
  assign n7428 = (n7421 & Ng6727) | (n7415 & (n7421 | ~Ng6727));
  assign n7429 = (n7427 & n9279) | (n7424 & (n7427 | ~n9279));
  assign n7430 = ~Ng6727 | ~Pg17722 | n7414;
  assign n7431 = n7428 & n7429 & (n7430 | ~Ng6657);
  assign n7432 = Pg35 | ~Ng6505;
  assign n7433 = ~Pg35 | ~n5884_1 | n7431;
  assign n7434 = ~Ng6195 | ~n8382 | ~n8386;
  assign n7435 = ~Ng6215 | n8217;
  assign n7436 = (n7438 & (n8443 | Ng6181)) | (n8443 & ~Ng6181);
  assign n7437 = Ng6173 | Ng6167 | n8443;
  assign n7438 = ~Pg35 | ~n8442;
  assign n7439 = ~Ng6159 | Ng6154 | n8443;
  assign n7440 = (~Pg17743 | ~Ng6303) & (~Pg17685 | ~Ng6251);
  assign n7441 = (~Pg13085 | ~Ng6247) & (~Ng6259 | ~Ng6377);
  assign n7442 = (~Pg17845 | ~Ng6271) & (~Pg12422 | ~Ng6255);
  assign n7443 = ~Ng6287 | ~Pg14705 | n7457;
  assign n7444 = (n7441 | n7454) & (n7440 | n6502_1);
  assign n7445 = ~Ng6395 | ~Ng6336;
  assign n7446 = n7443 & n7444 & (n7442 | n7445);
  assign n7447 = (~Pg13085 | ~Ng6235) & (~Ng6243 | ~Ng6377);
  assign n7448 = (~Pg17845 | ~Ng6263) & (~Pg12422 | ~Ng6239);
  assign n7449 = ~Ng6295 | ~Pg17743 | n7445;
  assign n7450 = ~Ng6279 | ~Pg14705 | n7454;
  assign n7451 = (n7448 | n6502_1) & (n7447 | n7457);
  assign n7452 = n7449 & n7450 & n7451;
  assign n7453 = n9125 & (~Pg17760 | n6502_1 | ~Ng6291);
  assign n7454 = Ng6395 | ~Ng6336;
  assign n7455 = n7453 & (~Pg17649 | n7454 | ~Ng6307);
  assign n7456 = n9124 & (~Pg14779 | n7454 | ~Ng6267);
  assign n7457 = Ng6336 | Ng6395;
  assign n7458 = n7456 & (~Pg17649 | n7457 | ~Ng6299);
  assign n7459 = (n7452 & Ng6381) | (n7446 & (n7452 | ~Ng6381));
  assign n7460 = (n7458 & n9283) | (n7455 & (n7458 | ~n9283));
  assign n7461 = ~Ng6381 | ~Pg17685 | n7445;
  assign n7462 = n7459 & n7460 & (n7461 | ~Ng6311);
  assign n7463 = Pg35 | ~Ng6159;
  assign n7464 = ~Pg35 | ~n5952 | n7462;
  assign n7465 = ~Ng5849 | ~n8382 | ~n8390;
  assign n7466 = ~Ng5869 | n8223;
  assign n7467 = (n7469 & (n8445 | Ng5835)) | (n8445 & ~Ng5835);
  assign n7468 = Ng5827 | Ng5821 | n8445;
  assign n7469 = ~Pg35 | ~n8444;
  assign n7470 = ~Ng5813 | Ng5808 | n8445;
  assign n7471 = (~Pg13068 | ~Ng5901) & (~Ng5913 | ~Ng6031);
  assign n7472 = (~Pg17715 | ~Ng5957) & (~Pg17646 | ~Ng5905);
  assign n7473 = (~Pg17819 | ~Ng5925) & (~Pg12350 | ~Ng5909);
  assign n7474 = ~Ng5941 | ~Pg14673 | n7485;
  assign n7475 = (n7472 | n6508) & (n7471 | n7488);
  assign n7476 = ~Ng6049 | ~Ng5990;
  assign n7477 = n7474 & n7475 & (n7473 | n7476);
  assign n7478 = (~Pg13068 | ~Ng5889) & (~Ng5897 | ~Ng6031);
  assign n7479 = (~Pg17819 | ~Ng5917) & (~Pg12350 | ~Ng5893);
  assign n7480 = ~Ng5933 | ~Pg14673 | n7488;
  assign n7481 = ~Ng5949 | ~Pg17715 | n7476;
  assign n7482 = (n7479 | n6508) & (n7478 | n7485);
  assign n7483 = n7480 & n7481 & n7482;
  assign n7484 = n9127 & (~Pg17739 | n6508 | ~Ng5945);
  assign n7485 = Ng5990 | Ng6049;
  assign n7486 = n7484 & (~Pg14738 | n7485 | ~Ng5929);
  assign n7487 = n9126 & (~Pg17739 | n7476 | ~Ng5937);
  assign n7488 = Ng6049 | ~Ng5990;
  assign n7489 = n7487 & (~Pg14738 | n7488 | ~Ng5921);
  assign n7490 = (n7483 & Ng6035) | (n7477 & (n7483 | ~Ng6035));
  assign n7491 = (n7489 & n9287) | (n7486 & (n7489 | ~n9287));
  assign n7492 = ~Ng6035 | ~Pg17646 | n7476;
  assign n7493 = n7490 & n7491 & (n7492 | ~Ng5965);
  assign n7494 = Pg35 | ~Ng5813;
  assign n7495 = ~Pg35 | ~n5940 | n7493;
  assign n7496 = ~Ng5503 | ~n8382 | ~n8394;
  assign n7497 = ~Ng5523 | n8221;
  assign n7498 = (n7500 & (n8447 | Ng5489)) | (n8447 & ~Ng5489);
  assign n7499 = Ng5481 | Ng5475 | n8447;
  assign n7500 = ~Pg35 | ~n8446;
  assign n7501 = Ng5462 | n8447 | ~Ng5467;
  assign n7502 = (~Pg17678 | ~Ng5611) & (~Pg17604 | ~Ng5559);
  assign n7503 = (~Pg13049 | ~Ng5555) & (~Ng5567 | ~Ng5685);
  assign n7504 = (~Pg17813 | ~Ng5579) & (~Pg12300 | ~Ng5563);
  assign n7505 = ~Ng5595 | ~Pg14635 | n7516;
  assign n7506 = (n7503 | n7519) & (n7502 | n8321);
  assign n7507 = ~Ng5703 | ~Ng5644;
  assign n7508 = n7505 & n7506 & (n7504 | n7507);
  assign n7509 = (~Pg17813 | ~Ng5571) & (~Pg12300 | ~Ng5547);
  assign n7510 = (~Pg13049 | ~Ng5543) & (~Ng5551 | ~Ng5685);
  assign n7511 = ~Ng5603 | ~Pg17678 | n7507;
  assign n7512 = ~Ng5587 | ~Pg14635 | n7519;
  assign n7513 = (n7510 | n7516) & (n7509 | n8321);
  assign n7514 = n7511 & n7512 & n7513;
  assign n7515 = n9129 & (~Pg17711 | n8321 | ~Ng5599);
  assign n7516 = Ng5644 | Ng5703;
  assign n7517 = n7515 & (~Pg14694 | n7516 | ~Ng5583);
  assign n7518 = n9128 & (~Pg17711 | n7507 | ~Ng5591);
  assign n7519 = Ng5703 | ~Ng5644;
  assign n7520 = n7518 & (~Pg14694 | n7519 | ~Ng5575);
  assign n7521 = (n7514 & Ng5689) | (n7508 & (n7514 | ~Ng5689));
  assign n7522 = (n7520 & n9291) | (n7517 & (n7520 | ~n9291));
  assign n7523 = ~Ng5689 | ~Pg17604 | n7507;
  assign n7524 = n7521 & n7522 & (n7523 | ~Ng5619);
  assign n7525 = n8322 | Ng5462 | n7524;
  assign n7526 = ~n8382 | ~Ng5156 | n7934;
  assign n7527 = ~Ng5176 | n8225;
  assign n7528 = (n7530 & (n8450 | Ng5142)) | (n8450 & ~Ng5142);
  assign n7529 = Ng5134 | Ng5128 | n8450;
  assign n7530 = ~Pg35 | ~n8449;
  assign n7531 = ~Ng5120 | Ng5115 | n8450;
  assign n7532 = (~Pg17787 | ~Ng5232) & (~Pg12238 | ~Ng5216);
  assign n7533 = (~Pg13039 | ~Ng5208) & (~Ng5220 | ~Ng5339);
  assign n7534 = (~Pg17639 | ~Ng5264) & (~Pg17577 | ~Ng5212);
  assign n7535 = ~Ng5248 | ~Pg14597 | n7545;
  assign n7536 = (n7533 | n7548) & (n7532 | n8192);
  assign n7537 = n7535 & n7536 & (n7534 | n6516);
  assign n7538 = (~Pg17787 | ~Ng5224) & (~Pg12238 | ~Ng5200);
  assign n7539 = (~Pg13039 | ~Ng5196) & (~Ng5204 | ~Ng5339);
  assign n7540 = ~Ng5240 | ~Pg14597 | n7548;
  assign n7541 = ~Ng5256 | ~Pg17639 | n8192;
  assign n7542 = (n7539 | n7545) & (n7538 | n6516);
  assign n7543 = n7540 & n7541 & n7542;
  assign n7544 = n9131 & (~Pg17519 | n7548 | ~Ng5268);
  assign n7545 = Ng5297 | Ng5357;
  assign n7546 = n7544 & (~Pg14662 | n7545 | ~Ng5236);
  assign n7547 = n9130 & (~Pg17674 | n8192 | ~Ng5244);
  assign n7548 = Ng5357 | ~Ng5297;
  assign n7549 = n7547 & (~Pg14662 | n7548 | ~Ng5228);
  assign n7550 = (n7537 & (~\[4415]  | n7543)) | (\[4415]  & n7543);
  assign n7551 = (n7549 & n9295) | (n7546 & (n7549 | ~n9295));
  assign n7552 = n7550 & n7551 & (~Ng5272 | ~n8448);
  assign n7553 = Pg35 | ~Ng5120;
  assign n7554 = ~Pg35 | ~n4151_1 | n7552;
  assign n7555 = n5907 & n5888 & (Ng4927 | n5926);
  assign n7556 = Ng4975 | ~Ng4912 | Ng4899;
  assign n7557 = (n5888 | ~Ng4922) & (n5926 | ~Ng4917);
  assign n7558 = n7556 & n7557 & (n5907 | ~Ng4907);
  assign n7559 = ~Ng4966 & (~n5935 | ~Ng4983) & ~n9297;
  assign n7560 = n5939 & n5874_1 & (Ng4737 | n5951);
  assign n7561 = Ng4785 | ~Ng4722 | Ng4709;
  assign n7562 = (n5874_1 | ~Ng4717) & (n5951 | ~Ng4727);
  assign n7563 = n7561 & n7562 & (n5939 | ~Ng4732);
  assign n7564 = ~Ng4776 & (~n5949 | ~Ng4793) & ~n9299;
  assign n7565 = n8121 ^ Ng4087;
  assign n7566 = ~Pg35 | ~Ng2841;
  assign n7567 = ~Ng3849 | ~n8382 | ~n8401;
  assign n7568 = ~Ng3869 | n8219;
  assign n7569 = (n7571 & (n8452 | Ng3835)) | (n8452 & ~Ng3835);
  assign n7570 = Ng3827 | Ng3821 | n8452;
  assign n7571 = ~Pg35 | ~n8451;
  assign n7572 = ~Ng3813 | Ng3808 | n8452;
  assign n7573 = (~Pg14518 | ~Ng3901) & (~Ng3913 | ~Ng4031);
  assign n7574 = (~Pg16748 | ~Ng3957) & (~Pg16693 | ~Ng3905);
  assign n7575 = (~Pg16955 | ~Ng3925) & (~Pg11418 | ~Ng3909);
  assign n7576 = ~Ng3941 | ~Pg13906 | n7587;
  assign n7577 = (n7574 | n6525) & (n7573 | n7590);
  assign n7578 = ~Ng4054 | ~Ng3990;
  assign n7579 = n7576 & n7577 & (n7575 | n7578);
  assign n7580 = (~Pg16955 | ~Ng3917) & (~Pg11418 | ~Ng3893);
  assign n7581 = (~Pg14518 | ~Ng3889) & (~Ng3897 | ~Ng4031);
  assign n7582 = ~Ng3949 | ~Pg16748 | n7578;
  assign n7583 = ~Ng3933 | ~Pg13906 | n7590;
  assign n7584 = (n7581 | n7587) & (n7580 | n6525);
  assign n7585 = n7582 & n7583 & n7584;
  assign n7586 = n9137 & (~Pg16659 | n7590 | ~Ng3961);
  assign n7587 = Ng3990 | Ng4054;
  assign n7588 = n7586 & (~Pg13966 | n7587 | ~Ng3929);
  assign n7589 = n9136 & (~Pg16775 | n7578 | ~Ng3937);
  assign n7590 = Ng4054 | ~Ng3990;
  assign n7591 = n7589 & (~Pg13966 | n7590 | ~Ng3921);
  assign n7592 = (n7585 & Ng4040) | (n7579 & (n7585 | ~Ng4040));
  assign n7593 = (n7591 & n9303) | (n7588 & (n7591 | ~n9303));
  assign n7594 = ~Ng4040 | ~Pg16693 | n7578;
  assign n7595 = n7592 & n7593 & (n7594 | ~Ng3965);
  assign n7596 = Pg35 | ~Ng3813;
  assign n7597 = ~Pg35 | ~n5927 | n7595;
  assign n7598 = ~Ng3498 | ~n8382 | ~n8405;
  assign n7599 = ~Ng3518 | n8224;
  assign n7600 = (n7602 & (n8454 | Ng3484)) | (n8454 & ~Ng3484);
  assign n7601 = Ng3476 | Ng3470 | n8454;
  assign n7602 = ~Pg35 | ~n8453;
  assign n7603 = ~Ng3462 | Ng3457 | n8454;
  assign n7604 = (~Pg16924 | ~Ng3574) & (~Pg11388 | ~Ng3558);
  assign n7605 = (~Pg14451 | ~Ng3550) & (~Ng3562 | ~Ng3680);
  assign n7606 = (~Pg16722 | ~Ng3606) & (~Pg16656 | ~Ng3554);
  assign n7607 = ~Ng3590 | ~Pg13881 | n8455;
  assign n7608 = (n7605 | n8327) & (n7604 | n7619);
  assign n7609 = n7607 & n7608 & (n7606 | n6531_1);
  assign n7610 = (~Pg14451 | ~Ng3538) & (~Ng3546 | ~Ng3680);
  assign n7611 = (~Pg16924 | ~Ng3566) & (~Pg11388 | ~Ng3542);
  assign n7612 = ~Ng3582 | ~Pg13881 | n8327;
  assign n7613 = ~Ng3598 | ~Pg16722 | n7619;
  assign n7614 = (n7611 | n6531_1) & (n7610 | n8455);
  assign n7615 = n7612 & n7613 & n7614;
  assign n7616 = n9139 & (~Pg16627 | n8327 | ~Ng3610);
  assign n7617 = n7616 & (~Pg16744 | n6531_1 | ~Ng3594);
  assign n7618 = n9138 & (~Pg13926 | n8327 | ~Ng3570);
  assign n7619 = ~Ng3703 | ~Ng3639;
  assign n7620 = n7618 & (~Pg16744 | n7619 | ~Ng3586);
  assign n7621 = (n7615 & Ng3689) | (n7609 & (n7615 | ~Ng3689));
  assign n7622 = (n7620 & n9307) | (n7617 & (n7620 | ~n9307));
  assign n7623 = ~Ng3689 | ~Pg16656 | n7619;
  assign n7624 = n7621 & n7622 & (n7623 | ~Ng3614);
  assign n7625 = Pg35 | ~Ng3462;
  assign n7626 = ~Pg35 | ~n5889 | n7624;
  assign n7627 = ~Ng3147 | ~n8382 | ~n8409;
  assign n7628 = ~Ng3167 | n8216;
  assign n7629 = (n7631 & (n8457 | Ng3133)) | (n8457 & ~Ng3133);
  assign n7630 = Ng3125 | Ng3119 | n8457;
  assign n7631 = ~Pg35 | ~n8456;
  assign n7632 = Ng3106 | n8457 | ~Ng3111;
  assign n7633 = (~Pg16686 | ~Ng3255) & (~Pg16624 | ~Ng3203);
  assign n7634 = (~Pg16874 | ~Ng3223) & (~Pg11349 | ~Ng3207);
  assign n7635 = (~Pg14421 | ~Ng3199) & (~Ng3211 | ~Ng3329);
  assign n7636 = ~Ng3239 | ~Pg13865 | n7649;
  assign n7637 = (n7634 | n8189) & (n7633 | n6537);
  assign n7638 = Ng3352 | ~Ng3288;
  assign n7639 = n7636 & n7637 & (n7635 | n7638);
  assign n7640 = (~Pg16874 | ~Ng3215) & (~Pg11349 | ~Ng3191);
  assign n7641 = (~Pg14421 | ~Ng3187) & (~Ng3195 | ~Ng3329);
  assign n7642 = ~Ng3247 | ~Pg16686 | n8189;
  assign n7643 = ~Ng3231 | ~Pg13865 | n7638;
  assign n7644 = (n7641 | n7649) & (n7640 | n6537);
  assign n7645 = n7642 & n7643 & n7644;
  assign n7646 = n9141 & (~Pg16718 | n6537 | ~Ng3243);
  assign n7647 = n7646 & (~Pg16603 | n7638 | ~Ng3259);
  assign n7648 = n9140 & (~Pg13895 | n7638 | ~Ng3219);
  assign n7649 = Ng3288 | Ng3352;
  assign n7650 = n7648 & (~Pg16603 | n7649 | ~Ng3251);
  assign n7651 = (n7645 & Ng3338) | (n7639 & (n7645 | ~Ng3338));
  assign n7652 = (n7650 & n9311) | (n7647 & (n7650 | ~n9311));
  assign n7653 = ~Ng3338 | ~Pg16624 | n8189;
  assign n7654 = n7651 & n7652 & (n7653 | ~Ng3263);
  assign n7655 = n8328 | Ng3106 | n7654;
  assign n7656 = n9313 & (~Pg35 | ~Ng2735 | ~n7657);
  assign n7657 = ~Ng2729 | n8256;
  assign n7658 = n5920 & (~n7659 | ~n8415);
  assign n7659 = ~Ng2638 | ~Ng2652 | ~n8415;
  assign n7660 = Ng2638 & (~Pg35 | (n5920 & n7659));
  assign n7661 = (~Ng2619 | ~Ng2571) & (~Ng2579 | ~Ng2587);
  assign n7662 = Ng2587 | Ng2619 | ~Ng2575;
  assign n7663 = (n8205 | ~Ng2583) & (~Ng2563 | n8415);
  assign n7664 = n7662 & n7663 & (Ng2610 | n7661);
  assign n7665 = n6745 | ~Ng2638;
  assign n7666 = (Pg35 | ~Ng2619) & (n7664 | n8369);
  assign n7667 = n5919 & (~n7668 | ~n8419);
  assign n7668 = ~Ng2504 | ~Ng2518 | ~n8419;
  assign n7669 = Ng2504 & (~Pg35 | (n5919 & n7668));
  assign n7670 = (~Ng2485 | ~Ng2437) & (~Ng2445 | ~Ng2453);
  assign n7671 = Ng2453 | Ng2485 | ~Ng2441;
  assign n7672 = (n8203 | ~Ng2449) & (~Ng2429 | n8419);
  assign n7673 = n7671 & n7672 & (Ng2476 | n7670);
  assign n7674 = n6755 | ~Ng2504;
  assign n7675 = (Pg35 | ~Ng2485) & (n7673 | n8371);
  assign n7676 = n8422 & Ng2384 & Ng2370;
  assign n7677 = n5925 & (n7676 | ~n8422);
  assign n7678 = Ng2370 & (~Pg35 | (n5925 & ~n7676));
  assign n7679 = (~Ng2351 | ~Ng2303) & (~Ng2311 | ~Ng2319);
  assign n7680 = Ng2319 | Ng2351 | ~Ng2307;
  assign n7681 = (n8204 | ~Ng2315) & (~Ng2295 | n8422);
  assign n7682 = n7680 & n7681 & (Ng2342 | n7679);
  assign n7683 = n6765 | ~Ng2370;
  assign n7684 = (Pg35 | ~Ng2351) & (n7682 | n8372);
  assign n7685 = n8425 & Ng2250 & Ng2236;
  assign n7686 = n5878 & (n7685 | ~n8425);
  assign n7687 = Ng2236 & (~Pg35 | (n5878 & ~n7685));
  assign n7688 = (~Ng2217 | ~Ng2169) & (~Ng2177 | ~Ng2185);
  assign n7689 = Ng2185 | Ng2217 | ~Ng2173;
  assign n7690 = (n8197 | ~Ng2181) & (~Ng2161 | n8425);
  assign n7691 = n7689 & n7690 & (Ng2208 | n7688);
  assign n7692 = n6775 | ~Ng2236;
  assign n7693 = (Pg35 | ~Ng2217) & (n7691 | n8374);
  assign n7694 = n8429 & Ng2093 & Ng2079;
  assign n7695 = n5916 & (n7694 | ~n8429);
  assign n7696 = Ng2079 & (~Pg35 | (n5916 & ~n7694));
  assign n7697 = (~Ng2060 | ~Ng2012) & (~Ng2020 | ~Ng2028);
  assign n7698 = Ng2028 | Ng2060 | ~Ng2016;
  assign n7699 = (n8201 | ~Ng2024) & (~Ng2004 | n8429);
  assign n7700 = n7698 & n7699 & (Ng2051 | n7697);
  assign n7701 = n6785 | ~Ng2079;
  assign n7702 = (Pg35 | ~Ng2060) & (n7700 | n8375);
  assign n7703 = n8432 & Ng1959 & Ng1945;
  assign n7704 = n5899 & (n7703 | ~n8432);
  assign n7705 = Ng1945 & (~Pg35 | (n5899 & ~n7703));
  assign n7706 = (~Ng1926 | ~Ng1878) & (~Ng1886 | ~Ng1894);
  assign n7707 = Ng1894 | Ng1926 | ~Ng1882;
  assign n7708 = (n8202 | ~Ng1890) & (~Ng1870 | n8432);
  assign n7709 = n7707 & n7708 & (Ng1917 | n7706);
  assign n7710 = n6795 | ~Ng1945;
  assign n7711 = (Pg35 | ~Ng1926) & (n7709 | n8376);
  assign n7712 = n5941 & (~n7713 | ~n8435);
  assign n7713 = ~Ng1811 | ~Ng1825 | ~n8435;
  assign n7714 = Ng1811 & (~Pg35 | (n5941 & n7713));
  assign n7715 = (~Ng1792 | ~Ng1744) & (~Ng1752 | ~Ng1760);
  assign n7716 = Ng1760 | Ng1792 | ~Ng1748;
  assign n7717 = (n8199 | ~Ng1756) & (~Ng1736 | n8435);
  assign n7718 = n7716 & n7717 & (Ng1783 | n7715);
  assign n7719 = n6805 | ~Ng1811;
  assign n7720 = (Pg35 | ~Ng1792) & (n7718 | n8377);
  assign n7721 = n5868 & (~n7722 | ~n8438);
  assign n7722 = ~Ng1677 | ~Ng1691 | ~n8438;
  assign n7723 = Ng1677 & (~Pg35 | (n5868 & n7722));
  assign n7724 = (~Ng1657 | ~Ng1608) & (~Ng1616 | ~Ng1624);
  assign n7725 = Ng1624 | Ng1657 | ~Ng1612;
  assign n7726 = (n8207 | ~Ng1620) & (~Ng1600 | n8438);
  assign n7727 = n7725 & n7726 & (Ng1648 | n7724);
  assign n7728 = n6815 | ~Ng1677;
  assign n7729 = (Pg35 | ~Ng1657) & (n7727 | n8378);
  assign n7730 = (Pg35 & ~n8771) | (~Ng1472 & (~Pg35 | ~n8771));
  assign n7731 = ~Pg35 | n5170;
  assign n7732 = n8335 | ~Ng1256 | n8005;
  assign n7733 = Pg35 | ~Ng1252;
  assign n7734 = (Pg35 & ~n8779) | (~Ng1129 & (~Pg35 | ~n8779));
  assign n7735 = ~Pg35 | n4887;
  assign n7736 = n8341 | ~Ng911 | n8014;
  assign n7737 = Pg35 | ~Ng907;
  assign n7738 = ~Ng847 | ~Ng812;
  assign n7739 = n7738 & (Ng837 | ~Ng847);
  assign n7740 = ~n7739 | ~n9326 | Ng723;
  assign n7741 = ~Ng723 | n7904 | n9326;
  assign n7742 = ~n6091_1 ^ Ng739;
  assign n7743 = ~Pg35 | n8180;
  assign n7744 = ~Ng699 | ~Ng681 | n8465 | Ng645 | n8466 | Ng650;
  assign n7745 = Ng703 & (n7744 | ~n8122);
  assign n7746 = n9327 | ~n7745 | Ng714;
  assign n7747 = ~n9327 | n7751 | ~Ng714;
  assign n7748 = ~n8467 | ~n7745 | Ng676;
  assign n7749 = n8467 | n7751 | ~Ng676;
  assign n7750 = ~n8122 ^ Ng671;
  assign n7751 = ~Pg35 | ~n7745;
  assign n7752 = ~Ng586 | ~n7754 | n8183;
  assign n7753 = Pg35 | ~Ng572;
  assign n7754 = ~Ng572 | n7831;
  assign n7755 = ~Pg35 | n8468;
  assign n7756 = n9328 & (~Pg35 | ~Ng490 | n8470);
  assign n7757 = Ng417 | n9329 | n8027;
  assign n7758 = ~Pg35 | ~n7976;
  assign n7759 = n6500 | ~Ng5011;
  assign n7760 = n6506 | ~Ng4826;
  assign n7761 = n6512_1 | ~Ng4831;
  assign n7762 = (n7791 | ~Ng4821) & (n7524 | n8322);
  assign n7763 = ~\[4427]  | n6520;
  assign n7764 = (n7578 & Ng4049) | (n6525 & (n7578 | ~Ng4049));
  assign n7765 = (n7587 & (~Ng4045 | n7590)) | (Ng4045 & n7590);
  assign n7766 = ~Ng4961 & (~n5927 | (n7764 & n7765));
  assign n7767 = n6529 | ~Ng4961;
  assign n7768 = n8211 | n5888;
  assign n7769 = (~Ng3694 & n8455) | (n8327 & (Ng3694 | n8455));
  assign n7770 = (n7619 & Ng3698) | (n6531_1 & (n7619 | ~Ng3698));
  assign n7771 = ~Ng4950 & (~n5889 | (n7769 & n7770));
  assign n7772 = n6535 | ~Ng4950;
  assign n7773 = n8211 | n5907;
  assign n7774 = n8211 | Ng4975 | Ng4899;
  assign n7775 = ~Pg35 | n5908;
  assign n7776 = (n7423 & (~Ng6732 | n7426)) | (Ng6732 & n7426);
  assign n7777 = (n7414 & Ng6736) | (n6496 & (n7414 | ~Ng6736));
  assign n7778 = ~Ng4894 & (~n5884_1 | (n7776 & n7777));
  assign n7779 = n6500 | ~Ng4894;
  assign n7780 = (~Ng6386 & n7457) | (n7454 & (Ng6386 | n7457));
  assign n7781 = (n7445 & Ng6390) | (n6502_1 & (n7445 | ~Ng6390));
  assign n7782 = ~Ng4771 & (~n5952 | (n7780 & n7781));
  assign n7783 = n6506 | ~Ng4771;
  assign n7784 = n8209 | n5939;
  assign n7785 = (n7485 & (~Ng6040 | n7488)) | (Ng6040 & n7488);
  assign n7786 = (n7476 & Ng6044) | (n6508 & (n7476 | ~Ng6044));
  assign n7787 = ~Ng4760 & (~n5940 | (n7785 & n7786));
  assign n7788 = n6512_1 | ~Ng4760;
  assign n7789 = n8209 | n5874_1;
  assign n7790 = n8209 | Ng4785 | Ng4709;
  assign n7791 = ~Pg35 | n5876;
  assign n7792 = (n8192 & Ng5352) | (n6516 & (n8192 | ~Ng5352));
  assign n7793 = (n7545 & (~Ng5348 | n7548)) | (Ng5348 & n7548);
  assign n7794 = ~Ng4704 & (~n4151_1 | (n7792 & n7793));
  assign n7795 = n6520 | ~Ng4704;
  assign n7796 = n5951 | n8209;
  assign n7797 = Pg35 & (Ng4057 | Ng4064 | ~n8471);
  assign n7798 = Pg35 | ~Ng4119;
  assign n7799 = ~Pg35 | ~n7800 | ~Ng4122;
  assign n7800 = n8323 | ~n8471;
  assign n7801 = ~Pg35 | ~Ng4145;
  assign n7802 = Pg35 | ~Ng4116;
  assign n7803 = ~Ng4119 | ~Pg35 | n8472;
  assign n7804 = Pg35 | ~Ng4112;
  assign n7805 = ~Ng4116 | ~Pg35 | n8473;
  assign n7806 = n9336 & (~Pg35 | ~Ng4076 | ~n7807);
  assign n7807 = ~n8324 | ~Ng4082;
  assign n7808 = n6529 | ~Ng4035;
  assign n7809 = n6535 | ~Ng3684;
  assign n7810 = (n7775 | ~Ng3333) & (n7654 | n8328);
  assign n7811 = Pg35 | ~Ng2724;
  assign n7812 = n8256 ^ Ng2729;
  assign n7813 = n9337 & (~Pg35 | n6631 | ~Ng1345);
  assign n7814 = ~Pg35 | ~n8333;
  assign n7815 = ~Ng1252 | ~n7817 | n8005;
  assign n7816 = Pg35 | ~Ng1280;
  assign n7817 = n8334 | ~Ng1280;
  assign n7818 = n9338 & (~Pg35 | n6638_1 | ~Ng1002);
  assign n7819 = ~Pg35 | ~n8339;
  assign n7820 = ~Ng907 | ~n7822 | n8014;
  assign n7821 = Pg35 | ~Ng936;
  assign n7822 = n8340 | ~Ng936;
  assign n7823 = n8464 | ~n7739 | Ng827;
  assign n7824 = ~n8464 | n7904 | ~Ng827;
  assign n7825 = n7758 | ~Ng699;
  assign n7826 = ~Pg35 | n8474;
  assign n7827 = (n7826 | ~Ng681) & (~Ng650 | ~n8475);
  assign n7828 = ~n7986 & (~Ng703 | Ng714);
  assign n7829 = ~Ng572 | ~n7831 | n8183;
  assign n7830 = Pg35 | ~Ng568;
  assign n7831 = ~Ng568 | n7909;
  assign n7832 = Pg35 | ~Ng528;
  assign n7833 = ~n5934 ^ Ng482;
  assign n7834 = ~Pg35 | ~n8241;
  assign n7835 = n5881 | n5885;
  assign n7836 = n7835 & (n5918 | (n5881 & n5885));
  assign n7837 = ~n5905 & n5877 & ~n5902;
  assign n7838 = ~n8212 & (n5877 | (~n5902 & ~n5905));
  assign n7839 = Ng4531 & Ng4581;
  assign n7840 = Pg10306 & Pg35;
  assign n7841 = ~Pg35 | ~Ng4515 | ~Ng4521;
  assign n7842 = n7853 | Ng4392 | Ng4417;
  assign n7843 = (~Pg35 | n7842) & (~Ng4392 | ~n8479);
  assign n7844 = Ng4452 | Ng4438 | Ng4443 | Pg7245 | Pg7260;
  assign n7845 = Pg35 & (~Ng4392 | n7844);
  assign n7846 = ~Pg35 | Ng4392;
  assign n7847 = ~Pg35 | ~Ng4392 | n7844;
  assign n7848 = Pg35 | ~Ng4443;
  assign n7849 = ~Ng4438 | ~Pg35 | Ng4382;
  assign n7850 = Ng4401 ^ Ng4434;
  assign n7851 = Pg35 & (n7850 | (Ng4388 & ~Ng4430));
  assign n7852 = ~Pg35 | ~Ng4423;
  assign n7853 = Ng4411 | Ng4405 | Ng4375 | Pg7257 | Pg7243;
  assign n7854 = Pg35 & (~Ng4392 | n7853);
  assign n7855 = ~Ng4382 | ~n8479 | Ng4375;
  assign n7856 = ~Ng4375 | Ng4382 | ~n8479;
  assign n7857 = (n7842 & (Pg35 | ~Ng4388)) | (~Pg35 & ~Ng4388);
  assign n7858 = ~Pg35 | ~Ng4392 | n7853;
  assign n7859 = n7853 | n7846;
  assign n7860 = Pg35 | ~Ng4141;
  assign n7861 = ~n8324 ^ Ng4082;
  assign n7862 = (~n5995 | ~Ng2827) & (~n5996 | Ng2595);
  assign n7863 = (~n5995 | ~Ng2823) & (~n5996 | Ng2461);
  assign n7864 = (~n5995 | ~Ng2811) & (~n5996 | Ng2327);
  assign n7865 = (~n5995 | ~Ng2799) & (~n5996 | Ng2193);
  assign n7866 = (~n5995 | ~Ng2795) & (~n5996 | Ng2036);
  assign n7867 = (~n5995 | ~Ng2791) & (~n5996 | Ng1902);
  assign n7868 = (~n5995 | ~Ng2779) & (~n5996 | Ng1768);
  assign n7869 = (~n5995 | ~Ng2767) & (~n5996 | Ng1632);
  assign n7870 = ~n8255 | n7336 | ~Ng2724;
  assign n7871 = ~Ng2841 | Ng2724 | n8255;
  assign n7872 = Pg35 | ~Ng1437;
  assign n7873 = ~Pg35 | ~Ng1478 | n8481;
  assign n7874 = Pg35 | ~Ng1467;
  assign n7875 = ~Pg35 | ~Ng1472 | n8482;
  assign n7876 = ~Pg35 | ~Ng1448 | n8483;
  assign n7877 = Pg12923 & (Pg7946 | Pg19357 | Ng1333);
  assign n7878 = Ng1395 & n7877;
  assign n7879 = ~n5425 & (Ng1384 | ~Ng1351);
  assign n7880 = ~Ng1389 | ~Pg35 | n7879;
  assign n7881 = Ng1280 | n8334;
  assign n7882 = ~Ng1280 | n8005 | ~n8334;
  assign n7883 = Pg35 | ~Ng1094;
  assign n7884 = ~Pg35 | ~Ng1135 | n8486;
  assign n7885 = Pg35 | ~Ng1124;
  assign n7886 = ~Pg35 | ~Ng1129 | n8487;
  assign n7887 = ~Pg35 | ~Ng1105 | n8488;
  assign n7888 = Pg12919 & (Pg7916 | Pg19334 | Ng990);
  assign n7889 = (~Pg35 | ~Ng1061) & (~n7888 | ~Ng1052);
  assign n7890 = ~n4558 & (~Ng1008 | Ng1041);
  assign n7891 = ~Ng1046 | ~Pg35 | n7890;
  assign n7892 = Ng936 | n8340;
  assign n7893 = ~Ng936 | n8014 | ~n8340;
  assign n7894 = Pg35 & ~Ng890;
  assign n7895 = (n8492 | ~Ng872) & (~Ng446 | n8491);
  assign n7896 = (~Ng246 | n8491) & (~Pg14167 | n8492);
  assign n7897 = (~Ng269 | n8491) & (~Pg14147 | n8492);
  assign n7898 = (~Ng239 | n8491) & (~Pg14125 | n8492);
  assign n7899 = (~Ng262 | n8491) & (~Pg14096 | n8492);
  assign n7900 = (~Ng232 | n8491) & (~Pg14217 | n8492);
  assign n7901 = (~Ng255 | n8491) & (~Pg14201 | n8492);
  assign n7902 = (~Ng225 | n8491) & (~Pg14189 | n8492);
  assign n7903 = n8131 ^ Ng822;
  assign n7904 = ~Pg35 | ~n7739;
  assign n7905 = Pg35 & (~Ng847 | ~Ng843);
  assign n7906 = ~Pg35 | ~\[4435]  | n8122;
  assign n7907 = ~Ng568 | ~n7909 | n8183;
  assign n7908 = Pg35 | ~Ng562;
  assign n7909 = ~n5957 | ~Ng562 | n8182;
  assign n7910 = ~Ng355 & (~Pg35 | (Ng351 & ~Ng333));
  assign n7911 = ~\[4436]  & ~Ng351;
  assign n7912 = ~Ng305 & (Ng311 | ~Ng324);
  assign n7913 = ~Pg35 | ~Ng336 | ~n8493;
  assign n7914 = Pg35 | ~Ng311;
  assign n7915 = ~Pg35 | n8493;
  assign n7916 = (Pg35 & (Ng329 | n9349)) | (~Ng329 & n9349);
  assign n7917 = (~Ng305 & Ng336) | (~Ng311 & (~Ng305 | ~Ng336));
  assign n7918 = ~Ng311 & ~Ng305;
  assign n7919 = (~Ng6537 | ~n8381) & (n7404 | ~n8863);
  assign n7920 = Pg35 | ~Ng6509;
  assign n7921 = Ng6513 | ~Pg35 | n7404;
  assign n7922 = (~Ng6191 | ~n8386) & (n7435 | ~n8873);
  assign n7923 = Pg35 | ~Ng6163;
  assign n7924 = Ng6167 | ~Pg35 | n7435;
  assign n7925 = (~Ng5845 | ~n8390) & (n7466 | ~n8883);
  assign n7926 = Pg35 | ~Ng5817;
  assign n7927 = Ng5821 | ~Pg35 | n7466;
  assign n7928 = (~Ng5499 | ~n8394) & (n7497 | ~n8893);
  assign n7929 = Pg35 | ~Ng5471;
  assign n7930 = Ng5475 | ~Pg35 | n7497;
  assign n7931 = (~Ng5152 | n7934) & (n7527 | ~n8903);
  assign n7932 = Pg35 | ~Ng5124;
  assign n7933 = Ng5128 | ~Pg35 | n7527;
  assign n7934 = ~Pg35 | ~n7527;
  assign n7935 = Pg35 | ~Ng5097;
  assign n7936 = ~Ng5097 | ~n8494;
  assign n7937 = Pg35 | ~Ng5092;
  assign n7938 = ~Pg35 | ~Ng5097 | n8494;
  assign n7939 = Ng5092 & Pg35;
  assign n7940 = ~Ng5077 | ~Pg35 | Ng5073;
  assign n7941 = Pg35 & ~Ng5084;
  assign n7942 = Ng4098 & ~Ng4093;
  assign n7943 = n7942 & Ng4076 & ~Ng4064 & n6260_1 & Ng4087 & ~Ng4057;
  assign n7944 = ~Ng2841 | n8323 | Ng4141;
  assign n7945 = ~Ng4141 | n7566 | ~n8323;
  assign n7946 = (Ng4064 & (Pg35 | ~Ng4072)) | (~Pg35 & ~Ng4072);
  assign n7947 = n7946 & n6521;
  assign n7948 = (~Ng3845 | ~n8401) & (n7568 | ~n8919);
  assign n7949 = Pg35 | ~Ng3817;
  assign n7950 = Ng3821 | ~Pg35 | n7568;
  assign n7951 = (~Ng3494 | ~n8405) & (n7599 | ~n8929);
  assign n7952 = Pg35 | ~Ng3466;
  assign n7953 = Ng3470 | ~Pg35 | n7599;
  assign n7954 = (n7628 | ~n8939) & (~n8409 | ~Ng3143);
  assign n7955 = Pg35 | ~Ng3115;
  assign n7956 = Ng3119 | ~Pg35 | n7628;
  assign n7957 = ~Ng2715 | Ng2719;
  assign n7958 = (Pg35 & n8370) | (~Ng2715 & (~Pg35 | n8370));
  assign n7959 = n7957 & n6333 & n7958;
  assign n7960 = Pg35 | ~Ng1484;
  assign n7961 = ~Pg35 | ~Ng1300 | n8496;
  assign n7962 = ~Pg35 | ~n5425 | ~Ng1384;
  assign n7963 = n8484 | Ng1384 | n5425;
  assign n7964 = ~Ng1361 | ~Ng1373;
  assign n7965 = ~n8484 & (~n6631 | (n7964 & ~n9355));
  assign n7966 = Pg35 & (~Pg12923 | Ng1266);
  assign n7967 = Ng1249 | n8005;
  assign n7968 = Pg35 | ~Ng1141;
  assign n7969 = ~Pg35 | ~Ng956 | n8498;
  assign n7970 = ~Pg35 | ~n4558 | ~Ng1041;
  assign n7971 = n8489 | Ng1041 | n4558;
  assign n7972 = ~Ng1018 | ~Ng1030;
  assign n7973 = ~n8489 & (~n6638_1 | (n7972 & ~n9360));
  assign n7974 = Pg35 & (~Pg12919 | Ng921);
  assign n7975 = Ng904 | n8014;
  assign n7976 = ~Ng370 | ~Ng385 | n7993;
  assign n7977 = Pg35 & (~n7739 | Ng832 | n7976);
  assign n7978 = n8533 | n8534;
  assign n7979 = n8138 | n8139;
  assign n7980 = n5960 | ~Ng732;
  assign n7981 = ~n8123 | ~Pg35 | n7986;
  assign n7982 = Pg35 | ~Ng691;
  assign n7983 = ~Pg35 | ~n7986;
  assign n7984 = n5957 ^ Ng562;
  assign n7985 = n7984 & (~Ng632 | ~Ng626) & ~n8183;
  assign n7986 = ~Ng358 | ~Ng385 | Ng376;
  assign n7987 = Pg35 & (n7986 | ~n8468);
  assign n7988 = (~n7983 & ~Ng504) | (~Ng499 & (n7983 | ~Ng504));
  assign n7989 = (~Ng246 | n8499) & (~n8500 | ~Ng460);
  assign n7990 = (~Ng446 | n8499) & (~Ng182 | ~n8500);
  assign n7991 = Pg35 | ~Ng376;
  assign n7992 = ~Pg35 | ~Ng385 | ~n7993;
  assign n7993 = ~Ng376 | ~Ng358;
  assign n7994 = Ng4322 | ~Pg35 | Ng4332 | Ng4311 | n8191;
  assign n7995 = Ng4340 | ~Ng4643;
  assign n7996 = Ng4593 | n8232 | Ng4584 | Ng4608 | ~Ng4633 | Ng4616 | n7994 | Ng4601;
  assign n7997 = ~Pg35 | Ng4258;
  assign n7998 = n7997 & (~Pg35 | Ng4264);
  assign n7999 = n7998 & (~Pg35 | Ng4269);
  assign n8000 = Pg35 & (~Ng4264 | Ng4273 | ~Ng4258);
  assign n8001 = (Ng2715 & (Pg35 | ~Ng2712)) | (~Pg35 & ~Ng2712);
  assign n8002 = n8001 & n6333;
  assign n8003 = Pg35 | ~Ng1548;
  assign n8004 = ~Pg35 | ~Ng1564 | n8495;
  assign n8005 = ~Pg35 | ~Pg12923;
  assign n8006 = Ng1548 & Pg35;
  assign n8007 = n8140 & ~n5425 & ~n5965;
  assign n8008 = n8007 & Pg35;
  assign n8009 = Pg35 | ~Ng1589;
  assign n8010 = ~Pg10527 | ~Pg35 | Pg17423;
  assign n8011 = Pg35 & ~Pg12923;
  assign n8012 = Pg35 | ~Ng1205;
  assign n8013 = ~Pg35 | ~Ng1221 | n8497;
  assign n8014 = ~Pg35 | ~Pg12919;
  assign n8015 = Ng1205 & Pg35;
  assign n8016 = n8141 & n5036_1;
  assign n8017 = n8016 & Pg35;
  assign n8018 = Pg35 | ~Ng1246;
  assign n8019 = ~Pg10500 | ~Pg35 | Pg17400;
  assign n8020 = Pg35 & ~Pg12919;
  assign n8021 = Pg35 & n7738 & (~Ng832 | ~Ng827);
  assign n8022 = ~n7976 & Ng847;
  assign n8023 = Ng703 & (~Pg35 | (~Ng837 & n8022));
  assign n8024 = n7758 & (~Pg35 | (Ng837 & ~n7738));
  assign n8025 = (Pg35 & (Ng847 | n9398)) | (~Ng847 & n9398);
  assign n8026 = Ng691 & ~Ng542;
  assign n8027 = ~Pg35 | n7976;
  assign n8028 = (n7758 | ~Ng475) & (n8027 | ~Ng246);
  assign n8029 = (n7758 | ~Ng433) & (n8027 | ~Ng269);
  assign n8030 = n7758 | ~Ng392;
  assign n8031 = ~Ng854 | Ng703 | n8027;
  assign n8032 = Pg35 & (Ng4269 | ~Ng4258);
  assign n8033 = Ng4264 & Pg35;
  assign n8034 = ~Ng4349 | n8063;
  assign n8035 = Pg35 & n8034;
  assign n8036 = ~n8126 & ~Ng2988;
  assign n8037 = ~Ng4564 | ~Ng4555 | ~Ng4561 | ~Ng4558;
  assign n8038 = n8037 & ~Ng2988;
  assign n8039 = Pg35 & ~Ng2667;
  assign n8040 = Pg35 & ~Ng2527;
  assign n8041 = Pg35 & ~Ng2399;
  assign n8042 = Pg35 & ~Ng2265;
  assign n8043 = Pg35 & ~Ng2102;
  assign n8044 = Pg35 & ~Ng1968;
  assign n8045 = Pg35 & ~Ng1840;
  assign n8046 = Pg35 & ~Ng1706;
  assign n8047 = n8115 | ~Ng1542;
  assign n8048 = Pg35 & n8047;
  assign n8049 = n8117 | ~Ng1199;
  assign n8050 = Pg35 & n8049;
  assign n8051 = Pg35 & ~Ng6533;
  assign n8052 = Pg35 & ~Ng6187;
  assign n8053 = Pg35 & ~Ng5841;
  assign n8054 = Pg35 & ~Ng5495;
  assign n8055 = Pg35 & ~Ng5148;
  assign n8056 = Pg35 & ~Ng3841;
  assign n8057 = Pg35 & ~Ng3490;
  assign n8058 = Pg35 & ~Ng3139;
  assign n8059 = ~n6252 & (Pg35 | ~Ng385);
  assign n1117 = ~n8059;
  assign n8061 = ~Ng4593 | ~n8234;
  assign n8062 = Ng4332 & Ng4322 & n8233;
  assign n8063 = ~Ng4628 | n8232;
  assign n8064 = Ng4349 ^ n8063;
  assign n8065 = ~Ng4688 | n8208;
  assign n8066 = Ng2599 | ~Ng2629;
  assign n8067 = ~n8066 ^ Ng112;
  assign n8068 = Ng2465 | ~Ng2495;
  assign n8069 = ~n8068 ^ Ng112;
  assign n8070 = Ng2331 | ~Ng2361;
  assign n8071 = ~n8070 ^ Ng112;
  assign n8072 = Ng2197 | ~Ng2227;
  assign n8073 = ~n8072 ^ Ng112;
  assign n8074 = Ng2040 | ~Ng2070;
  assign n8075 = ~n8074 ^ Ng112;
  assign n8076 = Ng1906 | ~Ng1936;
  assign n8077 = ~n8076 ^ Ng112;
  assign n8078 = Ng1772 | ~Ng1802;
  assign n8079 = ~n8078 ^ Ng112;
  assign n8080 = Ng1636 | ~Ng1668;
  assign n8081 = ~n8080 ^ Ng112;
  assign n8082 = ~Ng1339 ^ Ng1322;
  assign n8083 = ~Ng996 ^ Ng979;
  assign n8084 = Ng2610 | ~Ng2619;
  assign n8085 = Ng110 ^ n8084;
  assign n8086 = Ng2476 | ~Ng2485;
  assign n8087 = Ng110 ^ n8086;
  assign n8088 = Ng2342 | ~Ng2351;
  assign n8089 = Ng110 ^ n8088;
  assign n8090 = Ng2208 | ~Ng2217;
  assign n8091 = Ng110 ^ n8090;
  assign n8092 = Ng2051 | ~Ng2060;
  assign n8093 = Ng110 ^ n8092;
  assign n8094 = Ng1917 | ~Ng1926;
  assign n8095 = Ng110 ^ n8094;
  assign n8096 = Ng1783 | ~Ng1792;
  assign n8097 = Ng110 ^ n8096;
  assign n8098 = Ng1648 | ~Ng1657;
  assign n8099 = Ng110 ^ n8098;
  assign n8100 = Pg35 & Ng5471;
  assign n8101 = (n6884 | n6883) & (n8100 | n6887);
  assign n8102 = n6883 | n8100 | n6884;
  assign n8103 = n6890 & n8102;
  assign n8104 = n6889 & (n6890 | n8102);
  assign n8105 = Pg35 & Ng3466;
  assign n8106 = ~Ng2735 | n7657;
  assign n8107 = ~Ng2652 ^ Ng2648;
  assign n8108 = ~Ng2514 ^ Ng2518;
  assign n8109 = ~Ng2384 ^ Ng2380;
  assign n8110 = ~Ng2250 ^ Ng2246;
  assign n8111 = ~Ng2089 ^ Ng2093;
  assign n8112 = ~Ng1955 ^ Ng1959;
  assign n8113 = ~Ng1821 ^ Ng1825;
  assign n8114 = ~Ng1687 ^ Ng1691;
  assign n8115 = ~Pg7946 | ~Ng1526 | n5963 | Ng1514;
  assign n8116 = n8115 ^ Ng1542;
  assign n8117 = ~Pg7916 | Ng1171 | ~Ng1183 | n8439;
  assign n8118 = n8117 ^ Ng1199;
  assign n8119 = ~n5935 ^ n7558;
  assign n8120 = ~n5949 ^ n7563;
  assign n8121 = ~Ng4076 | n7807;
  assign n8122 = ~Ng504 & Ng499 & n5933 & ~n7976;
  assign n8123 = Ng691 | ~Ng703 | n7744;
  assign n8124 = (n7828 | ~Ng691) & (n7986 | n8123);
  assign n8125 = (n5918 | n7835) & (n5865 | n7836);
  assign n8126 = Ng4489 & Ng4483 & Ng4486 & Ng4492;
  assign n8127 = ~Ng4521 & ~n9340 & (n8126 | Ng4527);
  assign n8128 = ~n5958 & (~Ng1536 | (~n8047 & Ng1413));
  assign n8129 = ~n7878 ^ Ng1404;
  assign n8130 = ~n5959 & (~Ng1193 | (~n8049 & Ng1070));
  assign n8131 = ~Ng817 | ~Ng832 | n7976;
  assign n8132 = n8122 & (Ng728 | (Ng661 & Pg35));
  assign n8133 = n8495 & Ng1564;
  assign n8134 = ~n8133 ^ Ng1559;
  assign n8135 = n8497 & Ng1221;
  assign n8136 = ~n8135 ^ Ng1216;
  assign n8137 = Ng232 ^ Ng255;
  assign n8138 = ~Ng246 ^ Ng269;
  assign n8139 = ~Ng239 ^ Ng262;
  assign n8140 = Ng1322 ^ Ng1579;
  assign n8141 = Ng1236 ^ Ng979;
  assign n8142 = ~Pg54 | Pg57 | Pg56 | Pg53 | Ng55;
  assign n8143 = ~Ng50 | Ng16;
  assign n8144 = Ng46 & Ng48 & Ng45 & Ng8 & ~Ng52;
  assign n8145 = Ng45 | Ng46 | Ng8;
  assign n8146 = Ng52 | ~Ng51 | n8145;
  assign n8147 = Ng48 | n8146;
  assign n8148 = Ng50 | ~Ng16;
  assign n8149 = n8147 | n8148;
  assign n8150 = Ng16 | Ng50;
  assign n8151 = ~Ng52 | Ng48 | n8145;
  assign n3827_1 = ~n8142;
  assign n8153 = Pg53 | ~n8142;
  assign n8154 = n8145 | Ng51 | Ng52;
  assign n8155 = n8142 | n6080;
  assign n8156 = Ng48 | n8154;
  assign n8157 = n8151 | Ng51 | n8143;
  assign n8158 = n8157 & n6063 & n6027_1;
  assign n8159 = n8150 | n8156;
  assign n8160 = n8148 | n8156;
  assign n8161 = n8142 | n8160;
  assign n8162 = n8143 | n8147;
  assign n8163 = n8142 | n8162;
  assign n8164 = ~Ng48 | n8143;
  assign n8165 = n8146 | n8164;
  assign n8166 = n8142 | n8165;
  assign n8167 = n8142 | Ng48 | ~Ng50 | ~Ng16;
  assign n8168 = n8146 | n8167;
  assign n8169 = n8154 | n8167;
  assign n8170 = n8154 | n8164;
  assign n8171 = n8142 | n8170;
  assign n8172 = Ng51 | n8145 | ~Ng52 | n8164;
  assign n8173 = n8142 | n8172;
  assign n8174 = n8148 | ~n8144 | Ng51;
  assign n8175 = Ng1291 | n8161;
  assign n8176 = Ng947 | n8163;
  assign n8177 = n6087 | n6088;
  assign n8178 = Ng4322 ^ Pg72;
  assign n8179 = Ng4332 ^ Pg73;
  assign n8180 = Pg11678 & ~Ng736;
  assign n8181 = Ng370 | ~Ng385 | n7993;
  assign n8182 = Pg9048 & ~Ng559;
  assign n8183 = ~Pg35 | n8182;
  assign n8184 = Ng490 ^ Pg73;
  assign n8185 = Ng482 ^ Pg72;
  assign n8186 = Ng518 | n5931;
  assign n8187 = n5931 | ~Ng518;
  assign n8188 = ~Ng4349 | Ng4358;
  assign n8189 = ~Ng3352 | ~Ng3288;
  assign n8190 = Ng4349 | ~Ng4358;
  assign n8191 = Ng4358 | Ng4349;
  assign n8192 = ~Ng5357 | ~Ng5297;
  assign n8193 = Ng2759 ^ Pg72;
  assign n8194 = Ng2763 ^ Pg73;
  assign n8195 = n8193 | n8194;
  assign n8196 = n8195 | ~Ng2756 | Ng2748;
  assign n8197 = ~Ng2208 | Ng2217;
  assign n8198 = ~Ng2741 | Ng2756 | Ng2748;
  assign n8199 = ~Ng1783 | Ng1792;
  assign n8200 = ~Ng2748 | n8195;
  assign n8201 = ~Ng2051 | Ng2060;
  assign n8202 = ~Ng1917 | Ng1926;
  assign n8203 = ~Ng2476 | Ng2485;
  assign n8204 = ~Ng2342 | Ng2351;
  assign n8205 = ~Ng2610 | Ng2619;
  assign n8206 = ~Ng2741 & ~Ng2756 & ~Ng2748;
  assign n8207 = ~Ng1648 | Ng1657;
  assign n8208 = ~Ng4669 | ~Ng4659 | ~Ng4653;
  assign n8209 = ~Ng4793 | ~Ng4776 | Ng4801;
  assign n8210 = ~Ng4859 | ~Ng4843 | ~Ng4849;
  assign n8211 = ~Ng4983 | ~Ng4966 | Ng4991;
  assign n8212 = n7835 | n5865 | n5918;
  assign n8213 = Pg35 & Ng6509;
  assign n8214 = n8102 | n5880 | n6890 | n8105 | n6889 | n8213;
  assign n8215 = ~n8212 & ~n5906 & ~n5905 & n5877 & ~n5902;
  assign n8216 = ~Ng3171 | ~Ng3179;
  assign n8217 = ~Ng6219 | ~Ng6227;
  assign n8218 = ~Ng4098 & Ng4093;
  assign n8219 = ~Ng3873 | ~Ng3881;
  assign n8220 = Ng4098 & Ng4093;
  assign n8221 = ~Ng5527 | ~Ng5535;
  assign n8222 = ~Ng6565 | ~Ng6573;
  assign n8223 = ~Ng5873 | ~Ng5881;
  assign n8224 = ~Ng3522 | ~Ng3530;
  assign n8225 = ~Ng5180 | ~Ng5188;
  assign n8226 = Ng4108 ^ Pg72;
  assign n8227 = Ng4104 ^ Pg73;
  assign n8228 = n6126 & ~n8251;
  assign n8229 = ~Ng4878 | ~Ng4843;
  assign n8230 = n8065 & ~n8253;
  assign n8231 = ~Ng4688 | ~Ng4653;
  assign n8232 = ~Ng4340 | ~Ng4621 | Ng4639;
  assign n8233 = ~n8034 & Ng4358;
  assign n8234 = Ng4584 & n8062;
  assign n8235 = ~Pg35 | n6216_1;
  assign n8236 = Ng4311 & n8233;
  assign n8237 = n5924 | Ng4818 | \[4661] ;
  assign n8238 = ~n8237 & Ng71;
  assign n8239 = n5924 | Ng4818 | \[4661] ;
  assign n8240 = (~Ng278 & n4385) | (~n4384 & (Ng278 | n4385));
  assign n8241 = n8240 & ~n5962 & Ng691;
  assign n8242 = Ng287 & Ng283 & n8241;
  assign n8243 = ~n8242 | ~Ng291;
  assign n8244 = ~Ng294 | n8243;
  assign n8245 = ~Ng298 | n8244;
  assign n8246 = ~Ng691 | n5962 | n6300;
  assign n8247 = n4520 & Ng146 & ~n8246;
  assign n8248 = Ng164 & n8247;
  assign n8249 = ~n8248 | ~Ng150;
  assign n8250 = ~Ng153 | n8249;
  assign n8251 = Ng63 & n5966 & ~n6124;
  assign n8252 = ~n6316 & Ng4966;
  assign n8253 = Ng63 & n5966 & ~n6090;
  assign n8254 = ~n6327 & Ng4776;
  assign n8255 = ~Ng2715 | ~Ng2719;
  assign n8256 = ~Ng2724 | n8255;
  assign n8257 = n8106 | ~Ng2741;
  assign n8258 = ~Ng2748 | n8257;
  assign n8259 = ~Ng1322 | Ng1564 | Ng1548 | ~Ng1404 | Ng1559 | Ng1554;
  assign n8260 = ~Ng2629 & ~Ng2555;
  assign n8261 = ~n8260 | ~n8263;
  assign n8262 = n8261 & Pg35;
  assign n8263 = n5911 | ~n5999;
  assign n8264 = Ng2599 & ~Ng2555;
  assign n8265 = n8263 & n8264;
  assign n8266 = ~n8263 | ~Ng2555;
  assign n8267 = ~Ng2495 & ~Ng2421;
  assign n8268 = ~n8267 | ~n8270;
  assign n8269 = n8268 & Pg35;
  assign n8270 = n5872 | ~n6001;
  assign n8271 = Ng2465 & ~Ng2421;
  assign n8272 = n8270 & n8271;
  assign n8273 = ~n8270 | ~Ng2421;
  assign n8274 = ~Ng2361 & ~Ng2287;
  assign n8275 = ~n8274 | ~n8277;
  assign n8276 = n8275 & Pg35;
  assign n8277 = n5910 | ~n6011;
  assign n8278 = Ng2331 & ~Ng2287;
  assign n8279 = n8277 & n8278;
  assign n8280 = ~n8277 | ~Ng2287;
  assign n8281 = ~Ng2227 & ~Ng2153;
  assign n8282 = ~n8281 | ~n8284;
  assign n8283 = n8282 & Pg35;
  assign n8284 = n5873 | ~n6007;
  assign n8285 = ~Ng2227 | ~n8284;
  assign n8286 = Ng2197 & ~Ng2153;
  assign n8287 = n8284 & n8286;
  assign n8288 = ~Ng979 | Ng1221 | Ng1205 | Ng1211 | ~Ng1061 | Ng1216;
  assign n8289 = ~Ng2070 & ~Ng1996;
  assign n8290 = ~n8289 | ~n8292;
  assign n8291 = n8290 & Pg35;
  assign n8292 = n5921 | ~n6003;
  assign n8293 = ~Ng2070 | ~n8292;
  assign n8294 = Ng2040 & ~Ng1996;
  assign n8295 = n8292 & n8294;
  assign n8296 = ~Ng1936 & ~Ng1862;
  assign n8297 = ~n8296 | ~n8299;
  assign n8298 = n8297 & Pg35;
  assign n8299 = n5887 | ~n6005;
  assign n8300 = ~Ng1936 | ~n8299;
  assign n8301 = Ng1906 & ~Ng1862;
  assign n8302 = n8299 & n8301;
  assign n8303 = ~Ng1802 & ~Ng1728;
  assign n8304 = ~n8303 | ~n8306;
  assign n8305 = n8304 & Pg35;
  assign n8306 = n5894 | ~n5997;
  assign n8307 = Ng1772 & ~Ng1728;
  assign n8308 = n8306 & n8307;
  assign n8309 = ~n8306 | ~Ng1728;
  assign n8310 = ~Ng1592 & ~Ng1668;
  assign n8311 = ~n8310 | ~n8313;
  assign n8312 = n8311 & Pg35;
  assign n8313 = n4162 | ~n6009;
  assign n8314 = ~Ng1636 | ~n8313;
  assign n8315 = ~Ng1592 | ~n8313;
  assign n8316 = Ng4801 | Ng4793 | ~Ng4776;
  assign n8317 = Ng4991 | Ng4983 | ~Ng4966;
  assign n8318 = n5966 & Ng93;
  assign n8319 = n6124 | ~n8318;
  assign n8320 = n6090 | ~n8318;
  assign n8321 = ~Ng5703 | Ng5644;
  assign n8322 = ~Pg35 | ~n5876;
  assign n8323 = ~Ng4057 | ~Ng4064;
  assign n8324 = ~n8323 & Ng4141;
  assign n8325 = ~Ng4087 | n8121;
  assign n8326 = ~Ng4093 | n8325;
  assign n8327 = Ng3703 | ~Ng3639;
  assign n8328 = ~Pg35 | ~n5908;
  assign n8329 = Pg35 & n5966;
  assign n8330 = n5966 & Ng112;
  assign n8331 = n8082 | Ng1351;
  assign n8332 = ~n8082 | n7964 | ~Ng1351;
  assign n8333 = ~n9355 & n8332 & ~Ng1312 & n8331;
  assign n8334 = ~Pg12923 | ~Ng1266 | ~Ng1249;
  assign n8335 = Ng1252 & ~n7817;
  assign n8336 = Ng1259 & ~n7384;
  assign n8337 = n8083 | Ng1008;
  assign n8338 = ~n8083 | ~Ng1008 | n7972;
  assign n8339 = ~n9360 & n8338 & ~Ng969 & n8337;
  assign n8340 = ~Pg12919 | ~Ng921 | ~Ng904;
  assign n8341 = Ng907 & ~n7822;
  assign n8342 = Ng914 & ~n7394;
  assign n8343 = Ng43 & ~n5947 & n5966;
  assign n8344 = ~Ng4087 & n8343;
  assign n4287_1 = Pg35 & Ng6573;
  assign n8346 = ~Ng6565 | Ng6573;
  assign n8347 = Ng4087 & n8343;
  assign n8348 = ~Ng6219 | Ng6227;
  assign n1064_1 = Pg35 & Ng5881;
  assign n8350 = ~Ng5873 | Ng5881;
  assign n8351 = ~Ng5527 | Ng5535;
  assign n8352 = ~Ng5180 | Ng5188;
  assign n8353 = ~Ng5029 | ~Ng5016 | ~Ng5062;
  assign n8354 = ~Ng5033 | n8353 | ~Ng5037;
  assign n8355 = ~Ng5022 | Ng5029 | Ng5016;
  assign n8356 = n8355 | Ng5033 | Ng5037;
  assign n8357 = n8356 | Ng5046 | Ng5041;
  assign n8358 = Ng5057 & ~Ng5046 & Ng5022;
  assign n8359 = Ng5062 & Ng5046 & ~Ng5057;
  assign n8360 = n8358 & Pg84 & ~Ng5041;
  assign n8361 = n8359 & ~Pg84 & Ng5052;
  assign n8362 = n8358 & ~Pg84 & ~Ng5052;
  assign n8363 = Pg84 & Ng5041 & n8359;
  assign n8364 = n8360 | n8361 | n8362 | n8363;
  assign n8365 = ~Ng3873 | Ng3881;
  assign n8366 = ~Ng3522 | Ng3530;
  assign n8367 = ~Ng3171 | Ng3179;
  assign n8368 = n5966 & Ng110;
  assign n8369 = ~Pg35 | ~n5920;
  assign n8370 = Ng2715 | ~Ng2719;
  assign n8371 = ~Pg35 | ~n5919;
  assign n8372 = ~Pg35 | ~n5925;
  assign n8373 = Ng2719 | Ng2715;
  assign n8374 = ~Pg35 | ~n5878;
  assign n8375 = ~Pg35 | ~n5916;
  assign n8376 = ~Pg35 | ~n5899;
  assign n8377 = ~Pg35 | ~n5941;
  assign n8378 = ~Pg35 | ~n5868;
  assign n8379 = n8356 & n8354;
  assign n8380 = Ng5062 | Ng5022;
  assign n8381 = n7404 & Pg35;
  assign n8382 = Ng4180 & ~Ng4284;
  assign n8383 = Ng6565 | ~Ng6573;
  assign n8384 = Ng6565 | Ng6573;
  assign n8385 = Ng6555 | Ng6549 | Ng6561;
  assign n8386 = n7435 & Pg35;
  assign n8387 = Ng6219 | ~Ng6227;
  assign n8388 = Ng6219 | Ng6227;
  assign n8389 = Ng6203 | Ng6215 | Ng6209;
  assign n8390 = n7466 & Pg35;
  assign n8391 = Ng5873 | ~Ng5881;
  assign n8392 = Ng5873 | Ng5881;
  assign n8393 = Ng5863 | Ng5857 | Ng5869;
  assign n8394 = n7497 & Pg35;
  assign n8395 = Ng5527 | ~Ng5535;
  assign n8396 = Ng5527 | Ng5535;
  assign n8397 = Ng5517 | Ng5511 | Ng5523;
  assign n8398 = Ng5180 | ~Ng5188;
  assign n8399 = Ng5180 | Ng5188;
  assign n8400 = Ng5170 | Ng5164 | Ng5176;
  assign n8401 = n7568 & Pg35;
  assign n8402 = Ng3873 | ~Ng3881;
  assign n8403 = Ng3873 | Ng3881;
  assign n8404 = Ng3857 | Ng3869 | Ng3863;
  assign n8405 = n7599 & Pg35;
  assign n8406 = Ng3522 | ~Ng3530;
  assign n8407 = Ng3522 | Ng3530;
  assign n8408 = Ng3512 | Ng3506 | Ng3518;
  assign n8409 = n7628 & Pg35;
  assign n8410 = Ng3171 | ~Ng3179;
  assign n8411 = Ng3171 | Ng3179;
  assign n8412 = Ng3161 | Ng3155 | Ng3167;
  assign n8413 = Ng2619 & n5920 & Ng2587;
  assign n8414 = Pg35 & n8413;
  assign n8415 = ~Ng2610 | Ng2587;
  assign n8416 = Ng2485 & n5919;
  assign n8417 = Ng2453 & n8416;
  assign n8418 = Pg35 & n8417;
  assign n8419 = ~Ng2476 | Ng2453;
  assign n8420 = Ng2351 & n5925 & Ng2319;
  assign n8421 = Pg35 & n8420;
  assign n8422 = ~Ng2342 | Ng2319;
  assign n8423 = Ng2217 & n5878 & Ng2185;
  assign n8424 = Pg35 & n8423;
  assign n8425 = ~Ng2208 | Ng2185;
  assign n8426 = Ng2060 & n5916;
  assign n8427 = Ng2028 & n8426;
  assign n8428 = Pg35 & n8427;
  assign n8429 = ~Ng2051 | Ng2028;
  assign n8430 = Ng1926 & n5899 & Ng1894;
  assign n8431 = Pg35 & n8430;
  assign n8432 = ~Ng1917 | Ng1894;
  assign n8433 = Ng1792 & n5941 & Ng1760;
  assign n8434 = Pg35 & n8433;
  assign n8435 = ~Ng1783 | Ng1760;
  assign n8436 = Ng1657 & n5868 & Ng1624;
  assign n8437 = Pg35 & n8436;
  assign n8438 = ~Ng1648 | Ng1624;
  assign n8439 = Ng996 & Ng1178 & ~Ng1189;
  assign n8440 = ~n5884_1 | n7430;
  assign n8441 = ~Pg35 | n8440;
  assign n8442 = ~n5952 | n7461;
  assign n8443 = ~Pg35 | n8442;
  assign n8444 = ~n5940 | n7492;
  assign n8445 = ~Pg35 | n8444;
  assign n8446 = ~n5876 | n7523;
  assign n8447 = ~Pg35 | n8446;
  assign n8448 = \[4415]  & Pg17577 & ~n8192;
  assign n8449 = ~n4151_1 | ~n8448;
  assign n8450 = ~Pg35 | n8449;
  assign n8451 = ~n5927 | n7594;
  assign n8452 = ~Pg35 | n8451;
  assign n8453 = ~n5889 | n7623;
  assign n8454 = ~Pg35 | n8453;
  assign n8455 = Ng3639 | Ng3703;
  assign n8456 = ~n5908 | n7653;
  assign n8457 = ~Pg35 | n8456;
  assign n8458 = Pg13272 & Ng1526 & ~Ng1514;
  assign n8459 = Ng1514 & Ng1526 & Pg13272;
  assign n8460 = Ng1514 & Pg13272 & ~Ng1526;
  assign n8461 = Ng1183 & Pg13259 & ~Ng1171;
  assign n8462 = Ng1183 & Ng1171 & Pg13259;
  assign n8463 = Pg13259 & Ng1171 & ~Ng1183;
  assign n8464 = n8131 | ~Ng822;
  assign n8465 = Ng661 ^ Ng728;
  assign n8466 = Ng655 ^ Ng718;
  assign n8467 = n8122 & Ng671;
  assign n8468 = ~Ng667 | Ng686;
  assign n8469 = Ng513 | n7986 | ~Ng518;
  assign n8470 = Ng482 & n5934;
  assign n8471 = ~Ng4076 & ~n6261 & n6260_1 & ~Ng4087;
  assign n8472 = n8471 & Ng4057 & ~Ng4064;
  assign n8473 = n8471 & ~Ng4057 & Ng4064;
  assign n8474 = n8181 | n8476 | n8477;
  assign n8475 = n8474 & Pg35;
  assign n8476 = ~Ng691 & (Ng411 | Ng424 | ~Ng417);
  assign n8477 = Ng691 & (Ng499 | Ng518);
  assign n8478 = n5091 & Pg35;
  assign n8479 = n7853 & Pg35;
  assign n8480 = Ng1442 & ~Ng1495;
  assign n8481 = Ng1437 & n8460 & n8480;
  assign n8482 = Ng1467 & n8459 & n8480;
  assign n8483 = Ng1454 & n8458 & n8480;
  assign n8484 = ~Pg35 | ~Ng1351;
  assign n8485 = Ng1099 & ~Ng1152;
  assign n8486 = Ng1094 & n8463 & n8485;
  assign n8487 = Ng1124 & n8462 & n8485;
  assign n8488 = Ng1111 & n8461 & n8485;
  assign n8489 = ~Pg35 | ~Ng1008;
  assign n8490 = ~Ng862 & Ng890 & ~Ng896;
  assign n8491 = ~Pg35 | n8490;
  assign n8492 = ~Pg35 | ~n8490;
  assign n8493 = (Ng324 & ~Ng305) | (~Ng311 & (~Ng324 | ~Ng305));
  assign n8494 = Ng5084 & Ng5092;
  assign n8495 = Ng1430 & Ng1548;
  assign n8496 = Ng1484 & n5170 & n8480;
  assign n8497 = Ng1087 & Ng1205;
  assign n8498 = Ng1141 & n4887 & n8485;
  assign n8499 = ~Pg35 | n8181;
  assign n8500 = n8181 & Pg35;
  assign n8501 = Pg8291 & Ng218;
  assign n8502 = Pg17688 & Pg17778 & Pg14828 & Pg12470;
  assign n8503 = ~Pg17760 | ~Pg17649 | ~Pg14779 | ~Pg12422;
  assign n8504 = Pg17607 & Pg17739 & Pg14738 & Pg12350;
  assign n8505 = Pg17580 & Pg17711 & Pg14694 & Pg12300;
  assign n8506 = ~Pg17674 | ~Pg17519 | ~Pg14662 | ~Pg12238;
  assign n8507 = ~Pg16775 | ~Pg16659 | ~Pg13966 | ~Pg11418;
  assign n8508 = ~Pg16744 | ~Pg16627 | ~Pg13926 | ~Pg11388;
  assign n8509 = ~Pg16718 | ~Pg16603 | ~Pg13895 | ~Pg11349;
  assign n8510 = n8133 & Ng1554;
  assign n8511 = n8135 & Ng1211;
  assign n8512 = ~n7430 ^ n7431;
  assign n8513 = n7461 ^ n7462;
  assign n8514 = ~n7492 ^ n7493;
  assign n8515 = ~n7523 ^ n7524;
  assign n8516 = n8448 ^ n7552;
  assign n8517 = ~n7594 ^ n7595;
  assign n8518 = ~n7623 ^ n7624;
  assign n8519 = ~n7653 ^ n7654;
  assign n8520 = Ng1319 | n5091;
  assign n8521 = ~Ng1448 ^ n8520;
  assign n8522 = ~Ng1300 ^ n8520;
  assign n8523 = ~Ng1472 ^ n8520;
  assign n8524 = ~Ng1478 ^ n8520;
  assign n8525 = ~n6128 | Ng976;
  assign n8526 = ~Ng1105 ^ n8525;
  assign n8527 = ~Ng956 ^ n8525;
  assign n8528 = ~Ng1129 ^ n8525;
  assign n8529 = ~Ng1135 ^ n8525;
  assign n6560 = Ng4534 ^ n7840;
  assign n4047_1 = Ng862 ^ n7894;
  assign n1777 = Ng5084 ^ n7939;
  assign n8533 = Ng246 ^ Ng269;
  assign n8534 = Ng239 ^ Ng262;
  assign n8535 = n5985 ^ n7980;
  assign n6452 = Ng1430 ^ n8006;
  assign n4627 = Ng1333 ^ n8008;
  assign n1087_1 = Ng1087 ^ n8015;
  assign n5768 = Ng990 ^ n8017;
  assign n8540 = ~Pg9019 ^ Ng4291;
  assign n8541 = ~Pg9019 ^ n8540;
  assign n8542 = ~Pg8839 ^ Ng4281;
  assign n8543 = ~Pg8839 ^ n8542;
  assign n8544 = ~n9153 & (Pg35 | ~Ng2980);
  assign n2483 = ~n8544;
  assign n8546 = (Pg35 & n9162) | (~Ng4366 & (~Pg35 | n9162));
  assign n800_1 = ~n8546;
  assign n8548 = ~n9164 & (Pg35 | ~Ng2955);
  assign n3760 = ~n8548;
  assign n8550 = ~n9166 & (Pg35 | ~Ng2941);
  assign n1112_1 = ~n8550;
  assign n8552 = ~n9168 & (Pg35 | ~Ng2927);
  assign n1372_1 = ~n8552;
  assign n8554 = ~n9169 & (Pg35 | ~Ng2965);
  assign n2423 = ~n8554;
  assign n8556 = ~n9171 & (Pg35 | ~Ng2917);
  assign n4244 = ~n8556;
  assign n8558 = ~n9172 & (Pg35 | ~Ng2902);
  assign n4460 = ~n8558;
  assign n8560 = ~n9174 & (Pg35 | ~Ng2970);
  assign n2946_1 = ~n8560;
  assign n8562 = Ng55 | Ng2980;
  assign n8563 = (Pg35 & ~n8562) | (~Ng2886 & (~Pg35 | ~n8562));
  assign n1552_1 = ~n8563;
  assign n8565 = ~Pg44 | Ng2890;
  assign n8566 = (Pg35 & ~n8565) | (~Ng2873 & (~Pg35 | ~n8565));
  assign n5633 = ~n8566;
  assign n8568 = Ng2946 | Ng2886;
  assign n8569 = (Pg35 & ~n8568) | (~Ng2878 & (~Pg35 | ~n8568));
  assign n1752 = ~n8569;
  assign n8571 = ~Pg91 | Ng2878;
  assign n8572 = (Pg35 & ~n8571) | (~Ng2882 & (~Pg35 | ~n8571));
  assign n3832_1 = ~n8572;
  assign n8574 = ~n9176 & (Pg35 | ~Ng2898);
  assign n3871_1 = ~n8574;
  assign n8576 = Ng2898 | ~n8215;
  assign n8577 = (Pg35 & ~n8576) | (~Ng2864 & (~Pg35 | ~n8576));
  assign n1664_1 = ~n8577;
  assign n8579 = Ng2864 | n8214;
  assign n8580 = (Pg35 & ~n8579) | (~Ng2856 & (~Pg35 | ~n8579));
  assign n3975 = ~n8580;
  assign n8582 = ~n9178 & (Pg35 | ~Ng2848);
  assign n5653 = ~n8582;
  assign n8584 = ~n9180 & (Pg35 | ~\[4433] );
  assign n2280_1 = ~n8584;
  assign n8586 = Ng4242 | Ng4300;
  assign n8587 = (~Pg35 & ~Ng4297) | (~n8586 & (Pg35 | ~Ng4297));
  assign n6646 = ~n8587;
  assign n8589 = Ng4176 | Ng4072;
  assign n8590 = (Pg35 & ~n8589) | (~Ng4172 & (~Pg35 | ~n8589));
  assign n4882 = ~n8590;
  assign n8592 = Ng1283 | Ng1277;
  assign n8593 = (Pg35 & ~n8592) | (~Ng1296 & (~Pg35 | ~n8592));
  assign n2111 = ~n8593;
  assign n8595 = Ng933 | Ng939;
  assign n8596 = (Pg35 & ~n8595) | (~Ng952 & (~Pg35 | ~n8595));
  assign n1247 = ~n8596;
  assign n8598 = Ng534 | Ng301;
  assign n8599 = (Pg35 & ~n8598) | (~Ng542 & (~Pg35 | ~n8598));
  assign n6536 = ~n8599;
  assign n8601 = ~Ng691 | Ng546;
  assign n8602 = (Pg35 & ~n8601) | (~Ng538 & (~Pg35 | ~n8601));
  assign n5956 = ~n8602;
  assign n8604 = Ng199 | Ng222;
  assign n8605 = (Pg35 & ~n8604) | (~\[4426]  & (~Pg35 | ~n8604));
  assign n3675 = ~n8605;
  assign n8607 = ~\[4435]  | Ng550;
  assign n8608 = (Pg35 & ~n8607) | (~Ng534 & (~Pg35 | ~n8607));
  assign n3927 = ~n8608;
  assign n8610 = (~Pg35 & ~Ng37) | (~\[4433]  & (Pg35 | ~Ng37));
  assign n6160 = ~n8610;
  assign n4667_1 = ~n9188;
  assign n5913_1 = ~n9189;
  assign n8614 = (~Pg35 & ~Ng550) | (~\[4426]  & (Pg35 | ~Ng550));
  assign n2793_1 = ~n8614;
  assign n8616 = ~n9190 & (Ng4878 | n6193 | ~Ng4843);
  assign n6260 = ~n8616;
  assign n8618 = ~n9191 & (Ng4688 | n6198 | ~Ng4653);
  assign n1868 = ~n8618;
  assign n8620 = (Pg35 & n9192) | (~Ng4643 & (~Pg35 | n9192));
  assign n4249 = ~n8620;
  assign n8622 = (n6254 & (Pg35 | ~Ng446)) | (~Pg35 & ~Ng446);
  assign n3775 = ~n8622;
  assign n8624 = (Pg35 & n9206) | (~Ng4961 & (~Pg35 | n9206));
  assign n4554 = ~n8624;
  assign n8626 = (Pg35 & n9208) | (~Ng4950 & (~Pg35 | n9208));
  assign n3548 = ~n8626;
  assign n8628 = (Pg35 & n9210) | (~Ng4894 & (~Pg35 | n9210));
  assign n2065_1 = ~n8628;
  assign n8630 = (Pg35 & n9212) | (~Ng4771 & (~Pg35 | n9212));
  assign n4909_1 = ~n8630;
  assign n8632 = (Pg35 & n9214) | (~Ng4760 & (~Pg35 | n9214));
  assign n1591_1 = ~n8632;
  assign n8634 = (Pg35 & n9216) | (~Ng4704 & (~Pg35 | n9216));
  assign n6201_1 = ~n8634;
  assign n8636 = (n8035 & Ng4358) | (~n8034 & (n8035 | ~Ng4358));
  assign n8637 = n9217 & (~Pg35 | n5968 | n8064);
  assign n5613_1 = ~n8637;
  assign n8639 = (Pg35 & n6291) | (~Ng4369 & (~Pg35 | n6291));
  assign n4953_1 = ~n8639;
  assign n8641 = n9219 & (\[4437]  | n5967 | ~Ng4581);
  assign n8642 = (Pg35 & n9220) | (~Ng4492 & (~Pg35 | n9220));
  assign n6008 = ~n8642;
  assign n8644 = n9221 & (n5967 | ~Ng4581 | Ng4575);
  assign n8645 = (Pg35 & n9222) | (~Ng4564 & (~Pg35 | n9222));
  assign n1689_1 = ~n8645;
  assign n8647 = n8263 & (n6338 | n8260 | ~Ng2643);
  assign n8648 = n8647 & (~n9106 | (n5999 & ~Ng1589));
  assign n8649 = n8270 & (n6357 | n8267 | ~Ng2509);
  assign n8650 = n8649 & ((n6001 & Ng1589) | ~n9107);
  assign n8651 = n8277 & (n6375 | n8274 | ~Ng2375);
  assign n8652 = n8651 & (~n9108 | (n6011 & ~Ng1589));
  assign n8653 = n8284 & (n6393 | n8281 | ~Ng2241);
  assign n8654 = n8653 & ((n6007 & Ng1589) | ~n9109);
  assign n8655 = n8292 & (n6412 | n8289 | ~Ng2084);
  assign n8656 = n8655 & (~n9110 | (n6003 & ~Ng1246));
  assign n8657 = n8299 & (n6431 | n8296 | ~Ng1950);
  assign n8658 = n8657 & ((n6005 & Ng1246) | ~n9111);
  assign n8659 = n8306 & (n6450 | n8303 | ~Ng1816);
  assign n8660 = n8659 & (~n9112 | (n5997 & ~Ng1246));
  assign n8661 = n8313 & (n6468 | n8310 | ~Ng1682);
  assign n8662 = n8661 & ((n6009 & Ng1246) | ~n9113);
  assign n8663 = (n5967 | Ng269) & (~Pg72 | Ng262);
  assign n8664 = n8663 & (~Pg73 | (~Pg72 & Ng255));
  assign n8665 = (Pg35 & ~n8664) | (~\[4432]  & (~Pg35 | ~n8664));
  assign n1317_1 = ~n8665;
  assign n8667 = Ng239 | Pg73 | ~Pg72;
  assign n8668 = Ng246 | n5967;
  assign n8669 = (Ng232 & (~Pg72 | Ng225)) | (Pg72 & Ng225);
  assign n8670 = n8667 & n8668 & (~Pg73 | n8669);
  assign n8671 = (Pg35 & ~n8670) | (~Ng479 & (~Pg35 | ~n8670));
  assign n2247 = ~n8671;
  assign n8673 = (n5876 & n8321) | (~Ng5644 & (~n5876 | n8321));
  assign n8674 = ~n9225 & (Pg35 | ~Ng5703);
  assign n6086_1 = ~n8674;
  assign n8676 = (Pg35 & ~n8644) | (~Ng4552 & (~Pg35 | ~n8644));
  assign n6413 = ~n8676;
  assign n8678 = (Pg35 & ~n8641) | (~Ng4515 & (~Pg35 | ~n8641));
  assign n6340 = ~n8678;
  assign n8680 = (Ng2667 & Ng2661) | (n8039 & (Ng2667 | ~Ng2661));
  assign n8681 = (~n8262 & ~Ng2661) | (~Ng2667 & (n8262 | ~Ng2661));
  assign n3623 = ~n8681;
  assign n8683 = (~n8262 & ~Ng2643) | (~Ng2648 & (n8262 | ~Ng2643));
  assign n3538 = ~n8683;
  assign n8685 = (n8040 & (~Ng2533 | Ng2527)) | (Ng2533 & Ng2527);
  assign n8686 = (~n8269 & ~Ng2527) | (~Ng2533 & (n8269 | ~Ng2527));
  assign n6022_1 = ~n8686;
  assign n8688 = (~n8269 & ~Ng2509) | (~Ng2514 & (n8269 | ~Ng2509));
  assign n2590_1 = ~n8688;
  assign n8690 = (Ng2399 & Ng2393) | (n8041 & (Ng2399 | ~Ng2393));
  assign n8691 = (~n8276 & ~Ng2393) | (~Ng2399 & (n8276 | ~Ng2393));
  assign n1636_1 = ~n8691;
  assign n8693 = (~n8276 & ~Ng2375) | (~Ng2380 & (n8276 | ~Ng2375));
  assign n3360 = ~n8693;
  assign n8695 = (Ng2265 & Ng2259) | (n8042 & (Ng2265 | ~Ng2259));
  assign n8696 = (~n8283 & ~Ng2259) | (~Ng2265 & (n8283 | ~Ng2259));
  assign n4480 = ~n8696;
  assign n8698 = (~n8283 & ~Ng2241) | (~Ng2246 & (n8283 | ~Ng2241));
  assign n5111 = ~n8698;
  assign n8700 = (n8043 & (~Ng2108 | Ng2102)) | (Ng2108 & Ng2102);
  assign n8701 = (~n8291 & ~Ng2102) | (~Ng2108 & (n8291 | ~Ng2102));
  assign n5261 = ~n8701;
  assign n8703 = (~n8291 & ~Ng2084) | (~Ng2089 & (n8291 | ~Ng2084));
  assign n1026_1 = ~n8703;
  assign n8705 = (n8044 & (~Ng1974 | Ng1968)) | (Ng1974 & Ng1968);
  assign n8706 = (~n8298 & ~Ng1968) | (~Ng1974 & (n8298 | ~Ng1968));
  assign n4509_1 = ~n8706;
  assign n8708 = (~n8298 & ~Ng1950) | (~Ng1955 & (n8298 | ~Ng1950));
  assign n4164 = ~n8708;
  assign n8710 = (Ng1840 & Ng1834) | (n8045 & (Ng1840 | ~Ng1834));
  assign n8711 = (~n8305 & ~Ng1834) | (~Ng1840 & (n8305 | ~Ng1834));
  assign n3411 = ~n8711;
  assign n8713 = (~n8305 & ~Ng1816) | (~Ng1821 & (n8305 | ~Ng1816));
  assign n5366_1 = ~n8713;
  assign n8715 = (Ng1706 & Ng1700) | (n8046 & (Ng1706 | ~Ng1700));
  assign n8716 = (~n8312 & ~Ng1700) | (~Ng1706 & (n8312 | ~Ng1700));
  assign n1616 = ~n8716;
  assign n8718 = (~n8312 & ~Ng1682) | (~Ng1687 & (n8312 | ~Ng1682));
  assign n6012 = ~n8718;
  assign n8720 = n9228 & (~Pg35 | n8245 | ~Ng142);
  assign n1826_1 = ~n8720;
  assign n8722 = (n8354 & (Ng5041 | n8356)) | (~Ng5041 & n8356);
  assign n8723 = (n8353 & (Ng5033 | n8355)) | (~Ng5033 & n8355);
  assign n8724 = ~n9238 & (Ng283 | n7834 | ~Ng287);
  assign n3812_1 = ~n8724;
  assign n8726 = (n7168 & (Pg35 | ~Ng4122)) | (~Pg35 & ~Ng4122);
  assign n1201_1 = ~n8726;
  assign n8728 = (~n7338 & ~Ng2681) | (~Ng2675 & (n7338 | ~Ng2681));
  assign n6017 = ~n8728;
  assign n8730 = (~n7343 & ~Ng2547) | (~Ng2541 & (n7343 | ~Ng2547));
  assign n712 = ~n8730;
  assign n8732 = (~n7348 & ~Ng2413) | (~Ng2407 & (n7348 | ~Ng2413));
  assign n6056 = ~n8732;
  assign n8734 = (~n7353 & ~Ng2279) | (~Ng2273 & (n7353 | ~Ng2279));
  assign n3047 = ~n8734;
  assign n8736 = (~n7358 & ~Ng2122) | (~Ng2116 & (n7358 | ~Ng2122));
  assign n1844_1 = ~n8736;
  assign n8738 = (~n7363 & ~Ng1988) | (~Ng1982 & (n7363 | ~Ng1988));
  assign n6442 = ~n8738;
  assign n8740 = (~n7368 & ~Ng1854) | (~Ng1848 & (n7368 | ~Ng1854));
  assign n4379_1 = ~n8740;
  assign n8742 = (~n7373 & ~Ng1720) | (~Ng1714 & (n7373 | ~Ng1720));
  assign n5850_1 = ~n8742;
  assign n8744 = (n8048 & Ng1413) | (~n8047 & (n8048 | ~Ng1413));
  assign n8745 = n9275 & (~Pg35 | n5559 | n8116);
  assign n5681_1 = ~n8745;
  assign n8747 = (n8050 & Ng1070) | (~n8049 & (n8050 | ~Ng1070));
  assign n8748 = n9276 & (~Pg35 | n4474 | n8118);
  assign n4622 = ~n8748;
  assign n8750 = (~n7407 & ~Ng6519) | (~Ng6513 & (n7407 | ~Ng6519));
  assign n2560_1 = ~n8750;
  assign n8752 = (~n7438 & ~Ng6173) | (~Ng6167 & (n7438 | ~Ng6173));
  assign n4452 = ~n8752;
  assign n8754 = (~n7469 & ~Ng5827) | (~Ng5821 & (n7469 | ~Ng5827));
  assign n3340_1 = ~n8754;
  assign n8756 = (~n7500 & ~Ng5481) | (~Ng5475 & (n7500 | ~Ng5481));
  assign n5806 = ~n8756;
  assign n8758 = (~n7530 & ~Ng5134) | (~Ng5128 & (n7530 | ~Ng5134));
  assign n1327_1 = ~n8758;
  assign n8760 = ~n7559 & n8211 & (n8119 | n8317);
  assign n8761 = ~n7564 & n8209 & (n8120 | n8316);
  assign n8762 = (~n7571 & ~Ng3827) | (~Ng3821 & (n7571 | ~Ng3827));
  assign n3586_1 = ~n8762;
  assign n8764 = (~n7602 & ~Ng3476) | (~Ng3470 & (n7602 | ~Ng3476));
  assign n2178 = ~n8764;
  assign n8766 = (~n7631 & ~Ng3125) | (~Ng3119 & (n7631 | ~Ng3125));
  assign n6395 = ~n8766;
  assign n8768 = ~n9315 & (Pg35 | ~Ng1478);
  assign n1532_1 = ~n8768;
  assign n8770 = ~Ng1489 & ~Ng1442;
  assign n8771 = n8522 & n5170 & (Ng1484 | n8770);
  assign n8772 = ~n9317 & (Pg35 | ~Ng1448);
  assign n2530 = ~n8772;
  assign n8774 = ~n9319 & (Pg35 | ~Ng1442);
  assign n1433_1 = ~n8774;
  assign n8776 = ~n9321 & (Pg35 | ~Ng1135);
  assign n6114_1 = ~n8776;
  assign n8778 = ~Ng1146 & ~Ng1099;
  assign n8779 = n8527 & n4887 & (Ng1141 | n8778);
  assign n8780 = ~n9323 & (Pg35 | ~Ng1105);
  assign n4549 = ~n8780;
  assign n8782 = ~n9325 & (Pg35 | ~Ng1099);
  assign n6502 = ~n8782;
  assign n8784 = n9331 & (~Pg35 | n8360 | n8362);
  assign n5411_1 = ~n8784;
  assign n8786 = n9332 & (~Pg35 | n8361 | n8363);
  assign n5376_1 = ~n8786;
  assign n8788 = n9333 & (~Ng4521 | (Pg35 & n9334));
  assign n4099 = ~n8788;
  assign n8790 = n9335 & (Pg35 | ~Ng2841);
  assign n5753 = ~n8790;
  assign n8792 = (~n7797 & ~Ng4145) | (~Ng4112 & (n7797 | ~Ng4145));
  assign n5481_1 = ~n8792;
  assign n8794 = (~Ng661 & ~n8475) | (~Ng728 & (~Ng661 | n8475));
  assign n6427 = ~n8794;
  assign n8796 = (~Ng718 & ~n8475) | (~Ng661 & (~Ng718 | n8475));
  assign n3106 = ~n8796;
  assign n8798 = (~Ng655 & ~n8475) | (~Ng718 & (~Ng655 | n8475));
  assign n1287_1 = ~n8798;
  assign n8800 = (~Ng650 & ~n8475) | (~Ng655 & (~Ng650 | n8475));
  assign n3439 = ~n8800;
  assign n8802 = (Pg35 & n8124) | (~\[4435]  & (~Pg35 | n8124));
  assign n6531 = ~n8802;
  assign n8804 = (~Ng645 & ~n8475) | (~Ng681 & (~Ng645 | n8475));
  assign n1732_1 = ~n8804;
  assign n8806 = (n7839 & (Pg35 | ~Ng4512)) | (~Pg35 & ~Ng4512);
  assign n1036_1 = ~n8806;
  assign n8808 = (~Pg35 & ~Ng4459) | (~Ng4473 & (Pg35 | ~Ng4459));
  assign n2570 = ~n8808;
  assign n8810 = (Pg35 & n9339) | (~Ng4462 & (~Pg35 | n9339));
  assign n3720_1 = ~n8810;
  assign n8812 = (~Pg35 & ~Ng4558) | (~Pg6749 & (Pg35 | ~Ng4558));
  assign n4075 = ~n8812;
  assign n8814 = (~Pg35 & ~Ng4561) | (~Pg6750 & (Pg35 | ~Ng4561));
  assign n2803_1 = ~n8814;
  assign n8816 = (~Pg35 & ~Ng4555) | (~Pg6748 & (Pg35 | ~Ng4555));
  assign n1224_1 = ~n8816;
  assign n8818 = (~Pg35 & ~Ng4489) | (~Pg6750 & (Pg35 | ~Ng4489));
  assign n1257_1 = ~n8818;
  assign n8820 = (~Pg35 & ~Ng4486) | (~Pg6749 & (Pg35 | ~Ng4486));
  assign n4504 = ~n8820;
  assign n8822 = (~Pg35 & ~Ng4483) | (~Pg6748 & (Pg35 | ~Ng4483));
  assign n2354_1 = ~n8822;
  assign n8824 = (n9241 & (Pg35 | ~Ng4153)) | (~Pg35 & ~Ng4153);
  assign n1925_1 = ~n8824;
  assign n8826 = (Pg35 & n9240) | (~Ng4104 & (~Pg35 | n9240));
  assign n5864 = ~n8826;
  assign n8828 = n9341 & (Pg35 | ~Ng2841);
  assign n4211_1 = ~n8828;
  assign n8830 = (n8128 & (Pg35 | ~Ng1532)) | (~Pg35 & ~Ng1532);
  assign n5558_1 = ~n8830;
  assign n8832 = n9342 & (~Pg35 | n8129 | Ng1322);
  assign n3792 = ~n8832;
  assign n8834 = (n8130 & (Pg35 | ~Ng1189)) | (~Pg35 & ~Ng1189);
  assign n5898 = ~n8834;
  assign n8836 = (Pg35 & n9343) | (~Ng890 & (~Pg35 | n9343));
  assign n3490 = ~n8836;
  assign n8838 = n9344 & (Ng812 | (n8022 & Ng843));
  assign n8839 = (~Ng732 & n9345) | (~Ng753 & (~Ng732 | ~n9345));
  assign n1537_1 = ~n8839;
  assign n8841 = n8468 & ~n9346 & (~Ng528 | n8469);
  assign n8842 = (Pg35 & ~n8841) | (~Ng518 & (~Pg35 | ~n8841));
  assign n2232_1 = ~n8842;
  assign n8844 = Pg35 & (Ng333 | Ng355);
  assign n8845 = (~Ng351 & ~n8844) | (Pg35 & (Ng351 | ~n8844));
  assign n1979_1 = ~n8845;
  assign n8847 = n9347 & (Pg35 | ~Ng347);
  assign n1742_1 = ~n8847;
  assign n8849 = (Ng347 & (Pg35 | ~Ng333)) | (~Pg35 & ~Ng333);
  assign n3558 = ~n8849;
  assign n8851 = n9348 & (Pg35 | ~\[4436] );
  assign n5151_1 = ~n8851;
  assign n8853 = (Pg35 & ~Ng316) | (~\[4431]  & (~Pg35 | ~Ng316));
  assign n3651_1 = ~n8853;
  assign n8855 = (n7912 & (Pg35 | ~Ng336)) | (~Pg35 & ~Ng336);
  assign n6027 = ~n8855;
  assign n8857 = (n7918 & (Pg35 | ~Ng316)) | (~Pg35 & ~Ng316);
  assign n6275 = ~n8857;
  assign n8859 = (~Pg35 & ~Ng305) | (~Pg6744 & (Pg35 | ~Ng305));
  assign n895_1 = ~n8859;
  assign n8861 = (n8381 & ~Ng6505) | (~Ng6541 & (~n8381 | ~Ng6505));
  assign n5136_1 = ~n8861;
  assign n8863 = (Ng6533 & Ng6527) | (n8051 & (Ng6533 | ~Ng6527));
  assign n8864 = (~n8381 & ~Ng6527) | (~Ng6533 & (n8381 | ~Ng6527));
  assign n5541_1 = ~n8864;
  assign n8866 = ~Pg9817 & (Ng6444 | (Pg9743 & ~Ng6494));
  assign n8867 = (~Pg35 & ~Ng6494) | (~n8866 & (Pg35 | ~Ng6494));
  assign n3755_1 = ~n8867;
  assign n8869 = (Pg35 & ~Ng6727) | (~Ng6444 & (~Pg35 | ~Ng6727));
  assign n2306 = ~n8869;
  assign n8871 = (n8386 & ~Ng6159) | (~Ng6195 & (~n8386 | ~Ng6159));
  assign n2007_1 = ~n8871;
  assign n8873 = (Ng6187 & Ng6181) | (n8052 & (Ng6187 | ~Ng6181));
  assign n8874 = (~n8386 & ~Ng6181) | (~Ng6187 & (n8386 | ~Ng6181));
  assign n1893_1 = ~n8874;
  assign n8876 = ~Pg9741 & (Ng6098 | (Pg9682 & ~Ng6148));
  assign n8877 = (~Pg35 & ~Ng6148) | (~n8876 & (Pg35 | ~Ng6148));
  assign n4187 = ~n8877;
  assign n8879 = (Pg35 & ~Ng6381) | (~Ng6098 & (~Pg35 | ~Ng6381));
  assign n1068_1 = ~n8879;
  assign n8881 = (n8390 & ~Ng5813) | (~Ng5849 & (~n8390 | ~Ng5813));
  assign n741_1 = ~n8881;
  assign n8883 = (Ng5841 & Ng5835) | (n8053 & (Ng5841 | ~Ng5835));
  assign n8884 = (~n8390 & ~Ng5835) | (~Ng5841 & (n8390 | ~Ng5835));
  assign n6289 = ~n8884;
  assign n8886 = ~Pg9680 & (Ng5752 | (Pg9617 & ~Ng5802));
  assign n8887 = (~Pg35 & ~Ng5802) | (~n8886 & (Pg35 | ~Ng5802));
  assign n2408_1 = ~n8887;
  assign n8889 = (Pg35 & ~Ng6035) | (~Ng5752 & (~Pg35 | ~Ng6035));
  assign n2328_1 = ~n8889;
  assign n8891 = (n8394 & ~Ng5467) | (~Ng5503 & (~n8394 | ~Ng5467));
  assign n3416 = ~n8891;
  assign n8893 = (Ng5495 & Ng5489) | (n8054 & (Ng5495 | ~Ng5489));
  assign n8894 = (~n8394 & ~Ng5489) | (~Ng5495 & (n8394 | ~Ng5489));
  assign n2379_1 = ~n8894;
  assign n8896 = ~Pg9615 & (Ng5406 | (Pg9555 & ~Ng5456));
  assign n8897 = (~Pg35 & ~Ng5456) | (~n8896 & (Pg35 | ~Ng5456));
  assign n2984_1 = ~n8897;
  assign n8899 = (Pg35 & ~Ng5689) | (~Ng5406 & (~Pg35 | ~Ng5689));
  assign n2848_1 = ~n8899;
  assign n8901 = (~n7934 & ~Ng5120) | (~Ng5156 & (n7934 | ~Ng5120));
  assign n4574 = ~n8901;
  assign n8903 = (Ng5148 & Ng5142) | (n8055 & (Ng5148 | ~Ng5142));
  assign n8904 = (n7934 & ~Ng5142) | (~Ng5148 & (~n7934 | ~Ng5142));
  assign n6565 = ~n8904;
  assign n8906 = ~Pg9497 & (Ng5022 | (Pg9553 & ~Ng5112));
  assign n8907 = (~Pg35 & ~Ng5112) | (~n8906 & (Pg35 | ~Ng5112));
  assign n2285_1 = ~n8907;
  assign n8909 = ~Pg9553 & (Ng5062 | (Pg9497 & ~Ng5109));
  assign n8910 = (~Pg35 & ~Ng5109) | (~n8909 & (Pg35 | ~Ng5109));
  assign n5175_1 = ~n8910;
  assign n8912 = (~Pg35 & ~Ng5062) | (~\[4415]  & (Pg35 | ~Ng5062));
  assign n3009_1 = ~n8912;
  assign n8914 = (Ng5069 & Ng5084) | (Ng5073 & (Ng5069 | ~Ng5084));
  assign n8915 = ~n9351 & (n7566 | ~Ng4057 | Ng4064);
  assign n6250 = ~n8915;
  assign n8917 = (n8401 & ~Ng3813) | (~Ng3849 & (~n8401 | ~Ng3813));
  assign n1072_1 = ~n8917;
  assign n8919 = (Ng3841 & Ng3835) | (n8056 & (Ng3841 | ~Ng3835));
  assign n8920 = (~n8401 & ~Ng3835) | (~Ng3841 & (n8401 | ~Ng3835));
  assign n6507 = ~n8920;
  assign n8922 = ~Pg8398 & (Ng3752 | (Pg8344 & ~Ng3802));
  assign n8923 = (~Pg35 & ~Ng3802) | (~n8922 & (Pg35 | ~Ng3802));
  assign n2743 = ~n8923;
  assign n8925 = (Pg35 & ~Ng4040) | (~Ng3752 & (~Pg35 | ~Ng4040));
  assign n2668_1 = ~n8925;
  assign n8927 = (n8405 & ~Ng3462) | (~Ng3498 & (~n8405 | ~Ng3462));
  assign n5456_1 = ~n8927;
  assign n8929 = (Ng3490 & Ng3484) | (n8057 & (Ng3490 | ~Ng3484));
  assign n8930 = (~n8405 & ~Ng3484) | (~Ng3490 & (n8405 | ~Ng3484));
  assign n815_1 = ~n8930;
  assign n8932 = ~Pg8342 & (Ng3401 | (Pg8279 & ~Ng3451));
  assign n8933 = (~Pg35 & ~Ng3451) | (~n8932 & (Pg35 | ~Ng3451));
  assign n6147 = ~n8933;
  assign n8935 = (Pg35 & ~Ng3689) | (~Ng3401 & (~Pg35 | ~Ng3689));
  assign n6634 = ~n8935;
  assign n8937 = (n8409 & ~Ng3111) | (~Ng3147 & (~n8409 | ~Ng3111));
  assign n1232_1 = ~n8937;
  assign n8939 = (Ng3139 & Ng3133) | (n8058 & (Ng3139 | ~Ng3133));
  assign n8940 = (~n8409 & ~Ng3133) | (~Ng3139 & (n8409 | ~Ng3133));
  assign n2242_1 = ~n8940;
  assign n8942 = ~Pg8277 & (Ng3050 | (Pg8215 & ~Ng3100));
  assign n8943 = (~Pg35 & ~Ng3100) | (~n8942 & (Pg35 | ~Ng3100));
  assign n1831_1 = ~n8943;
  assign n8945 = (Pg35 & ~Ng3338) | (~Ng3050 & (~Pg35 | ~Ng3338));
  assign n5971_1 = ~n8945;
  assign n8947 = n9352 & (~Pg35 | n8134 | n8510);
  assign n6211 = ~n8947;
  assign n8949 = ~n8510 & ((n8133 & Ng1559) | Ng1554);
  assign n8950 = (Pg35 & ~n8949) | (~Ng1559 & (~Pg35 | ~n8949));
  assign n5705_1 = ~n8950;
  assign n8952 = (Pg35 & n9354) | (~Ng1521 & (~Pg35 | n9354));
  assign n5446_1 = ~n8952;
  assign n8954 = n9357 & (~Pg35 | n8136 | n8511);
  assign n2275 = ~n8954;
  assign n8956 = ~n8511 & ((n8135 & Ng1216) | Ng1211);
  assign n8957 = (Pg35 & ~n8956) | (~Ng1216 & (~Pg35 | ~n8956));
  assign n5326_1 = ~n8957;
  assign n8959 = (Pg35 & n9359) | (~Ng1178 & (~Pg35 | n9359));
  assign n2493 = ~n8959;
  assign n8961 = (~n8027 & ~Ng817) | (~n7758 & (~n8027 | Ng817));
  assign n8962 = (n7983 & ~Ng686) | (~Ng667 & (~n7983 | ~Ng686));
  assign n4311_1 = ~n8962;
  assign n8964 = (n8500 & ~Ng452) | (~Ng460 & (~n8500 | ~Ng452));
  assign n726_1 = ~n8964;
  assign n8966 = (~Ng174 & n8500) | (~Ng182 & (~Ng174 | ~n8500));
  assign n1969_1 = ~n8966;
  assign n8968 = (~Ng168 & n8500) | (~Ng174 & (~Ng168 | ~n8500));
  assign n2956_1 = ~n8968;
  assign n8970 = (Pg35 & n9362) | (~Ng358 & (~Pg35 | n9362));
  assign n5568_1 = ~n8970;
  assign n8972 = (Pg35 & n9363) | (~Ng370 & (~Pg35 | n9363));
  assign n5874 = ~n8972;
  assign n8974 = (n9365 & (Pg35 | ~Ng191)) | (~Pg35 & ~Ng191);
  assign n4707_1 = ~n8974;
  assign n8976 = (Pg35 & n9367) | (~Ng222 & (~Pg35 | n9367));
  assign n4138_1 = ~n8976;
  assign n8978 = (Pg35 & Ng218) | (~Ng209 & (~Pg35 | Ng218));
  assign n3267 = ~n8978;
  assign n8980 = n9368 & (~Pg35 | ~n5006 | Ng6736);
  assign n5441_1 = ~n8980;
  assign n8982 = (Pg35 & n9369) | (~Ng6723 & (~Pg35 | n9369));
  assign n1557_1 = ~n8982;
  assign n8984 = n9370 & (~Pg35 | ~n5604 | Ng6390);
  assign n1792 = ~n8984;
  assign n8986 = (Pg35 & n9371) | (~Ng6377 & (~Pg35 | n9371));
  assign n4904 = ~n8986;
  assign n8988 = n9372 & (~Pg35 | ~n5069_1 | Ng6044);
  assign n2999_1 = ~n8988;
  assign n8990 = (Pg35 & n9373) | (~Ng6031 & (~Pg35 | n9373));
  assign n6240 = ~n8990;
  assign n8992 = n9374 & (~Pg35 | ~n5837 | Ng5698);
  assign n5573_1 = ~n8992;
  assign n8994 = (Pg35 & n9375) | (~Ng5685 & (~Pg35 | n9375));
  assign n3215 = ~n8994;
  assign n8996 = n9376 & (~Pg35 | ~n5715 | Ng5352);
  assign n6575 = ~n8996;
  assign n8998 = (Pg35 & n9377) | (~Ng5339 & (~Pg35 | n9377));
  assign n1307_1 = ~n8998;
  assign n9000 = (Pg35 & n9378) | (~Ng4308 & (~Pg35 | n9378));
  assign n2212 = ~n9000;
  assign n9002 = (Pg35 & ~n9383) | (~Ng4235 & (~Pg35 | ~n9383));
  assign n4539 = ~n9002;
  assign n9004 = n9384 & (~Pg35 | ~n4631_1 | Ng4049);
  assign n2525 = ~n9004;
  assign n9006 = (Pg35 & n9385) | (~Ng4031 & (~Pg35 | n9385));
  assign n707_1 = ~n9006;
  assign n9008 = n9386 & (~Pg35 | ~n4267 | Ng3698);
  assign n5801 = ~n9008;
  assign n9010 = (Pg35 & n9387) | (~Ng3680 & (~Pg35 | n9387));
  assign n3476_1 = ~n9010;
  assign n9012 = n9388 & (~Pg35 | ~n5184 | Ng3347);
  assign n1669_1 = ~n9012;
  assign n9014 = (Pg35 & n9389) | (~Ng3329 & (~Pg35 | n9389));
  assign n2979_1 = ~n9014;
  assign n9016 = (Pg35 & ~Ng496) | (~Ng1554 & (~Pg35 | ~Ng496));
  assign n6052_1 = ~n9016;
  assign n9018 = (Pg35 & n9391) | (~Ng1339 & (~Pg35 | n9391));
  assign n944_1 = ~n9018;
  assign n9020 = (Pg35 & n9392) | (~Ng1306 & (~Pg35 | n9392));
  assign n1572_1 = ~n9020;
  assign n9022 = (Pg35 & n9393) | (~Ng1526 & (~Pg35 | n9393));
  assign n6600 = ~n9022;
  assign n9024 = (n7731 & ~Ng1495) | (~Ng1442 & (~n7731 | ~Ng1495));
  assign n1485_1 = ~n9024;
  assign n9026 = (~n7731 & ~Ng1495) | (~Ng1489 & (n7731 | ~Ng1495));
  assign n1428_1 = ~n9026;
  assign n9028 = (~Pg35 & ~Ng1211) | (~\[4432]  & (Pg35 | ~Ng1211));
  assign n2169_1 = ~n9028;
  assign n9030 = (Pg35 & n9395) | (~Ng996 & (~Pg35 | n9395));
  assign n3515 = ~n9030;
  assign n9032 = (Pg35 & n9396) | (~Ng962 & (~Pg35 | n9396));
  assign n1596_1 = ~n9032;
  assign n9034 = (Pg35 & n9397) | (~Ng1183 & (~Pg35 | n9397));
  assign n1277_1 = ~n9034;
  assign n9036 = (n7735 & ~Ng1152) | (~Ng1099 & (~n7735 | ~Ng1152));
  assign n1122_1 = ~n9036;
  assign n9038 = (~n7735 & ~Ng1152) | (~Ng1146 & (n7735 | ~Ng1152));
  assign n5298 = ~n9038;
  assign n9040 = (n7758 & ~Ng854) | (~Ng847 & (~n7758 | ~Ng854));
  assign n785_1 = ~n9040;
  assign n9042 = (~n7758 & ~Ng441) | (~Ng475 & (n7758 | ~Ng441));
  assign n3004_1 = ~n9042;
  assign n9044 = (n7758 & ~Ng441) | (~Ng437 & (~n7758 | ~Ng441));
  assign n1737_1 = ~n9044;
  assign n9046 = (~n7758 & ~Ng429) | (~Ng433 & (n7758 | ~Ng429));
  assign n4777_1 = ~n9046;
  assign n9048 = (n7758 & ~Ng429) | (~Ng401 & (~n7758 | ~Ng429));
  assign n2994_1 = ~n9048;
  assign n9050 = (~n7758 & ~Ng424) | (~Ng411 & (n7758 | ~Ng424));
  assign n5344_1 = ~n9050;
  assign n9052 = (~n7758 & ~Ng405) | (~Ng392 & (n7758 | ~Ng405));
  assign n3223_1 = ~n9052;
  assign n9054 = (Pg35 & n9401) | (~Ng2946 & (~Pg35 | n9401));
  assign n5884 = ~n9054;
  assign n9056 = (Pg35 & n9402) | (~Ng4239 & (~Pg35 | n9402));
  assign n3788_1 = ~n9056;
  assign n9058 = (n8540 & (Pg35 | ~Ng4291)) | (~Pg35 & ~Ng4291);
  assign n4272_1 = ~n9058;
  assign n9060 = (n8541 & (Pg35 | ~Ng4284)) | (~Pg35 & ~Ng4284);
  assign n5007 = ~n9060;
  assign n9062 = (n8542 & (Pg35 | ~Ng4281)) | (~Pg35 & ~Ng4281);
  assign n6512 = ~n9062;
  assign n9064 = (Pg35 & n8543) | (~Ng4245 & (~Pg35 | n8543));
  assign n4160_1 = ~n9064;
  assign n9066 = (Pg35 & Ng4239) | (~Ng4273 & (~Pg35 | Ng4239));
  assign n6522 = ~n9066;
  assign n9068 = (Pg35 & n9379) | (~Ng4180 & (~Pg35 | n9379));
  assign n2384_1 = ~n9068;
  assign n9070 = n6045 | ~Ng2882;
  assign n9071 = ~Ng534 | n8159;
  assign n9072 = (n8153 | ~Ng16) & (n6020 | n8142);
  assign n9073 = n6015 | ~Ng790;
  assign n9074 = ~n5992 & n9073 & (n6027_1 | ~Ng749);
  assign n9075 = (n6063 | ~Ng608) & (n8159 | Ng550);
  assign n9076 = n9075 & (~Ng572 | n8157);
  assign n9077 = (n8153 | ~Ng50) & (n6046 | n8142);
  assign n9078 = (n6045 | ~Ng2886) & (~Ng2980 | n8174);
  assign n9079 = n6063 | ~Ng604;
  assign n9080 = (n8153 | ~Ng51) & (n6032 | n8142);
  assign n9081 = (n8161 | ~Ng1283) & (n8171 | ~Ng2138);
  assign n9082 = n6063 | ~Ng599;
  assign n9083 = ~n5992 & n9082 & (n8157 | ~Ng562);
  assign n9084 = (n6015 | ~Ng781) & (n6027_1 | ~Ng739);
  assign n9085 = n9084 & (n8159 | ~Ng199);
  assign n9086 = (n8153 | ~Ng52) & (n6038 | n8142);
  assign n9087 = (n6045 | ~Ng2848) & (n6056_1 | ~Ng2902);
  assign n9088 = (n6031 | ~Ng2907) & (n6080 | ~Ng2844);
  assign n9089 = (~Ng1300 | n8175) & (~Ng956 | n8176);
  assign n9090 = (Pg35 | n8158) & (n6027_1 | ~Ng772);
  assign n9091 = (n6063 | ~Ng626) & (~Ng590 | n8157);
  assign n9092 = (~Ng1472 | n8175) & (~Ng1129 | n8176);
  assign n9093 = n6015 | ~Ng554;
  assign n9094 = (~Ng1448 | n8175) & (~Ng1105 | n8176);
  assign n9095 = (n8153 | ~Ng8) & (n8171 | ~Ng5507);
  assign n9096 = n6045 | ~Ng2898;
  assign n9097 = n6063 | ~Ng617;
  assign n9098 = (~Ng1478 | n8175) & (~Ng1135 | n8176);
  assign n9099 = (n8153 | ~Ng48) & (n8168 | ~Ng4912);
  assign n9100 = (n8188 | n8189) & (n8190 | n7619);
  assign n9101 = (n5730 | n7578) & (n8191 | n7414);
  assign n9102 = (n7404 | ~n7942) & (n7466 | ~n8218);
  assign n9103 = (n7599 | ~n8220) & (n6261 | n7527);
  assign n9104 = (n7435 | ~n8218) & (n7628 | ~n7942);
  assign n9105 = (n7568 | ~n8220) & (n6261 | n7497);
  assign n9106 = ~n5923 & (n8260 | ~Ng2643);
  assign n9107 = ~n5942 & (n8267 | ~Ng2509);
  assign n9108 = ~n5956_1 & (n8274 | ~Ng2375);
  assign n9109 = ~n5953 & (n8281 | ~Ng2241);
  assign n9110 = ~n5944 & (n8289 | ~Ng2084);
  assign n9111 = ~n5948 & (n8296 | ~Ng1950);
  assign n9112 = ~n5898_1 & (n8303 | ~Ng1816);
  assign n9113 = ~n5954 & (n8310 | ~Ng1682);
  assign n9114 = ~n6268 & n8330;
  assign n9115 = Pg35 & (~n6634_1 | (~Ng1373 & n8333));
  assign n9116 = Pg35 & (~n6641 | (~Ng1030 & n8339));
  assign n9117 = ~n8102 & (n6882 | (~n5880 & ~n8105));
  assign n9118 = (Ng2236 | n8373) & (Ng2370 | n7957);
  assign n9119 = (n7957 | ~Ng2807) & (~Ng2803 | n8373);
  assign n9120 = (Ng1945 | n8370) & (Ng2079 | n8255);
  assign n9121 = (n7957 | ~Ng2775) & (~Ng2771 | n8373);
  assign n9122 = ~Ng6645 | ~Pg17688 | n7423;
  assign n9123 = ~Ng6653 | ~Pg17688 | n7426;
  assign n9124 = ~Ng6283 | ~Pg17760 | n7445;
  assign n9125 = ~Ng6275 | ~Pg14779 | n7457;
  assign n9126 = ~Ng5953 | ~Pg17607 | n7485;
  assign n9127 = ~Ng5961 | ~Pg17607 | n7488;
  assign n9128 = ~Ng5607 | ~Pg17580 | n7516;
  assign n9129 = ~Ng5615 | ~Pg17580 | n7519;
  assign n9130 = ~Ng5260 | ~Pg17519 | n7545;
  assign n9131 = ~Ng5252 | ~Pg17674 | n6516;
  assign n9132 = (~Ng4836 | ~Ng5011) & (~Ng4864 | Ng3333);
  assign n9133 = (~Ng4871 | ~Ng3684) & (~Ng4878 | Ng4035);
  assign n9134 = (~\[4427]  | ~Ng4646) & (~Ng4674 | Ng4821);
  assign n9135 = (~Ng4681 | ~Ng4831) & (~Ng4688 | Ng4826);
  assign n9136 = ~Ng3953 | ~Pg16659 | n7587;
  assign n9137 = ~Ng3945 | ~Pg16775 | n6525;
  assign n9138 = ~Ng3602 | ~Pg16627 | n8455;
  assign n9139 = ~Ng3578 | ~Pg13926 | n8455;
  assign n9140 = ~Ng3235 | ~Pg16718 | n8189;
  assign n9141 = ~Ng3227 | ~Pg13895 | n7649;
  assign n9142 = (n6537 & (n8189 | Ng3347)) | (n8189 & ~Ng3347);
  assign n9143 = (n7638 & (~Ng3343 | n7649)) | (Ng3343 & n7649);
  assign n9144 = ~n8328 & (Ng4939 | (n9142 & n9143));
  assign n9145 = (~Ng5694 & n7519) | (n7516 & (Ng5694 | n7519));
  assign n9146 = (n8321 & Ng5698) | (n7507 & (n8321 | ~Ng5698));
  assign n9147 = ~n8322 & (Ng4749 | (n9145 & n9146));
  assign n9148 = ~Ng979 & (~n7888 | ~Ng1061 | ~Ng1052);
  assign n9149 = Ng832 & (~n7758 | (Pg35 & ~Ng817));
  assign n9150 = (~Pg35 | Pg19357) & (~Ng1395 | n8005);
  assign n9151 = Pg17316 | Pg17400 | Pg17291;
  assign n9152 = (n8014 | ~Ng1052) & (~Pg35 | Pg19334);
  assign n9153 = Pg35 & (n6089 | Ng2984);
  assign n9154 = Ng753 | Ng655 | Ng718;
  assign n9155 = ~Ng4332 & (n5967 | (Pg90 & ~Ng2994));
  assign n9156 = ~Ng4322 & (n9155 | (Ng4332 & Ng4311));
  assign n9157 = ~Ng4332 & Ng4322 & (n5967 | ~Ng4515);
  assign n9158 = Ng4608 | ~Ng4593 | Ng4601 | ~Ng4584;
  assign n9159 = ~Ng4349 & (Ng4340 | n9156 | n9157);
  assign n9160 = ~n9159 & (n5729 | Ng4340 | ~Ng4349);
  assign n9161 = (Ng4340 & ~Ng4349) | (n5729 & (~Ng4340 | ~Ng4349));
  assign n9162 = (n9160 & (~Ng4358 | n9161)) | (Ng4358 & n9161);
  assign n9163 = ~Pg91 | n4212 | n4213 | Ng2965;
  assign n9164 = n9163 & Pg35;
  assign n9165 = n4206_1 | n4207 | n4209 | n4210 | Ng2955 | n8214 | ~n8215 | Ng2946;
  assign n9166 = n9165 & Pg35;
  assign n9167 = Ng2941 | Ng4072 | Ng4153;
  assign n9168 = n9167 & Pg35;
  assign n9169 = Pg35 & ~n9426;
  assign n9170 = Ng2932 | ~Pg44 | Ng2927;
  assign n9171 = n9170 & Pg35;
  assign n9172 = Pg35 & ~n9427;
  assign n9173 = n5969 | Ng301 | Ng2902;
  assign n9174 = n9173 & Pg35;
  assign n9175 = Ng2882 | n4213 | n4212;
  assign n9176 = n9175 & Pg35;
  assign n9177 = Ng2856 | n4209 | n4210;
  assign n9178 = n9177 & Pg35;
  assign n9179 = Ng2848 | n4207 | n4206_1;
  assign n9180 = n9179 & Pg35;
  assign n9181 = n9103 & ~Ng4087 & n9102;
  assign n9182 = n9105 & n9104 & Ng4087;
  assign n9183 = (~Ng2724 & ~Ng2803) | (~Ng2807 & (Ng2724 | ~Ng2803));
  assign n9184 = (~Ng2724 & ~Ng2815) | (~Ng2819 & (Ng2724 | ~Ng2815));
  assign n9185 = (~Ng2724 & ~Ng2771) | (~Ng2775 & (Ng2724 | ~Ng2771));
  assign n9186 = (~Ng2724 & ~Ng2783) | (~Ng2787 & (Ng2724 | ~Ng2783));
  assign n9187 = Pg35 | ~Ng2894;
  assign n9188 = ~Pg35 | ~Ng1291;
  assign n9189 = ~Pg35 | ~Ng947;
  assign n9190 = Ng4878 & (~Pg35 | (~Ng4843 & n8228));
  assign n9191 = Ng4688 & (~Pg35 | (~Ng4653 & n8230));
  assign n9192 = (~n6203 & n6204) | (~Ng4340 & (n6203 | n6204));
  assign n9193 = Pg35 | ~Ng2827;
  assign n9194 = Pg35 | ~Ng2815;
  assign n9195 = Pg35 | ~Ng2819;
  assign n9196 = Pg35 | ~Ng2807;
  assign n9197 = Pg35 | ~Ng2795;
  assign n9198 = Pg35 | ~Ng2783;
  assign n9199 = Pg35 | ~Ng2787;
  assign n9200 = Pg35 | ~Ng2775;
  assign n9201 = (Ng392 & ~Ng452) | (~Ng174 & (~Ng392 | ~Ng452));
  assign n9202 = (~Ng405 & ~Ng424) | (~Ng437 & (Ng405 | ~Ng424));
  assign n9203 = (~Ng405 & ~Ng437) | (~Ng401 & (Ng405 | ~Ng437));
  assign n9204 = (n9202 & (~Ng392 | n9203)) | (Ng392 & n9203);
  assign n9205 = n7768 & n8237;
  assign n9206 = (~Ng4955 & n9205) | (n6274 & (~Ng4955 | ~n9205));
  assign n9207 = n7773 & n8237;
  assign n9208 = (~Ng4944 & n9207) | (n6275_1 & (~Ng4944 | ~n9207));
  assign n9209 = n6125 & n8237;
  assign n9210 = (~Ng4888 & n9209) | (n6280 & (~Ng4888 | ~n9209));
  assign n9211 = n7784 & n8239;
  assign n9212 = (~Ng4765 & n9211) | (n6282 & (~Ng4765 | ~n9211));
  assign n9213 = n7789 & n8239;
  assign n9214 = (~Ng4754 & n9213) | (n6283 & (~Ng4754 | ~n9213));
  assign n9215 = n7796 & n8239;
  assign n9216 = (~Ng4698 & n9215) | (n6288 & (~Ng4698 | ~n9215));
  assign n9217 = Pg35 | ~Ng4340;
  assign n9218 = ~Ng157 | n8250;
  assign n9219 = Ng4512 | Ng4581;
  assign n9220 = (n5967 & ~n8641) | (n8036 & (~n5967 | ~n8641));
  assign n9221 = Ng4552 | Ng4581;
  assign n9222 = (n5967 & ~n8644) | (n8038 & (~n5967 | ~n8644));
  assign n9223 = Pg35 | ~Ng2759;
  assign n9224 = n8320 | ~n5876 | n8188;
  assign n9225 = Pg35 & n9224 & (~n7519 | ~n8673);
  assign n9226 = Pg35 | ~Ng4108;
  assign n9227 = Pg35 | ~Ng2756;
  assign n9228 = Pg35 | ~Ng301;
  assign n9229 = ~Ng5046 | n8354 | ~Ng5041;
  assign n9230 = (n8357 & (~Ng5052 | n9229)) | (Ng5052 & n9229);
  assign n9231 = Pg35 | ~Ng4098;
  assign n9232 = ~Ng5033 & (~n8353 | (Pg35 & ~n8355));
  assign n9233 = ~Ng5052 & (~n9229 | (Pg35 & ~n8357));
  assign n9234 = Pg35 | ~Ng5041;
  assign n9235 = Pg35 | ~Ng5037;
  assign n9236 = Pg35 | ~Ng5033;
  assign n9237 = Pg35 | ~Ng5022;
  assign n9238 = Ng283 & (~Pg35 | (~Ng287 & n8241));
  assign n9239 = ~Ng4473 | Ng4459;
  assign n9240 = (~Pg120 & ~Ng4146) | (~Pg124 & (~Pg120 | Ng4146));
  assign n9241 = (~Pg114 & ~Ng4157) | (~Pg116 & (~Pg114 | Ng4157));
  assign n9242 = (~Ng2504 & ~Ng2715) | (~Ng2638 & (~Ng2504 | Ng2715));
  assign n9243 = (Ng2819 & (Ng2815 | Ng2715)) | (Ng2815 & ~Ng2715);
  assign n9244 = ~n8206 | n5866 | Ng2735;
  assign n9245 = n9244 & (~n9118 | (Ng2719 & n9242));
  assign n9246 = ~n9244 & (~n9119 | (Ng2719 & n9243));
  assign n9247 = (~Ng1677 & ~Ng2715) | (~Ng1811 & (~Ng1677 | Ng2715));
  assign n9248 = (Ng2787 & (Ng2783 | Ng2715)) | (Ng2783 & ~Ng2715);
  assign n9249 = n9244 & (~n9120 | (~Ng2719 & n9247));
  assign n9250 = ~n9244 & (~n9121 | (Ng2719 & n9248));
  assign n9251 = Ng2681 & (~Pg35 | (Ng2675 & n8413));
  assign n9252 = Pg35 & Ng2657 & (~n5920 | n8415);
  assign n9253 = Pg35 & Ng2595 & (~n5920 | n8205);
  assign n9254 = Ng2547 & (~Pg35 | (Ng2541 & n8417));
  assign n9255 = Pg35 & Ng2523 & (~n5919 | n8419);
  assign n9256 = Pg35 & Ng2461 & (~n5919 | n8203);
  assign n9257 = Ng2413 & (~Pg35 | (Ng2407 & n8420));
  assign n9258 = Pg35 & Ng2389 & (~n5925 | n8422);
  assign n9259 = Pg35 & Ng2327 & (~n5925 | n8204);
  assign n9260 = Ng2279 & (~Pg35 | (Ng2273 & n8423));
  assign n9261 = Pg35 & Ng2255 & (~n5878 | n8425);
  assign n9262 = Pg35 & Ng2193 & (~n5878 | n8197);
  assign n9263 = Ng2122 & (~Pg35 | (Ng2116 & n8427));
  assign n9264 = Pg35 & Ng2098 & (~n5916 | n8429);
  assign n9265 = Pg35 & Ng2036 & (~n5916 | n8201);
  assign n9266 = Ng1988 & (~Pg35 | (Ng1982 & n8430));
  assign n9267 = Pg35 & Ng1964 & (~n5899 | n8432);
  assign n9268 = Pg35 & Ng1902 & (~n5899 | n8202);
  assign n9269 = Ng1854 & (~Pg35 | (Ng1848 & n8433));
  assign n9270 = Pg35 & Ng1830 & (~n5941 | n8435);
  assign n9271 = Pg35 & Ng1768 & (~n5941 | n8199);
  assign n9272 = Ng1720 & (~Pg35 | (Ng1714 & n8436));
  assign n9273 = Pg35 & Ng1696 & (~n5868 | n8438);
  assign n9274 = Pg35 & Ng1632 & (~n5868 | n8207);
  assign n9275 = Pg35 | ~Ng1536;
  assign n9276 = Pg35 | ~Ng1193;
  assign n9277 = Ng6519 & (~Pg35 | (~n8440 & Ng6513));
  assign n9278 = Ng6500 & (~Pg35 | (~n8440 & ~Ng6505));
  assign n9279 = ~Pg12470 ^ Ng6727;
  assign n9280 = Pg35 & Ng6500 & (~n5884_1 | n8512);
  assign n9281 = Ng6173 & (~Pg35 | (~n8442 & Ng6167));
  assign n9282 = Ng6154 & (~Pg35 | (~n8442 & ~Ng6159));
  assign n9283 = ~Pg12422 ^ Ng6381;
  assign n9284 = Pg35 & Ng6154 & (~n5952 | ~n8513);
  assign n9285 = Ng5827 & (~Pg35 | (~n8444 & Ng5821));
  assign n9286 = Ng5808 & (~Pg35 | (~n8444 & ~Ng5813));
  assign n9287 = ~Pg12350 ^ Ng6035;
  assign n9288 = Pg35 & Ng5808 & (~n5940 | n8514);
  assign n9289 = Ng5481 & (~Pg35 | (~n8446 & Ng5475));
  assign n9290 = (~Pg35 | (~n8446 & ~Ng5467)) & Ng5462;
  assign n9291 = ~Pg12300 ^ Ng5689;
  assign n9292 = Pg35 & Ng5462 & (~n5876 | n8515);
  assign n9293 = Ng5134 & (~Pg35 | (~n8449 & Ng5128));
  assign n9294 = Ng5115 & (~Pg35 | (~n8449 & ~Ng5120));
  assign n9295 = ~\[4415]  ^ Pg12238;
  assign n9296 = Pg35 & Ng5115 & (~n4151_1 | n8516);
  assign n9297 = ~Ng4983 & (n7555 | Ng4991);
  assign n9298 = n9133 & n9132 & n4483;
  assign n9299 = ~Ng4793 & (n7560 | Ng4801);
  assign n9300 = n9135 & n9134 & n4637;
  assign n9301 = Ng3827 & (~Pg35 | (~n8451 & Ng3821));
  assign n9302 = Ng3808 & (~Pg35 | (~n8451 & ~Ng3813));
  assign n9303 = ~Pg11418 ^ Ng4040;
  assign n9304 = Pg35 & Ng3808 & (~n5927 | n8517);
  assign n9305 = Ng3476 & (~Pg35 | (~n8453 & Ng3470));
  assign n9306 = Ng3457 & (~Pg35 | (~n8453 & ~Ng3462));
  assign n9307 = ~Pg11388 ^ Ng3689;
  assign n9308 = Pg35 & Ng3457 & (~n5889 | n8518);
  assign n9309 = Ng3125 & (~Pg35 | (~n8456 & Ng3119));
  assign n9310 = (~Pg35 | (~n8456 & ~Ng3111)) & Ng3106;
  assign n9311 = ~Pg11349 ^ Ng3338;
  assign n9312 = Pg35 & Ng3106 & (~n5908 | n8519);
  assign n9313 = Pg35 | ~Ng2729;
  assign n9314 = n8521 & n8458 & (Ng1454 | n8770);
  assign n9315 = Pg35 & (n9314 | (~n8458 & Ng1454));
  assign n9316 = n8523 & n8459 & (Ng1467 | n8770);
  assign n9317 = Pg35 & (n9316 | (~n8459 & Ng1467));
  assign n9318 = n8524 & n8460 & (Ng1437 | n8770);
  assign n9319 = Pg35 & (n9318 | (~n8460 & Ng1437));
  assign n9320 = n8526 & n8461 & (Ng1111 | n8778);
  assign n9321 = Pg35 & (n9320 | (~n8461 & Ng1111));
  assign n9322 = n8528 & n8462 & (Ng1124 | n8778);
  assign n9323 = Pg35 & (n9322 | (~n8462 & Ng1124));
  assign n9324 = n8529 & n8463 & (Ng1094 | n8778);
  assign n9325 = Pg35 & (n9324 | (~n8463 & Ng1094));
  assign n9326 = Ng827 & ~n8464;
  assign n9327 = ~Ng676 | ~n8467;
  assign n9328 = Pg35 | ~Ng482;
  assign n9329 = ~Ng417 ^ n9204;
  assign n9330 = Ng417 & (~Pg35 | (~n7976 & n9329));
  assign n9331 = Pg35 | ~Ng5057;
  assign n9332 = Pg35 | ~Ng5069;
  assign n9333 = Ng4521 | ~Pg35 | n5729;
  assign n9334 = ~n8126 ^ Ng4527;
  assign n9335 = ~Ng26936 | ~Pg35 | Ng4125;
  assign n9336 = Pg35 | ~Ng4082;
  assign n9337 = Pg35 | ~Ng1351;
  assign n9338 = Pg35 | ~Ng1008;
  assign n9339 = Ng10384 | Ng4473;
  assign n9340 = n8126 & (~Pg35 | Ng4527);
  assign n9341 = ~Ng26936 | ~Pg35 | Ng2712;
  assign n9342 = Pg35 | ~Ng1395;
  assign n9343 = (~Ng896 & ~Ng862) | (Ng890 & (Ng896 | ~Ng862));
  assign n9344 = ~Ng812 | ~n7758 | n7905;
  assign n9345 = ~Pg35 | n5960;
  assign n9346 = ~Ng528 & (n5933 | n8469);
  assign n9347 = ~Pg35 | ~Pg7540 | Ng347;
  assign n9348 = ~Pg35 | ~Ng329 | ~n8493 | Ng341;
  assign n9349 = ~Pg35 | Ng311 | Ng305 | Ng26885;
  assign n9350 = n7941 & ~Ng5080 & (Ng5069 | ~Ng5077);
  assign n9351 = Ng4064 & (~Pg35 | (~Ng4057 & Ng2841));
  assign n9352 = Pg35 | ~Ng1564;
  assign n9353 = ~Ng1526 | n7379;
  assign n9354 = (~Ng1306 & n9353) | (~Ng1339 & (~Ng1306 | ~n9353));
  assign n9355 = ~n8082 & Ng1389;
  assign n9356 = Ng1351 & (n9355 | n7964);
  assign n9357 = Pg35 | ~Ng1221;
  assign n9358 = ~Ng1183 | n7389;
  assign n9359 = (~Ng962 & n9358) | (~Ng996 & (~Ng962 | ~n9358));
  assign n9360 = ~n8083 & Ng1046;
  assign n9361 = Ng1008 & (n9360 | n7972);
  assign n9362 = ~n6252 ^ Ng370;
  assign n9363 = ~Ng376 ^ Ng358;
  assign n9364 = ~Pg8358 ^ Ng191;
  assign n9365 = (~Ng209 & (~n8501 | n9364)) | (n8501 & n9364);
  assign n9366 = n8501 & n9364;
  assign n9367 = ~Pg8358 ^ n9366;
  assign n9368 = Pg35 | ~Ng6727;
  assign n9369 = ~Ng6727 ^ n8502;
  assign n9370 = Pg35 | ~Ng6381;
  assign n9371 = n8503 ^ Ng6381;
  assign n9372 = Pg35 | ~Ng6035;
  assign n9373 = ~Ng6035 ^ n8504;
  assign n9374 = Pg35 | ~Ng5689;
  assign n9375 = ~Ng5689 ^ n8505;
  assign n9376 = Pg35 | ~\[4415] ;
  assign n9377 = n8506 ^ \[4415] ;
  assign n9378 = ~Pg9251 ^ Ng4308;
  assign n9379 = (Ng4145 & (~Ng4253 | Ng4164)) | (Ng4253 & Ng4164);
  assign n9380 = ~Pg8870 | Ng4235;
  assign n9381 = Pg8918 | Pg8917 | Pg8920 | Pg8919 | Pg11770 | Pg8916 | Pg8915;
  assign n9382 = n9380 & (Pg8870 | (~Ng4235 & n9381));
  assign n9383 = n9382 ^ n9379;
  assign n9384 = Pg35 | ~Ng4040;
  assign n9385 = n8507 ^ Ng4040;
  assign n9386 = Pg35 | ~Ng3689;
  assign n9387 = n8508 ^ Ng3689;
  assign n9388 = Pg35 | ~Ng3338;
  assign n9389 = n8509 ^ Ng3338;
  assign n9390 = Pg13272 | Pg7946 | Pg19357 | Ng1333 | Pg8475;
  assign n9391 = n8007 ^ n9390;
  assign n9392 = (~Pg7946 & ~Ng1532) | (~Ng1521 & (Pg7946 | ~Ng1532));
  assign n9393 = (~Pg7946 & ~Ng1521) | (~Ng1339 & (Pg7946 | ~Ng1521));
  assign n9394 = Pg13259 | Pg7916 | Pg19334 | Ng990 | Pg8416;
  assign n9395 = n8016 ^ n9394;
  assign n9396 = (~Pg7916 & ~Ng1189) | (~Ng1178 & (Pg7916 | ~Ng1189));
  assign n9397 = (~Pg7916 & ~Ng1178) | (~Ng996 & (Pg7916 | ~Ng1178));
  assign n9398 = n8027 | ~Ng822 | ~Ng817 | ~Ng723;
  assign n9399 = ~Pg8786 | Ng4180;
  assign n9400 = Pg8785 | Pg8787 | Pg8783 | Pg8784 | Pg11447 | Pg8788 | Pg8789;
  assign n9401 = n9399 & (Pg8786 | (~Ng4180 & n9400));
  assign n9402 = Ng4297 | Pg10122;
  assign n1335_1 = ~n6714;
  assign n1472_1 = Pg35 & Pg113;
  assign n2083 = ~n6734;
  assign n2136 = ~n6202;
  assign n3336 = ~n6683;
  assign n3524 = ~n6693;
  assign n3847_1 = Pg35 & Pg64;
  assign n4156_1 = ~n6724;
  assign n4331_1 = ~n7967;
  assign n4369 = ~n7975;
  assign n4587_1 = ~n7852;
  assign n5686 = ~n7997;
  assign n6226 = ~n6664;
  assign n1242_1 = Pg35 & Pg125;
  assign n9417 = Ng4125 | n6263 | Ng4057 | Ng4064;
  assign n9418 = n5947 | n9181 | n9182;
  assign n9419 = n8319 | n5730 | ~n5927;
  assign n9420 = n8319 | ~n5884_1 | n8191;
  assign n9421 = n8320 | n5730 | ~n5952;
  assign n9422 = n8320 | ~n4151_1 | n8191;
  assign n9423 = n8320 | ~n5940 | n8190;
  assign n9424 = n8319 | ~n5889 | n8190;
  assign n9425 = n8319 | ~n5908 | n8188;
  assign n9426 = n4218 & n4219 & ~Ng2975;
  assign n9427 = ~n8478 & n4217 & ~Ng2917;
  assign n9428 = n8329 & n8067 & n5911 & ~n6273;
  assign n9429 = n8329 & n8069 & n5872 & ~n6269;
  assign n9430 = n8329 & n8071 & n5910 & ~n6270_1;
  assign n9431 = n8329 & n8073 & n5873 & ~n6271;
  assign n9432 = n8329 & n8075 & n5921 & ~n6267;
  assign n9433 = n8329 & n8077 & n5887 & ~n6272;
  assign n9434 = n8329 & n8079 & n5894 & ~n6266;
  assign n9435 = n8329 & n8081 & n4162 & ~n6268;
  assign n9436 = n7979 & n5983 & n7978 & n5984;
  assign n9437 = ~Ng1389 & n7879 & ~n8484;
  assign n9438 = ~Ng1046 & n7890 & ~n8489;
  assign n9439 = n8229 & ~n6193 & Ng4849;
  assign n9440 = n8231 & ~n6198 & Ng4659;
  assign n9441 = Ng608 & n6259 & ~n8183;
  assign n9442 = Ng604 & n6297_1 & ~n8183;
  assign n9443 = n6361 & Ng2449 & Pg35;
  assign n9444 = n6379 & Ng2315 & Pg35;
  assign n9445 = n6454 & Ng1756 & Pg35;
  assign n9446 = Ng599 & n6490 & ~n8183;
  assign n9447 = Ng595 & n6649 & ~n8183;
  assign n9448 = Ng590 & n6839 & ~n8183;
  assign n9449 = n6654 & Ng6597 & Pg35;
  assign n9450 = n6900 & Ng6653 & Pg35;
  assign n9451 = n6914 & Ng6633 & Pg35;
  assign n9452 = n6970 & Ng6287 & Pg35;
  assign n9453 = n6972 & Ng6283 & Pg35;
  assign n9454 = n6977 & Ng6275 & Pg35;
  assign n9455 = n6673 & Ng5905 & Pg35;
  assign n9456 = n7008 & Ng5961 & Pg35;
  assign n9457 = n7022 & Ng5941 & Pg35;
  assign n9458 = n6682 & Ng5559 & Pg35;
  assign n9459 = n7077 & Ng5595 & Pg35;
  assign n9460 = n7124 & Ng5260 & Pg35;
  assign n9461 = n7129 & Ng5252 & Pg35;
  assign n9462 = n7131 & Ng5248 & Pg35;
  assign n9463 = n7187 & Ng3953 & Pg35;
  assign n9464 = n7192 & Ng3945 & Pg35;
  assign n9465 = n7194 & Ng3941 & Pg35;
  assign n9466 = n7241 & Ng3602 & Pg35;
  assign n9467 = n7249 & Ng3590 & Pg35;
  assign n9468 = n7257 & Ng3578 & Pg35;
  assign n9469 = n7304 & Ng3239 & Pg35;
  assign n9470 = n7306 & Ng3235 & Pg35;
  assign n9471 = n7311 & Ng3227 & Pg35;
  assign n9472 = ~Pg35 & Ng1454;
  assign n9473 = ~Pg35 & Ng1111;
  assign n9474 = n7936 & \[4434]  & Pg35;
  assign n1457 = ~n6802;
  assign n5056_1 = ~n6812;
  assign n6335 = ~n6822;
  assign n4736_1 = ~n8002;
  assign n6137 = ~n6709;
  assign n1517 = ~n6752;
  assign n4020 = ~n6762;
  assign n1993_1 = ~n6772;
  assign n4412_1 = ~n6782;
  assign n5893_1 = ~n6792;
  assign n4422 = ~n7947;
  assign n4432_1 = ~n7959;
  assign n6359 = ~n6705;
  assign n6570 = ~n7163;
  assign Pg34956 = n4124_1;
  assign Pg34839 = n4124_1;
  assign Pg34788 = n4133;
  assign Pg34437 = n4135;
  assign Pg34436 = n4136;
  assign Pg33959 = n4151_1;
  assign Pg33894 = n4133;
  assign Pg33533 = n4162;
  assign Pg31861 = \[4415] ;
  assign Pg31665 = n4135;
  assign Pg31656 = n4136;
  assign Pg30332 = \[4421] ;
  assign Pg29221 = \[4426] ;
  assign Pg29220 = \[4427] ;
  assign Pg29219 = \[4428] ;
  assign Pg29218 = \[4507] ;
  assign Pg29217 = \[4430] ;
  assign Pg29216 = \[4431] ;
  assign Pg29215 = \[4432] ;
  assign Pg29214 = \[4433] ;
  assign Pg29213 = \[4434] ;
  assign Pg29212 = \[4435] ;
  assign Pg29211 = \[4436] ;
  assign Pg29210 = \[4437] ;
  assign Pg28753 = n4151_1;
  assign Pg27831 = n4162;
  assign Pg25219 = \[4415] ;
  assign Pg24185 = Pg44;
  assign Pg24184 = Pg135;
  assign Pg24183 = Pg134;
  assign Pg24182 = Pg127;
  assign Pg24181 = Pg126;
  assign Pg24180 = Pg125;
  assign Pg24179 = Pg124;
  assign Pg24178 = Pg120;
  assign Pg24177 = Pg116;
  assign Pg24176 = Pg115;
  assign Pg24175 = Pg114;
  assign Pg24174 = Pg113;
  assign Pg24173 = Pg100;
  assign Pg24172 = Pg99;
  assign Pg24171 = Pg92;
  assign Pg24170 = Pg91;
  assign Pg24169 = Pg90;
  assign Pg24168 = Pg84;
  assign Pg24167 = Pg73;
  assign Pg24166 = Pg72;
  assign Pg24165 = Pg64;
  assign Pg24164 = Pg57;
  assign Pg24163 = Pg56;
  assign Pg24162 = Pg54;
  assign Pg24161 = Pg53;
  assign Pg23683 = \[4421] ;
  assign Pg21698 = Pg36;
  assign Pg21292 = \[4426] ;
  assign Pg21270 = \[4430] ;
  assign Pg21245 = \[4427] ;
  assign Pg21176 = \[4431] ;
  assign Pg20901 = \[4432] ;
  assign Pg20899 = \[4435] ;
  assign Pg20763 = \[4436] ;
  assign Pg20654 = \[4428] ;
  assign Pg20652 = \[4433] ;
  assign Pg20557 = \[4434] ;
  assign Pg20049 = \[4437] ;
  assign Pg18881 = \[4507] ;
  assign Pg18101 = Pg6746;
  assign Pg18100 = Pg6751;
  assign Pg18099 = Pg6745;
  assign Pg18098 = Pg6744;
  assign Pg18097 = Pg6747;
  assign Pg18096 = Pg6750;
  assign Pg18095 = Pg6749;
  assign Pg18094 = Pg6748;
  assign Pg18092 = Pg6753;
  assign Pg8403 = \[4651] ;
  assign Pg8353 = \[4651] ;
  assign Pg8283 = \[4658] ;
  assign Pg8235 = \[4658] ;
  assign Pg8178 = \[4661] ;
  assign Pg8132 = \[4661] ;
  assign n716 = Pg9048;
  assign n780_1 = Pg17715;
  assign n823_1 = Pg8920;
  assign n837_1 = Pg16656;
  assign n851_1 = Ng4571;
  assign n914_1 = Pg17743;
  assign n1022_1 = Pg16874;
  assign n1045_1 = Pg16627;
  assign n1136_1 = Pg17580;
  assign n1174 = Pg12368;
  assign n1177 = Pg17739;
  assign n1205_1 = Pg14694;
  assign n1228_1 = Pg17649;
  assign n1331_1 = Pg17320;
  assign n1358_1 = Pg14217;
  assign n1411_1 = Pg17722;
  assign n1423 = Pg8215;
  assign n1442 = Pg10527;
  assign n1481 = Pg16775;
  assign n1495_1 = Ng26960;
  assign n1513 = Pg12422;
  assign n1650 = Pg16744;
  assign n1717_1 = Pg9617;
  assign n1816_1 = Pg11678;
  assign n1840 = Pg17711;
  assign n1912_1 = Pg14673;
  assign n1920_1 = Pg17639;
  assign n1959 = Pg16722;
  assign n1983_1 = Pg17400;
  assign n2002_1 = Pg8344;
  assign n2031 = Pg13966;
  assign n2074 = Pg17760;
  assign n2096_1 = Pg8839;
  assign n2120_1 = Pg10122;
  assign n2124 = Pg12350;
  assign n2127_1 = Pg19357;
  assign n2150 = Pg7946;
  assign n2261_1 = Pg14597;
  assign n2289_1 = Pg14518;
  assign n2297_1 = Pg16924;
  assign n2309_1 = Pg17423;
  assign n2313 = Pg7245;
  assign n2331_1 = Pg9682;
  assign n2345_1 = Pg14125;
  assign n2432 = Pg11418;
  assign n2445 = Pg14096;
  assign n2458 = Pg8475;
  assign n2502 = Pg8870;
  assign n2619_1 = Ng26936;
  assign n2663 = Pg9497;
  assign n2701_1 = Pg11388;
  assign n2729_1 = Pg14779;
  assign n2752_1 = Pg11447;
  assign n2755_1 = Pg12923;
  assign n2774_1 = Pg8915;
  assign n2876_1 = Pg9251;
  assign n2885_1 = Pg8416;
  assign n2934_1 = Ng6974;
  assign n2937_1 = Pg11349;
  assign n2941_1 = Ng26959;
  assign n2975_1 = Pg17787;
  assign n3061 = Pg14189;
  assign n3079 = Pg8784;
  assign n3082 = Pg17519;
  assign n3219_1 = Pg19334;
  assign n3232_1 = Pg9743;
  assign n3270 = Pg7257;
  assign n3279_1 = Ng10384;
  assign n3282_1 = Pg17577;
  assign n3379 = Pg16693;
  assign n3382_1 = Pg17291;
  assign n3435_1 = Pg12238;
  assign n3468_1 = Pg16955;
  assign n3471 = Pg10306;
  assign n3480_1 = Pg17678;
  assign n3561 = Pg7260;
  assign n3595 = Pg13049;
  assign n3608_1 = Pg13259;
  assign n3627 = Pg8788;
  assign n3779 = Pg17607;
  assign n3900_1 = Pg14147;
  assign n3903_1 = Pg13039;
  assign n3971_1 = Pg14749;
  assign n3984_1 = Pg14635;
  assign n3992 = Pg16659;
  assign n4010_1 = Pg10500;
  assign n4039_1 = Pg14738;
  assign n4042 = Pg8719;
  assign n4066 = Pg12470;
  assign n4084 = Pg8279;
  assign n4151 = Pg12919;
  assign n4178_1 = Pg17871;
  assign n4206 = Pg8358;
  assign n4235_1 = Pg13068;
  assign n4263_1 = Pg14421;
  assign n4340_1 = Pg14451;
  assign n4393_1 = Pg8917;
  assign n4456 = Pg14705;
  assign n4489 = Pg17845;
  assign n4492_1 = Pg17674;
  assign n4495 = Pg8783;
  assign n4578 = Pg14662;
  assign n4640_1 = Pg13926;
  assign n4648 = Pg8918;
  assign n4731_1 = \[4507] ;
  assign n4770_1 = Pg13085;
  assign n4773_1 = Pg13099;
  assign n4846_1 = Pg13272;
  assign n4851_1 = Ng6972;
  assign n4855_1 = Pg8916;
  assign n4868_1 = Pg16748;
  assign n4877 = \[4661] ;
  assign n4890 = Pg7243;
  assign n4894_1 = Pg14167;
  assign n4948_1 = Pg7540;
  assign n4987 = Pg17764;
  assign n5060 = Pg13895;
  assign n5083_1 = Pg9019;
  assign n5107 = Pg8787;
  assign n5160_1 = Pg8291;
  assign n5237_1 = Pg12184;
  assign n5265_1 = Pg17646;
  assign n5269_1 = Ng25;
  assign n5322 = Pg17819;
  assign n5335_1 = Pg14201;
  assign n5353_1 = Pg17404;
  assign n5356_1 = Pg33435;
  assign n5385_1 = \[4658] ;
  assign n5389_1 = Pg17685;
  assign n5402_1 = Pg17316;
  assign n5521_1 = Ng26885;
  assign n5545_1 = Pg16624;
  assign n5662 = Pg17688;
  assign n5690 = \[4651] ;
  assign n5714 = Pg14828;
  assign n5776 = Ng4520;
  assign n5825_1 = Pg13906;
  assign n5828_1 = Pg33079;
  assign n5842_1 = Pg8785;
  assign n5859 = Pg9553;
  assign n5937 = Pg17778;
  assign n5994_1 = Pg17813;
  assign n6100_1 = Pg11770;
  assign n6123_1 = Pg16718;
  assign n6156 = Pg13881;
  assign n6169 = Pg16686;
  assign n6192 = Pg7916;
  assign n6293 = Pg12300;
  assign n6306_1 = Pg8919;
  assign n6373 = Pg17604;
  assign n6376 = Pg16603;
  assign n6399 = Pg13865;
  assign n6526 = Pg8789;
  assign n6555 = Pg9555;
  assign n6642 = Pg8786;
  always @ (posedge clk) begin
    Ng5057 <= n687;
    Ng2771 <= n692_1;
    Ng1882 <= n697_1;
    Ng2299 <= n702_1;
    Ng4040 <= n707_1;
    Ng2547 <= n712;
    Ng559 <= n716;
    Ng3243 <= n721_1;
    Ng452 <= n726_1;
    Ng3542 <= n731_1;
    Ng5232 <= n736_1;
    Ng5813 <= n741_1;
    Ng2907 <= n746_1;
    Ng1744 <= n751_1;
    Ng5909 <= n756_1;
    Ng1802 <= n761_1;
    Ng3554 <= n766_1;
    Ng6219 <= n771_1;
    Ng807 <= n776_1;
    Ng6031 <= n780_1;
    Ng847 <= n785_1;
    Ng976 <= n790_1;
    Ng4172 <= n795_1;
    Ng4372 <= n800_1;
    Ng3512 <= n805_1;
    Ng749 <= n810_1;
    Ng3490 <= n815_1;
    Pg12350 <= n820_1;
    Ng4235 <= n823_1;
    Ng1600 <= n828_1;
    Ng1714 <= n833_1;
    Pg14451 <= n837_1;
    Ng3155 <= n841_1;
    Ng2236 <= n846_1;
    Ng4555 <= n851_1;
    Ng3698 <= n856_1;
    Ng1736 <= n861_1;
    Ng1968 <= n866_1;
    Ng4621 <= n871_1;
    Ng5607 <= n876_1;
    Ng2657 <= n881_1;
    Pg12300 <= n886_1;
    Ng490 <= n890_1;
    Ng311 <= n895_1;
    Ng772 <= n900_1;
    Ng5587 <= n905_1;
    Ng6177 <= n910_1;
    Ng6377 <= n914_1;
    Ng3167 <= n919_1;
    Ng5615 <= n924_1;
    Ng4567 <= n929;
    Ng3457 <= n934_1;
    Ng6287 <= n939_1;
    Pg7946 <= n944_1;
    Ng2563 <= n948_1;
    Ng4776 <= n953_1;
    Ng4593 <= n958_1;
    Ng6199 <= n963_1;
    Ng2295 <= n968_1;
    Ng1384 <= n973_1;
    Ng1339 <= n978_1;
    Ng5180 <= n983_1;
    Ng2844 <= n988_1;
    Ng1024 <= n993_1;
    Ng5591 <= n998_1;
    Ng3598 <= n1003_1;
    Ng4264 <= n1008_1;
    Ng767 <= n1013_1;
    Ng5853 <= n1018_1;
    Pg13865 <= n1022_1;
    Ng2089 <= n1026_1;
    Ng4933 <= n1031_1;
    Ng4521 <= n1036_1;
    Ng5507 <= n1041_1;
    Pg16656 <= n1045_1;
    Ng6291 <= n1049_1;
    Ng294 <= n1054_1;
    Ng5559 <= n1059_1;
    Pg9617 <= n1064_1;
    Pg9741 <= n1068_1;
    Ng3813 <= n1072_1;
    Ng562 <= n1077_1;
    Ng608 <= n1082;
    Ng1205 <= n1087_1;
    Ng3909 <= n1092_1;
    Ng6259 <= n1097_1;
    Ng5905 <= n1102;
    Ng921 <= n1107_1;
    Ng2955 <= n1112_1;
    Ng203 <= n1117;
    Ng1099 <= n1122_1;
    Ng4878 <= n1127;
    Ng5204 <= n1132_1;
    Pg17604 <= n1136_1;
    Ng3606 <= n1140_1;
    Ng1926 <= n1145_1;
    Ng6215 <= n1150_1;
    Ng3586 <= n1155_1;
    Ng291 <= n1160_1;
    Ng4674 <= n1165_1;
    Ng3570 <= n1170_1;
    Pg9048 <= n1174;
    Pg17607 <= n1177;
    Ng1862 <= n1181;
    Ng676 <= n1186;
    Ng843 <= n1191_1;
    Ng4332 <= n1196_1;
    Ng4153 <= n1201_1;
    Pg17711 <= n1205_1;
    Ng6336 <= n1209_1;
    Ng622 <= n1214;
    Ng3506 <= n1219_1;
    Ng4558 <= n1224_1;
    Pg17685 <= n1228_1;
    Ng3111 <= n1232_1;
    \[4430]  <= n1237_1;
    Ng26936 <= n1242_1;
    Ng939 <= n1247;
    Ng278 <= n1252;
    Ng4492 <= n1257_1;
    Ng4864 <= n1262;
    Ng1036 <= n1267_1;
    \[4427]  <= n1272_1;
    Ng1178 <= n1277_1;
    Ng3239 <= n1282_1;
    Ng718 <= n1287_1;
    Ng6195 <= n1292_1;
    Ng1135 <= n1297_1;
    Ng6395 <= n1302;
    \[4415]  <= n1307_1;
    Ng554 <= n1312_1;
    Ng496 <= n1317_1;
    Ng3853 <= n1322_1;
    Ng5134 <= n1327_1;
    Pg17404 <= n1331_1;
    Pg8344 <= n1335_1;
    Ng2485 <= n1339_1;
    Ng925 <= n1344;
    Ng48 <= n1349_1;
    Ng5555 <= n1354_1;
    Pg14096 <= n1358_1;
    Ng1798 <= n1362_1;
    Ng4076 <= n1367;
    Ng2941 <= n1372_1;
    Ng3905 <= n1377_1;
    Ng763 <= n1382_1;
    Ng6255 <= n1387_1;
    Ng4375 <= n1392_1;
    Ng4871 <= n1397_1;
    Ng4722 <= n1402_1;
    Ng590 <= n1407_1;
    Pg13099 <= n1411_1;
    Ng1632 <= n1415_1;
    Pg12238 <= n1420;
    Ng3100 <= n1423;
    Ng1495 <= n1428_1;
    Ng1437 <= n1433_1;
    Ng6154 <= n1438_1;
    Ng1579 <= n1442;
    Ng5567 <= n1447;
    Ng1752 <= n1452_1;
    Ng1917 <= n1457;
    Ng744 <= n1462_1;
    Ng4737 <= n1467;
    \[4661]  <= n1472_1;
    Ng6267 <= n1477;
    Pg16659 <= n1481;
    Ng1442 <= n1485_1;
    Ng5965 <= n1490;
    Ng4477 <= n1495_1;
    Pg10500 <= n1500;
    Ng4643 <= n1504;
    Ng5264 <= n1509;
    Pg14779 <= n1513;
    Ng2610 <= n1517;
    Ng5160 <= n1522_1;
    Ng5933 <= n1527;
    Ng1454 <= n1532_1;
    Ng753 <= n1537_1;
    Ng1296 <= n1542_1;
    Ng3151 <= n1547_1;
    Ng2980 <= n1552_1;
    Ng6727 <= n1557_1;
    Ng3530 <= n1562_1;
    Ng4104 <= n1567;
    Ng1532 <= n1572_1;
    Pg9251 <= n1577_1;
    Ng2177 <= n1581;
    Ng52 <= n1586;
    Ng4754 <= n1591_1;
    Ng1189 <= n1596_1;
    Ng2287 <= n1601_1;
    Ng4273 <= n1606_1;
    Ng1389 <= n1611_1;
    Ng1706 <= n1616;
    Ng5835 <= n1621_1;
    Ng1171 <= n1626_1;
    Ng4269 <= n1631_1;
    Ng2399 <= n1636_1;
    Ng4983 <= n1641_1;
    Ng5611 <= n1646_1;
    Pg16627 <= n1650;
    Ng4572 <= n1654;
    Ng3143 <= n1659;
    Ng2898 <= n1664_1;
    Ng3343 <= n1669_1;
    Ng3235 <= n1674;
    Ng4543 <= n1679_1;
    Ng3566 <= n1684_1;
    Ng4534 <= n1689_1;
    Ng4961 <= n1694_1;
    Ng4927 <= n1699_1;
    Ng2259 <= n1704_1;
    Ng2819 <= n1709_1;
    Pg7257 <= n1714;
    Ng5802 <= n1717_1;
    Ng2852 <= n1722_1;
    Ng417 <= n1727_1;
    Ng681 <= n1732_1;
    Ng437 <= n1737_1;
    Ng351 <= n1742_1;
    Ng5901 <= n1747_1;
    Ng2886 <= n1752;
    Ng3494 <= n1757_1;
    Ng5511 <= n1762_1;
    Ng3518 <= n1767_1;
    Ng1604 <= n1772;
    Ng5092 <= n1777;
    Ng4831 <= n1782_1;
    Ng4382 <= n1787_1;
    Ng6386 <= n1792;
    Ng479 <= n1797;
    Ng3965 <= n1802;
    Ng4749 <= n1807_1;
    Ng2008 <= n1812_1;
    Ng736 <= n1816_1;
    Ng3933 <= n1821_1;
    Ng222 <= n1826_1;
    Ng3050 <= n1831_1;
    Ng1052 <= n1836_1;
    Pg17580 <= n1840;
    Ng2122 <= n1844_1;
    Ng2465 <= n1849_1;
    Ng5889 <= n1854;
    Ng4495 <= n1859_1;
    Pg8719 <= n1864_1;
    Ng4653 <= n1868;
    Ng3179 <= n1873_1;
    Ng1728 <= n1878_1;
    Ng2433 <= n1883_1;
    Ng3835 <= n1888_1;
    Ng6187 <= n1893_1;
    Ng4917 <= n1898_1;
    Ng1070 <= n1903_1;
    Ng822 <= n1908_1;
    Pg17715 <= n1912_1;
    Ng914 <= n1916_1;
    Ng5339 <= n1920_1;
    Ng4164 <= n1925_1;
    Ng969 <= n1930_1;
    Ng2807 <= n1935_1;
    Ng4054 <= n1940_1;
    Ng6191 <= n1945_1;
    Ng5077 <= n1950_1;
    Ng5523 <= n1955;
    Ng3680 <= n1959;
    Ng6637 <= n1964;
    Ng174 <= n1969_1;
    Ng1682 <= n1974_1;
    Ng355 <= n1979_1;
    Ng1087 <= n1983_1;
    Ng1105 <= n1988;
    Ng2342 <= n1993_1;
    Ng6307 <= n1998_1;
    Ng3802 <= n2002_1;
    Ng6159 <= n2007_1;
    Ng2255 <= n2012_1;
    Ng2815 <= n2017_1;
    Ng911 <= n2022_1;
    Ng43 <= n2027_1;
    Pg16775 <= n2031;
    Ng1748 <= n2035;
    Ng5551 <= n2040;
    Ng3558 <= n2045;
    Ng5499 <= n2050;
    Ng2960 <= n2055_1;
    Ng3901 <= n2060;
    Ng4888 <= n2065_1;
    Ng6251 <= n2070;
    Pg17649 <= n2074;
    Ng1373 <= n2078_1;
    Pg8215 <= n2083;
    Ng157 <= n2087;
    Ng2783 <= n2092;
    Ng4281 <= n2096_1;
    Ng3574 <= n2101_1;
    Ng2112 <= n2106_1;
    Ng1283 <= n2111;
    Ng433 <= n2116;
    Ng4297 <= n2120_1;
    Pg14738 <= n2124;
    Pg13272 <= n2127_1;
    Ng758 <= n2131_1;
    Ng4639 <= n2136;
    Ng6537 <= n2141_1;
    Ng5543 <= n2146;
    Pg8475 <= n2150;
    Ng5961 <= n2154;
    Ng6243 <= n2159_1;
    Ng632 <= n2164_1;
    Pg12919 <= n2169_1;
    Ng3889 <= n2173_1;
    Ng3476 <= n2178;
    Ng1664 <= n2183_1;
    Ng1246 <= n2188_1;
    Ng6629 <= n2193;
    Ng246 <= n2198;
    Ng4049 <= n2203_1;
    Pg7260 <= n2208_1;
    Ng2932 <= n2212;
    Ng4575 <= n2217_1;
    Ng4098 <= n2222;
    Ng4498 <= n2227;
    Ng528 <= n2232_1;
    Ng16 <= n2237_1;
    Ng3139 <= n2242_1;
    \[4432]  <= n2247;
    Ng4584 <= n2252;
    Ng142 <= n2257;
    Pg17639 <= n2261_1;
    Ng5831 <= n2265;
    Ng239 <= n2270_1;
    Ng1216 <= n2275;
    Ng2848 <= n2280_1;
    Ng5022 <= n2285_1;
    Pg16955 <= n2289_1;
    Ng1030 <= n2293_1;
    Pg13881 <= n2297_1;
    Ng3231 <= n2301_1;
    Pg9817 <= n2306;
    Ng1430 <= n2309_1;
    Ng4452 <= n2313;
    Ng2241 <= n2318_1;
    Ng1564 <= n2323_1;
    Pg9680 <= n2328_1;
    Ng6148 <= n2331_1;
    Ng6649 <= n2336_1;
    Ng110 <= n2341_1;
    Pg14147 <= n2345_1;
    Ng225 <= n2349_1;
    Ng4486 <= n2354_1;
    Ng4504 <= n2359_1;
    Ng5873 <= n2364_1;
    Ng5037 <= n2369_1;
    Ng2319 <= n2374_1;
    Ng5495 <= n2379_1;
    Pg11770 <= n2384_1;
    Ng5208 <= n2388_1;
    Ng5579 <= n2393_1;
    Ng5869 <= n2398_1;
    Ng1589 <= n2403_1;
    Ng5752 <= n2408_1;
    Ng6279 <= n2413;
    Ng5917 <= n2418;
    Ng2975 <= n2423;
    Ng6167 <= n2428_1;
    Pg13966 <= n2432;
    Ng2599 <= n2436_1;
    Ng1448 <= n2441_1;
    Pg14125 <= n2445;
    Ng2370 <= n2449_1;
    Ng5164 <= n2454_1;
    Ng1333 <= n2458;
    Ng153 <= n2463_1;
    Ng6549 <= n2468_1;
    Ng4087 <= n2473_1;
    Ng4801 <= n2478_1;
    Ng2984 <= n2483;
    Ng3961 <= n2488_1;
    Ng962 <= n2493;
    Ng101 <= n2498_1;
    Pg8918 <= n2502;
    Ng6625 <= n2506;
    Ng51 <= n2511_1;
    Ng1018 <= n2516;
    Pg17320 <= n2521_1;
    Ng4045 <= n2525;
    Ng1467 <= n2530;
    Ng2461 <= n2535_1;
    Ng2756 <= n2540;
    Ng5990 <= n2545_1;
    Ng1256 <= n2550_1;
    Ng5029 <= n2555_1;
    Ng6519 <= n2560_1;
    Ng1816 <= n2565_1;
    Ng4369 <= n2570;
    Ng4578 <= n2575;
    Ng4459 <= n2580_1;
    Ng3831 <= n2585_1;
    Ng2514 <= n2590_1;
    Ng3288 <= n2595_1;
    Ng2403 <= n2600_1;
    Ng2145 <= n2605_1;
    Ng1700 <= n2610_1;
    Ng513 <= n2615_1;
    Ng2841 <= n2619_1;
    Ng5297 <= n2624_1;
    Ng2763 <= n2629_1;
    Ng4793 <= n2634_1;
    Ng952 <= n2639_1;
    Ng1263 <= n2644_1;
    Ng1950 <= n2649_1;
    Ng5138 <= n2654;
    Ng2307 <= n2659_1;
    Ng5109 <= n2663;
    Pg8398 <= n2668_1;
    Ng4664 <= n2672_1;
    Ng2223 <= n2677_1;
    Ng5808 <= n2682_1;
    Ng6645 <= n2687_1;
    Ng2016 <= n2692_1;
    Ng3873 <= n2697;
    Pg13926 <= n2701_1;
    Ng2315 <= n2705_1;
    Ng2811 <= n2710_1;
    Ng5957 <= n2715_1;
    Ng2047 <= n2720_1;
    Ng3869 <= n2725_1;
    Pg17760 <= n2729_1;
    Ng5575 <= n2733_1;
    Ng46 <= n2738_1;
    Ng3752 <= n2743;
    Ng3917 <= n2748_1;
    Pg8783 <= n2752_1;
    Ng1585 <= n2755_1;
    Ng4388 <= n2760_1;
    Ng6275 <= n2765_1;
    Ng6311 <= n2770;
    Pg8916 <= n2774_1;
    Ng1041 <= n2778_1;
    Ng2595 <= n2783_1;
    Ng2537 <= n2788_1;
    \[4426]  <= n2793_1;
    Ng4430 <= n2798_1;
    Ng4564 <= n2803_1;
    Ng4826 <= n2808_1;
    Ng6239 <= n2813_1;
    Ng232 <= n2818_1;
    Ng5268 <= n2823_1;
    Ng6545 <= n2828;
    Ng2417 <= n2833_1;
    Ng1772 <= n2838_1;
    Ng5052 <= n2843_1;
    Pg9615 <= n2848_1;
    Ng1890 <= n2852_1;
    Ng2629 <= n2857_1;
    Ng572 <= n2862_1;
    Ng2130 <= n2867_1;
    Ng4108 <= n2872_1;
    Ng4308 <= n2876_1;
    Ng475 <= n2881_1;
    Ng990 <= n2885_1;
    Ng45 <= n2890_1;
    Pg12184 <= n2895_1;
    Ng3990 <= n2899_1;
    Ng5881 <= n2904_1;
    Ng1992 <= n2909_1;
    Ng3171 <= n2914_1;
    Ng812 <= n2919_1;
    Ng832 <= n2924_1;
    Ng5897 <= n2929_1;
    Ng4571 <= n2934_1;
    Pg13895 <= n2937_1;
    Ng4455 <= n2941_1;
    Ng2902 <= n2946_1;
    Ng333 <= n2951_1;
    Ng168 <= n2956_1;
    Ng2823 <= n2961_1;
    Ng3684 <= n2966_1;
    Ng3639 <= n2971_1;
    Pg14597 <= n2975_1;
    Ng3338 <= n2979_1;
    Ng5406 <= n2984_1;
    Ng269 <= n2989_1;
    Ng401 <= n2994_1;
    Ng6040 <= n2999_1;
    Ng441 <= n3004_1;
    Pg9553 <= n3009_1;
    Ng3808 <= n3013_1;
    Ng10384 <= n3018_1;
    Ng3957 <= n3023_1;
    Ng4093 <= n3028_1;
    Ng1760 <= n3033_1;
    Pg12422 <= n3038_1;
    Ng160 <= n3042_1;
    Ng2279 <= n3047;
    Ng3498 <= n3052;
    Ng586 <= n3057;
    Pg14201 <= n3061;
    Ng2619 <= n3065_1;
    Ng1183 <= n3070;
    Ng1608 <= n3075;
    Pg8785 <= n3079;
    Pg17577 <= n3082;
    Ng1779 <= n3086_1;
    Ng2652 <= n3091;
    Ng2193 <= n3096_1;
    Ng2393 <= n3101_1;
    Ng661 <= n3106;
    Ng4950 <= n3111;
    Ng5535 <= n3116_1;
    Ng2834 <= n3121;
    Ng1361 <= n3126;
    Ng6235 <= n3131_1;
    Ng1146 <= n3136;
    Ng2625 <= n3141_1;
    Ng150 <= n3146;
    Ng1696 <= n3151_1;
    Ng6555 <= n3156_1;
    Pg14189 <= n3161;
    Ng3881 <= n3165;
    Ng6621 <= n3170_1;
    Ng3470 <= n3175_1;
    Ng3897 <= n3180_1;
    Ng518 <= n3185_1;
    Ng538 <= n3190;
    Ng2606 <= n3195;
    Ng1472 <= n3200;
    Ng542 <= n3205;
    Ng5188 <= n3210_1;
    Ng5689 <= n3215;
    Pg13259 <= n3219_1;
    Ng405 <= n3223_1;
    Ng5216 <= n3228;
    Ng6494 <= n3232_1;
    Ng4669 <= n3237;
    Ng996 <= n3242_1;
    Ng4531 <= n3247_1;
    Ng2860 <= n3252;
    Ng4743 <= n3257_1;
    Ng6593 <= n3262_1;
    Pg8291 <= n3267;
    Ng4411 <= n3270;
    Ng1413 <= n3275_1;
    Ng26960 <= n3279_1;
    Pg13039 <= n3282_1;
    Ng6641 <= n3286_1;
    Ng1936 <= n3291_1;
    Ng55 <= n3296_1;
    Ng504 <= n3301;
    Ng2587 <= n3306_1;
    Ng4480 <= n3311;
    Ng2311 <= n3316_1;
    Ng3602 <= n3321;
    Ng5571 <= n3326_1;
    Ng3578 <= n3331_1;
    Pg9555 <= n3336;
    Ng5827 <= n3340_1;
    Ng3582 <= n3345;
    Ng6271 <= n3350_1;
    Ng4688 <= n3355_1;
    Ng2380 <= n3360;
    Ng5196 <= n3365_1;
    Ng3227 <= n3370_1;
    Ng2020 <= n3375;
    Pg14518 <= n3379;
    Pg17316 <= n3382_1;
    Ng6541 <= n3386_1;
    Ng3203 <= n3391_1;
    Ng1668 <= n3396_1;
    Ng4760 <= n3401_1;
    Ng262 <= n3406_1;
    Ng1840 <= n3411;
    Ng5467 <= n3416;
    Ng460 <= n3421_1;
    Ng6209 <= n3426_1;
    \[4436]  <= n3431_1;
    Pg14662 <= n3435_1;
    Ng655 <= n3439;
    Ng3502 <= n3444_1;
    Ng2204 <= n3449;
    Ng5256 <= n3454;
    Ng4608 <= n3459_1;
    Ng794 <= n3464_1;
    Pg13906 <= n3468_1;
    Ng4423 <= n3471;
    Ng3689 <= n3476_1;
    Ng5685 <= n3480_1;
    Ng703 <= n3485_1;
    Ng862 <= n3490;
    Ng3247 <= n3495_1;
    Ng2040 <= n3500_1;
    Ng4146 <= n3505;
    Ng4633 <= n3510_1;
    Pg7916 <= n3515;
    Ng4732 <= n3519_1;
    Pg9497 <= n3524;
    Ng5817 <= n3528_1;
    Ng2351 <= n3533;
    Ng2648 <= n3538;
    Ng6736 <= n3543;
    Ng4944 <= n3548;
    Ng4072 <= n3553;
    Pg7540 <= n3558;
    Ng4443 <= n3561;
    Ng3466 <= n3566_1;
    Ng4116 <= n3571_1;
    Ng5041 <= n3576;
    Ng4434 <= n3581_1;
    Ng3827 <= n3586_1;
    Ng6500 <= n3591_1;
    Pg17813 <= n3595;
    Ng3133 <= n3599;
    Ng3333 <= n3604;
    Ng979 <= n3608_1;
    Ng4681 <= n3613_1;
    Ng298 <= n3618_1;
    Ng2667 <= n3623;
    Pg8789 <= n3627;
    Ng1894 <= n3631;
    Ng2988 <= n3636_1;
    Ng3538 <= n3641;
    Ng301 <= n3646_1;
    Ng341 <= n3651_1;
    Ng827 <= n3656_1;
    Pg17291 <= n3661;
    Ng2555 <= n3665_1;
    Ng5011 <= n3670_1;
    Ng199 <= n3675;
    Ng6523 <= n3680_1;
    Ng1526 <= n3685_1;
    Ng4601 <= n3690_1;
    Ng854 <= n3695;
    Ng1484 <= n3700;
    Ng4922 <= n3705;
    Ng5080 <= n3710_1;
    Ng5863 <= n3715_1;
    Ng4581 <= n3720_1;
    Ng2518 <= n3725;
    Ng2567 <= n3730;
    Ng568 <= n3735;
    Ng3263 <= n3740;
    Ng6613 <= n3745;
    Ng6044 <= n3750_1;
    Ng6444 <= n3755_1;
    Ng2965 <= n3760;
    Ng5857 <= n3765_1;
    Ng1616 <= n3770_1;
    Ng890 <= n3775;
    Pg17646 <= n3779;
    Ng3562 <= n3783_1;
    Pg10122 <= n3788_1;
    Ng1404 <= n3792;
    Ng3817 <= n3797_1;
    Ng93 <= n3802_1;
    Ng4501 <= n3807_1;
    Ng287 <= n3812_1;
    Ng2724 <= n3817_1;
    Ng4704 <= n3822_1;
    Ng22 <= n3827_1;
    Ng2878 <= n3832_1;
    Ng5220 <= n3837_1;
    Ng617 <= n3842_1;
    Pg12368 <= n3847_1;
    Ng316 <= n3851_1;
    Ng1277 <= n3856;
    Ng6513 <= n3861_1;
    Ng336 <= n3866_1;
    Ng2882 <= n3871_1;
    Ng933 <= n3876_1;
    Ng1906 <= n3881_1;
    Ng305 <= n3886;
    Ng8 <= n3891_1;
    Ng2799 <= n3896;
    Pg14167 <= n3900_1;
    Pg17787 <= n3903_1;
    Ng4912 <= n3907_1;
    Ng4157 <= n3912;
    Ng2541 <= n3917;
    Ng2153 <= n3922;
    Ng550 <= n3927;
    Ng255 <= n3932;
    Ng1945 <= n3937_1;
    Ng5240 <= n3942_1;
    Ng1478 <= n3947;
    Ng3863 <= n3952_1;
    Ng1959 <= n3957_1;
    Ng3480 <= n3962;
    Ng6653 <= n3967_1;
    Pg17764 <= n3971_1;
    Ng2864 <= n3975;
    Ng4894 <= n3980_1;
    Pg17678 <= n3984_1;
    Ng3857 <= n3988;
    Pg16693 <= n3992;
    Ng499 <= n3996_1;
    Ng1002 <= n4001;
    Ng776 <= n4006;
    Ng1236 <= n4010_1;
    Ng4646 <= n4015;
    Ng2476 <= n4020;
    Ng1657 <= n4025_1;
    Ng2375 <= n4030;
    Ng63 <= n4035_1;
    Pg17739 <= n4039_1;
    Ng358 <= n4042;
    Ng896 <= n4047_1;
    Ng283 <= n4052_1;
    Ng3161 <= n4057;
    Ng2384 <= n4062;
    Pg14828 <= n4066;
    Ng4616 <= n4070_1;
    Ng4561 <= n4075;
    Ng2024 <= n4080;
    Ng3451 <= n4084;
    Ng2795 <= n4089_1;
    Ng613 <= n4094_1;
    Ng4527 <= n4099;
    Ng1844 <= n4104;
    Ng5937 <= n4109;
    Ng4546 <= n4114_1;
    Ng2523 <= n4119;
    Pg11349 <= n4124;
    Ng2643 <= n4128;
    Ng1489 <= n4133_1;
    Pg8358 <= n4138_1;
    Ng2551 <= n4142_1;
    Ng5156 <= n4147;
    \[4421]  <= n4151;
    Pg8279 <= n4156_1;
    Pg8839 <= n4160_1;
    Ng1955 <= n4164;
    Ng6049 <= n4169_1;
    Ng2273 <= n4174;
    Pg14749 <= n4178_1;
    Ng4771 <= n4182_1;
    Ng6098 <= n4187;
    Ng3147 <= n4192_1;
    Ng3347 <= n4197;
    Ng2269 <= n4202_1;
    Ng191 <= n4206;
    Ng2712 <= n4211_1;
    Ng626 <= n4216;
    Ng2729 <= n4221_1;
    Ng5357 <= n4226_1;
    Ng4991 <= n4231_1;
    Pg17819 <= n4235_1;
    Ng4709 <= n4239_1;
    Ng2927 <= n4244;
    Ng4340 <= n4249;
    Ng5929 <= n4254;
    Ng4907 <= n4259_1;
    Pg16874 <= n4263_1;
    Ng4035 <= n4267_1;
    Ng2946 <= n4272_1;
    Ng918 <= n4277_1;
    Ng4082 <= n4282;
    Pg9743 <= n4287_1;
    Ng2036 <= n4291_1;
    Ng577 <= n4296_1;
    Ng1620 <= n4301_1;
    Ng2831 <= n4306;
    Ng667 <= n4311_1;
    Ng930 <= n4316_1;
    Ng3937 <= n4321_1;
    Ng817 <= n4326_1;
    Ng1249 <= n4331_1;
    Ng837 <= n4336_1;
    Pg16924 <= n4340_1;
    Ng599 <= n4344_1;
    Ng5475 <= n4349_1;
    Ng739 <= n4354_1;
    Ng5949 <= n4359_1;
    Ng6682 <= n4364_1;
    Ng904 <= n4369;
    Ng2873 <= n4374_1;
    Ng1854 <= n4379_1;
    Ng5084 <= n4384_1;
    Ng5603 <= n4389_1;
    Pg8870 <= n4393_1;
    Ng2495 <= n4397_1;
    Ng2437 <= n4402_1;
    Ng2102 <= n4407_1;
    Ng2208 <= n4412_1;
    Ng2579 <= n4417_1;
    Ng4064 <= n4422;
    Ng4899 <= n4427_1;
    Ng2719 <= n4432_1;
    Ng4785 <= n4437;
    Ng5583 <= n4442_1;
    Ng781 <= n4447;
    Ng6173 <= n4452;
    Pg17743 <= n4456;
    Ng2917 <= n4460;
    Ng686 <= n4465_1;
    Ng1252 <= n4470;
    Ng671 <= n4475;
    Ng2265 <= n4480;
    Ng6283 <= n4485;
    Pg14705 <= n4489;
    Pg17519 <= n4492_1;
    Pg8784 <= n4495;
    Ng5527 <= n4499;
    Ng4489 <= n4504;
    Ng1974 <= n4509_1;
    Ng1270 <= n4514;
    Ng4966 <= n4519;
    Ng6227 <= n4524;
    Ng3929 <= n4529;
    Ng5503 <= n4534;
    Ng4242 <= n4539;
    Ng5925 <= n4544_1;
    Ng1124 <= n4549;
    Ng4955 <= n4554;
    Ng5224 <= n4559_1;
    Ng2012 <= n4564_1;
    Ng6203 <= n4569_1;
    Ng5120 <= n4574;
    Pg17674 <= n4578;
    Ng2389 <= n4582_1;
    Ng4438 <= n4587_1;
    Ng2429 <= n4592;
    Ng2787 <= n4597_1;
    Ng1287 <= n4602;
    Ng2675 <= n4607;
    \[4507]  <= n4612;
    Ng4836 <= n4617;
    Ng1199 <= n4622;
    Pg19357 <= n4627;
    Ng5547 <= n4631;
    Ng2138 <= n4636;
    Pg16744 <= n4640_1;
    Ng2338 <= n4644;
    Pg8919 <= n4648;
    Ng6247 <= n4652_1;
    Ng2791 <= n4657_1;
    Ng3949 <= n4662;
    Ng1291 <= n4667_1;
    Ng5945 <= n4672_1;
    Ng5244 <= n4677_1;
    Ng2759 <= n4682;
    Ng6741 <= n4687;
    Ng785 <= n4692_1;
    Ng1259 <= n4697_1;
    Ng3484 <= n4702_1;
    Ng209 <= n4707_1;
    Ng6609 <= n4712_1;
    Ng5517 <= n4717_1;
    Ng2449 <= n4722_1;
    Ng2575 <= n4727_1;
    Ng65 <= n4731_1;
    Ng2715 <= n4736_1;
    Ng936 <= n4741_1;
    Ng2098 <= n4746;
    Ng4462 <= n4751_1;
    Ng604 <= n4756;
    Ng6589 <= n4761_1;
    Ng1886 <= n4766;
    Pg17845 <= n4770_1;
    Pg17871 <= n4773_1;
    Ng429 <= n4777_1;
    Ng1870 <= n4782;
    Ng4249 <= n4787_1;
    Ng1825 <= n4792_1;
    Ng1008 <= n4797;
    Ng4392 <= n4802;
    Ng3546 <= n4807_1;
    Ng5236 <= n4812;
    Ng1768 <= n4817;
    Ng4854 <= n4822;
    Ng3925 <= n4827;
    Ng6509 <= n4832_1;
    Ng732 <= n4837_1;
    Ng2504 <= n4842_1;
    Ng1322 <= n4846_1;
    Ng4520 <= n4851_1;
    Pg8917 <= n4855_1;
    Ng2185 <= n4859_1;
    Ng37 <= n4864_1;
    Ng4031 <= n4868_1;
    Ng2070 <= n4873_1;
    \[4658]  <= n4877;
    Ng4176 <= n4882;
    Pg11418 <= n4887_1;
    Ng4405 <= n4890;
    Ng872 <= n4894_1;
    Ng6181 <= n4899;
    Ng6381 <= n4904;
    Ng4765 <= n4909_1;
    Ng5563 <= n4914_1;
    Ng1395 <= n4919_1;
    Ng1913 <= n4924_1;
    Ng2331 <= n4929_1;
    Ng6263 <= n4934_1;
    Ng50 <= n4939;
    Ng3945 <= n4944;
    Ng347 <= n4948_1;
    Ng4473 <= n4953_1;
    Ng1266 <= n4958_1;
    Ng5489 <= n4963_1;
    Ng714 <= n4968_1;
    Ng2748 <= n4973;
    Ng5471 <= n4978;
    Ng4540 <= n4983_1;
    Ng6723 <= n4987;
    Ng6605 <= n4992;
    Ng2445 <= n4997;
    Ng2173 <= n5002;
    Pg9019 <= n5007;
    Ng2491 <= n5011_1;
    Ng4849 <= n5016;
    Ng2169 <= n5021;
    Ng2283 <= n5026;
    Ng6585 <= n5031_1;
    \[4428]  <= n5036;
    Ng2407 <= n5041;
    Ng2868 <= n5046_1;
    Ng2767 <= n5051_1;
    Ng1783 <= n5056_1;
    Pg16718 <= n5060;
    Ng1312 <= n5064;
    Ng5212 <= n5069;
    Ng4245 <= n5074_1;
    Ng645 <= n5079_1;
    Ng4291 <= n5083_1;
    \[4435]  <= n5088_1;
    Ng182 <= n5093_1;
    Ng1129 <= n5098;
    Ng2227 <= n5103;
    Pg8788 <= n5107;
    Ng2246 <= n5111;
    Ng1830 <= n5116;
    Ng3590 <= n5121;
    Ng392 <= n5126;
    Ng1592 <= n5131;
    Ng6505 <= n5136_1;
    Ng1221 <= n5141;
    Ng5921 <= n5146;
    \[4431]  <= n5151_1;
    Ng146 <= n5156;
    Ng218 <= n5160_1;
    Ng1932 <= n5165_1;
    Ng1624 <= n5170_1;
    Ng5062 <= n5175_1;
    Ng5462 <= n5180_1;
    Ng2689 <= n5185_1;
    Ng6573 <= n5190_1;
    Ng1677 <= n5195_1;
    Ng2028 <= n5200_1;
    Ng2671 <= n5205_1;
    Pg10527 <= n5210_1;
    Pg7243 <= n5214_1;
    Ng1848 <= n5218_1;
    \[4434]  <= n5223_1;
    Ng5485 <= n5228_1;
    Ng2741 <= n5233_1;
    Pg11678 <= n5237_1;
    Ng2638 <= n5241_1;
    Ng4122 <= n5246_1;
    Ng4322 <= n5251;
    Ng5941 <= n5256_1;
    Ng2108 <= n5261;
    Pg13068 <= n5265_1;
    Ng25 <= n5269_1;
    Ng1644 <= n5273;
    Ng595 <= n5278_1;
    Ng2217 <= n5283_1;
    Ng1319 <= n5288_1;
    Ng2066 <= n5293_1;
    Ng1152 <= n5298;
    Ng5252 <= n5303_1;
    Ng2165 <= n5308_1;
    Ng2571 <= n5313_1;
    Ng5176 <= n5318;
    Pg14673 <= n5322;
    Ng1211 <= n5326_1;
    Ng2827 <= n5331_1;
    Pg14217 <= n5335_1;
    Ng4859 <= n5339_1;
    Ng424 <= n5344_1;
    Ng1274 <= n5349;
    Pg17423 <= n5353_1;
    Ng85 <= n5356_1;
    Ng2803 <= n5361_1;
    Ng1821 <= n5366_1;
    Ng2509 <= n5371_1;
    Ng5073 <= n5376_1;
    Ng1280 <= n5381_1;
    \[4651]  <= n5385_1;
    Pg13085 <= n5389_1;
    Ng6633 <= n5393_1;
    Ng5124 <= n5398_1;
    Pg17400 <= n5402_1;
    Ng6303 <= n5406_1;
    Ng5069 <= n5411_1;
    Ng2994 <= n5416;
    Ng650 <= n5421_1;
    Ng1636 <= n5426_1;
    Ng3921 <= n5431_1;
    Ng2093 <= n5436;
    Ng6732 <= n5441_1;
    Ng1306 <= n5446_1;
    Ng1061 <= n5451_1;
    Ng3462 <= n5456_1;
    Ng2181 <= n5461;
    Ng956 <= n5466_1;
    Ng1756 <= n5471_1;
    Ng5849 <= n5476_1;
    Ng4112 <= n5481_1;
    Ng2685 <= n5486_1;
    Ng2197 <= n5491_1;
    Ng2421 <= n5496_1;
    Ng1046 <= n5501_1;
    Ng482 <= n5506_1;
    Ng4401 <= n5511_1;
    Ng1514 <= n5516_1;
    Ng329 <= n5521_1;
    Ng6565 <= n5526_1;
    Ng2950 <= n5531_1;
    Ng1345 <= n5536_1;
    Ng6533 <= n5541_1;
    Pg14421 <= n5545_1;
    Ng4727 <= n5549_1;
    Pg12470 <= n5554_1;
    Ng1536 <= n5558_1;
    Ng3941 <= n5563_1;
    Ng370 <= n5568_1;
    Ng5694 <= n5573_1;
    Ng1858 <= n5578_1;
    Ng446 <= n5583_1;
    Ng3219 <= n5588_1;
    Ng1811 <= n5593_1;
    Ng6601 <= n5598;
    Ng2441 <= n5603_1;
    Ng1874 <= n5608_1;
    Ng4349 <= n5613_1;
    Ng6581 <= n5618_1;
    Ng6597 <= n5623_1;
    Ng3610 <= n5628;
    Ng2890 <= n5633;
    Ng1978 <= n5638;
    Ng1612 <= n5643_1;
    Ng112 <= n5648_1;
    Ng2856 <= n5653;
    Ng1982 <= n5658_1;
    Pg17722 <= n5662;
    Ng5228 <= n5666_1;
    Ng4119 <= n5671;
    Ng6390 <= n5676_1;
    Ng1542 <= n5681_1;
    Ng4258 <= n5686;
    Ng4818 <= n5690;
    Ng5033 <= n5695;
    Ng4717 <= n5700_1;
    Ng1554 <= n5705_1;
    Ng3849 <= n5710_1;
    Pg17778 <= n5714;
    Ng3199 <= n5718;
    Ng5845 <= n5723_1;
    Ng4975 <= n5728;
    Ng790 <= n5733_1;
    Ng5913 <= n5738_1;
    Ng1902 <= n5743_1;
    Ng6163 <= n5748;
    Ng4125 <= n5753;
    Ng4821 <= n5758_1;
    Ng4939 <= n5763;
    Pg19334 <= n5768;
    Ng3207 <= n5772;
    Ng4483 <= n5776;
    Ng3259 <= n5781_1;
    Ng5142 <= n5786;
    Ng5248 <= n5791;
    Ng2126 <= n5796;
    Ng3694 <= n5801;
    Ng5481 <= n5806;
    Ng1964 <= n5811;
    Ng5097 <= n5816_1;
    Ng3215 <= n5821_1;
    Pg16748 <= n5825_1;
    Ng111 <= n5828_1;
    Ng4427 <= n5833_1;
    Ng2779 <= n5838_1;
    Pg8786 <= n5842_1;
    Pg7245 <= n5846;
    Ng1720 <= n5850_1;
    Ng1367 <= n5855_1;
    Ng5112 <= n5859;
    Ng4145 <= n5864;
    Ng2161 <= n5869;
    Ng376 <= n5874;
    Ng2361 <= n5879_1;
    Pg11447 <= n5884;
    Ng582 <= n5888_1;
    Ng2051 <= n5893_1;
    Ng1193 <= n5898;
    Ng2327 <= n5903_1;
    Ng907 <= n5908_1;
    Ng947 <= n5913_1;
    Ng1834 <= n5918_1;
    Ng3594 <= n5923_1;
    Ng2999 <= n5928_1;
    Ng2303 <= n5933_1;
    Pg17688 <= n5937;
    Ng699 <= n5941_1;
    Ng723 <= n5946_1;
    Ng5703 <= n5951_1;
    Ng546 <= n5956;
    Ng2472 <= n5961_1;
    Ng5953 <= n5966_1;
    Pg8277 <= n5971_1;
    Ng1740 <= n5975_1;
    Ng3550 <= n5980_1;
    Ng3845 <= n5985_1;
    Ng2116 <= n5990;
    Pg14635 <= n5994_1;
    Ng3195 <= n5998;
    Ng3913 <= n6003_1;
    Pg10306 <= n6008;
    Ng1687 <= n6012;
    Ng2681 <= n6017;
    Ng2533 <= n6022_1;
    Ng324 <= n6027;
    Ng2697 <= n6032_1;
    Ng4417 <= n6037_1;
    Ng6561 <= n6042;
    Ng1141 <= n6047_1;
    Pg12923 <= n6052_1;
    Ng2413 <= n6056;
    Ng1710 <= n6061;
    Ng6527 <= n6066_1;
    Ng3255 <= n6071_1;
    Ng1691 <= n6076_1;
    Ng2936 <= n6081;
    Ng5644 <= n6086_1;
    Ng5152 <= n6091;
    Ng5352 <= n6096;
    Pg8915 <= n6100_1;
    Ng2775 <= n6104;
    Ng2922 <= n6109_1;
    Ng1111 <= n6114_1;
    Ng5893 <= n6119_1;
    Pg16603 <= n6123_1;
    Ng6617 <= n6127;
    Ng2060 <= n6132_1;
    Ng4512 <= n6137;
    Ng5599 <= n6142;
    Ng3401 <= n6147;
    Ng4366 <= n6152;
    Pg16722 <= n6156;
    \[4433]  <= n6160;
    Ng3129 <= n6165;
    Ng3329 <= n6169;
    Ng5170 <= n6174_1;
    Ng26959 <= n6179;
    Ng5821 <= n6183;
    Ng6299 <= n6188_1;
    Pg8416 <= n6192;
    Ng2079 <= n6196;
    Ng4698 <= n6201_1;
    Ng3703 <= n6206;
    Ng1559 <= n6211;
    Ng943 <= n6216;
    Ng411 <= n6221;
    Pg9682 <= n6226;
    Ng3953 <= n6230;
    Ng2704 <= n6235;
    Ng6035 <= n6240;
    Ng1300 <= n6245;
    Ng4057 <= n6250;
    Ng5200 <= n6255;
    Ng4843 <= n6260;
    Ng5046 <= n6265;
    Ng2250 <= n6270;
    Ng26885 <= n6275;
    Ng4549 <= n6279;
    Ng2453 <= n6284;
    Ng5841 <= n6289;
    Pg14694 <= n6293;
    Ng2912 <= n6297;
    Ng2357 <= n6302;
    Pg8920 <= n6306_1;
    Ng164 <= n6310;
    Ng4253 <= n6315;
    Ng5016 <= n6320;
    Ng3119 <= n6325_1;
    Ng1351 <= n6330;
    Ng1648 <= n6335;
    Ng6972 <= n6340;
    Ng5115 <= n6344_1;
    Ng3352 <= n6349;
    Ng6657 <= n6354;
    Ng4552 <= n6359;
    Ng3893 <= n6364_1;
    Ng3211 <= n6369;
    Pg13049 <= n6373;
    Pg16624 <= n6376;
    Ng5595 <= n6380;
    Ng3614 <= n6385;
    Ng2894 <= n6390;
    Ng3125 <= n6395;
    Pg16686 <= n6399;
    Ng3821 <= n6403;
    Ng4141 <= n6408_1;
    Ng6974 <= n6413;
    Ng5272 <= n6417;
    Ng2735 <= n6422;
    Ng728 <= n6427;
    Ng6295 <= n6432;
    Ng2661 <= n6437;
    Ng1988 <= n6442;
    Ng5128 <= n6447;
    Ng1548 <= n6452;
    Ng3106 <= n6457;
    Ng4659 <= n6462;
    Ng4358 <= n6467;
    Ng1792 <= n6472;
    Ng2084 <= n6477;
    Ng3187 <= n6482;
    Ng4311 <= n6487;
    Ng2583 <= n6492;
    Ng3003 <= n6497;
    Ng1094 <= n6502;
    Ng3841 <= n6507;
    Ng4284 <= n6512;
    Ng3191 <= n6517;
    Ng4239 <= n6522;
    Ng4180 <= n6526;
    Ng691 <= n6531;
    Ng534 <= n6536;
    Ng385 <= n6541;
    Ng2004 <= n6546;
    Ng2527 <= n6551;
    Ng5456 <= n6555;
    Ng4420 <= n6560;
    Ng5148 <= n6565;
    Ng4507 <= n6570;
    Ng5348 <= n6575;
    Ng3223 <= n6580;
    Ng2970 <= n6585;
    Ng5698 <= n6590;
    Ng5260 <= n6595;
    Ng1521 <= n6600;
    Ng3522 <= n6605;
    Ng3115 <= n6610;
    Ng3251 <= n6615;
    Pg12832 <= n6620;
    Ng4628 <= n6624;
    Ng1996 <= n6629;
    Pg8342 <= n6634;
    Ng4515 <= n6638;
    Pg8787 <= n6642;
    Ng4300 <= n6646;
    Ng1724 <= n6651;
    Ng1379 <= n6656;
    Pg11388 <= n6661;
    Ng1878 <= n6665;
    Ng5619 <= n6670;
    Ng71 <= n6675;
    \[4437]  <= n6680;
  end
endmodule


