*****************************
*     FPGA SPICE Netlist    *
* Description: Channel Y-direction  [1][1] in FPGA *
*    Author: Xifan TANG     *
* Organization: EPFL/IC/LSI *
* Date: Thu Nov 15 14:26:04 2018
 *
*****************************
***** Subckt for Channel Y [1][1] *****
.subckt chany[1][1] 
+ in0 out1 in2 out3 in4 out5 in6 out7 in8 out9 in10 out11 in12 out13 in14 out15 in16 out17 in18 out19 in20 out21 in22 out23 in24 out25 in26 out27 in28 out29 
+ out0 in1 out2 in3 out4 in5 out6 in7 out8 in9 out10 in11 out12 in13 out14 in15 out16 in17 out18 in19 out20 in21 out22 in23 out24 in25 out26 in27 out28 in29 
+ mid_out0 mid_out1 mid_out2 mid_out3 mid_out4 mid_out5 mid_out6 mid_out7 mid_out8 mid_out9 mid_out10 mid_out11 mid_out12 mid_out13 mid_out14 mid_out15 mid_out16 mid_out17 mid_out18 mid_out19 mid_out20 mid_out21 mid_out22 mid_out23 mid_out24 mid_out25 mid_out26 mid_out27 mid_out28 mid_out29 
+ svdd sgnd
Xtrack_seg[90] in0 out0 mid_out0 svdd sgnd chan_segment_seg0
Xtrack_seg[91] in1 out1 mid_out1 svdd sgnd chan_segment_seg0
Xtrack_seg[92] in2 out2 mid_out2 svdd sgnd chan_segment_seg0
Xtrack_seg[93] in3 out3 mid_out3 svdd sgnd chan_segment_seg0
Xtrack_seg[94] in4 out4 mid_out4 svdd sgnd chan_segment_seg0
Xtrack_seg[95] in5 out5 mid_out5 svdd sgnd chan_segment_seg0
Xtrack_seg[96] in6 out6 mid_out6 svdd sgnd chan_segment_seg0
Xtrack_seg[97] in7 out7 mid_out7 svdd sgnd chan_segment_seg0
Xtrack_seg[98] in8 out8 mid_out8 svdd sgnd chan_segment_seg0
Xtrack_seg[99] in9 out9 mid_out9 svdd sgnd chan_segment_seg0
Xtrack_seg[100] in10 out10 mid_out10 svdd sgnd chan_segment_seg0
Xtrack_seg[101] in11 out11 mid_out11 svdd sgnd chan_segment_seg0
Xtrack_seg[102] in12 out12 mid_out12 svdd sgnd chan_segment_seg1
Xtrack_seg[103] in13 out13 mid_out13 svdd sgnd chan_segment_seg1
Xtrack_seg[104] in14 out14 mid_out14 svdd sgnd chan_segment_seg1
Xtrack_seg[105] in15 out15 mid_out15 svdd sgnd chan_segment_seg1
Xtrack_seg[106] in16 out16 mid_out16 svdd sgnd chan_segment_seg1
Xtrack_seg[107] in17 out17 mid_out17 svdd sgnd chan_segment_seg1
Xtrack_seg[108] in18 out18 mid_out18 svdd sgnd chan_segment_seg1
Xtrack_seg[109] in19 out19 mid_out19 svdd sgnd chan_segment_seg1
Xtrack_seg[110] in20 out20 mid_out20 svdd sgnd chan_segment_seg1
Xtrack_seg[111] in21 out21 mid_out21 svdd sgnd chan_segment_seg1
Xtrack_seg[112] in22 out22 mid_out22 svdd sgnd chan_segment_seg2
Xtrack_seg[113] in23 out23 mid_out23 svdd sgnd chan_segment_seg2
Xtrack_seg[114] in24 out24 mid_out24 svdd sgnd chan_segment_seg2
Xtrack_seg[115] in25 out25 mid_out25 svdd sgnd chan_segment_seg2
Xtrack_seg[116] in26 out26 mid_out26 svdd sgnd chan_segment_seg2
Xtrack_seg[117] in27 out27 mid_out27 svdd sgnd chan_segment_seg2
Xtrack_seg[118] in28 out28 mid_out28 svdd sgnd chan_segment_seg2
Xtrack_seg[119] in29 out29 mid_out29 svdd sgnd chan_segment_seg2
.eom
