*****************************
*     FPGA SPICE Netlist    *
* Description: Connection Block X-channel  [1][1] in FPGA *
*    Author: Xifan TANG     *
* Organization: EPFL/IC/LSI *
* Date: Thu Nov 15 14:26:08 2018
 *
*****************************
.subckt cbx[1][1] 
+ chanx[1][1]_midout[0] 
+ chanx[1][1]_midout[1] 
+ chanx[1][1]_midout[2] 
+ chanx[1][1]_midout[3] 
+ chanx[1][1]_midout[4] 
+ chanx[1][1]_midout[5] 
+ chanx[1][1]_midout[6] 
+ chanx[1][1]_midout[7] 
+ chanx[1][1]_midout[8] 
+ chanx[1][1]_midout[9] 
+ chanx[1][1]_midout[10] 
+ chanx[1][1]_midout[11] 
+ chanx[1][1]_midout[12] 
+ chanx[1][1]_midout[13] 
+ chanx[1][1]_midout[14] 
+ chanx[1][1]_midout[15] 
+ chanx[1][1]_midout[16] 
+ chanx[1][1]_midout[17] 
+ chanx[1][1]_midout[18] 
+ chanx[1][1]_midout[19] 
+ chanx[1][1]_midout[20] 
+ chanx[1][1]_midout[21] 
+ chanx[1][1]_midout[22] 
+ chanx[1][1]_midout[23] 
+ chanx[1][1]_midout[24] 
+ chanx[1][1]_midout[25] 
+ chanx[1][1]_midout[26] 
+ chanx[1][1]_midout[27] 
+ chanx[1][1]_midout[28] 
+ chanx[1][1]_midout[29] 
+ chanx[1][1]_midout[30] 
+ chanx[1][1]_midout[31] 
+ chanx[1][1]_midout[32] 
+ chanx[1][1]_midout[33] 
+ chanx[1][1]_midout[34] 
+ chanx[1][1]_midout[35] 
+ chanx[1][1]_midout[36] 
+ chanx[1][1]_midout[37] 
+ chanx[1][1]_midout[38] 
+ chanx[1][1]_midout[39] 
+ chanx[1][1]_midout[40] 
+ chanx[1][1]_midout[41] 
+ chanx[1][1]_midout[42] 
+ chanx[1][1]_midout[43] 
+ chanx[1][1]_midout[44] 
+ chanx[1][1]_midout[45] 
+ chanx[1][1]_midout[46] 
+ chanx[1][1]_midout[47] 
+ chanx[1][1]_midout[48] 
+ chanx[1][1]_midout[49] 
+ chanx[1][1]_midout[50] 
+ chanx[1][1]_midout[51] 
+ chanx[1][1]_midout[52] 
+ chanx[1][1]_midout[53] 
+ chanx[1][1]_midout[54] 
+ chanx[1][1]_midout[55] 
+ chanx[1][1]_midout[56] 
+ chanx[1][1]_midout[57] 
+ chanx[1][1]_midout[58] 
+ chanx[1][1]_midout[59] 
+ chanx[1][1]_midout[60] 
+ chanx[1][1]_midout[61] 
+ chanx[1][1]_midout[62] 
+ chanx[1][1]_midout[63] 
+ chanx[1][1]_midout[64] 
+ chanx[1][1]_midout[65] 
+ chanx[1][1]_midout[66] 
+ chanx[1][1]_midout[67] 
+ chanx[1][1]_midout[68] 
+ chanx[1][1]_midout[69] 
+ chanx[1][1]_midout[70] 
+ chanx[1][1]_midout[71] 
+ chanx[1][1]_midout[72] 
+ chanx[1][1]_midout[73] 
+ chanx[1][1]_midout[74] 
+ chanx[1][1]_midout[75] 
+ chanx[1][1]_midout[76] 
+ chanx[1][1]_midout[77] 
+ chanx[1][1]_midout[78] 
+ chanx[1][1]_midout[79] 
+ chanx[1][1]_midout[80] 
+ chanx[1][1]_midout[81] 
+ chanx[1][1]_midout[82] 
+ chanx[1][1]_midout[83] 
+ chanx[1][1]_midout[84] 
+ chanx[1][1]_midout[85] 
+ chanx[1][1]_midout[86] 
+ chanx[1][1]_midout[87] 
+ chanx[1][1]_midout[88] 
+ chanx[1][1]_midout[89] 
+ chanx[1][1]_midout[90] 
+ chanx[1][1]_midout[91] 
+ chanx[1][1]_midout[92] 
+ chanx[1][1]_midout[93] 
+ chanx[1][1]_midout[94] 
+ chanx[1][1]_midout[95] 
+ chanx[1][1]_midout[96] 
+ chanx[1][1]_midout[97] 
+ chanx[1][1]_midout[98] 
+ chanx[1][1]_midout[99] 
+ grid[1][2]_pin[0][2][0] 
+ grid[1][2]_pin[0][2][2] 
+ grid[1][2]_pin[0][2][4] 
+ grid[1][2]_pin[0][2][6] 
+ grid[1][2]_pin[0][2][8] 
+ grid[1][2]_pin[0][2][10] 
+ grid[1][2]_pin[0][2][12] 
+ grid[1][2]_pin[0][2][14] 
+ grid[1][1]_pin[0][0][0] 
+ grid[1][1]_pin[0][0][4] 
+ grid[1][1]_pin[0][0][8] 
+ grid[1][1]_pin[0][0][12] 
+ grid[1][1]_pin[0][0][16] 
+ grid[1][1]_pin[0][0][20] 
+ grid[1][1]_pin[0][0][24] 
+ grid[1][1]_pin[0][0][28] 
+ grid[1][1]_pin[0][0][32] 
+ grid[1][1]_pin[0][0][36] 
+ svdd sgnd
Xmux_2level_tapbuf_size16[18] chanx[1][1]_midout[6] chanx[1][1]_midout[7] chanx[1][1]_midout[10] chanx[1][1]_midout[11] chanx[1][1]_midout[30] chanx[1][1]_midout[31] chanx[1][1]_midout[36] chanx[1][1]_midout[37] chanx[1][1]_midout[48] chanx[1][1]_midout[49] chanx[1][1]_midout[60] chanx[1][1]_midout[61] chanx[1][1]_midout[74] chanx[1][1]_midout[75] chanx[1][1]_midout[88] chanx[1][1]_midout[89] grid[1][2]_pin[0][2][0] sram[2226]->outb sram[2226]->out sram[2227]->out sram[2227]->outb sram[2228]->out sram[2228]->outb sram[2229]->out sram[2229]->outb sram[2230]->outb sram[2230]->out sram[2231]->out sram[2231]->outb sram[2232]->out sram[2232]->outb sram[2233]->out sram[2233]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[18], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2226] sram->in sram[2226]->out sram[2226]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2226]->out) 0
.nodeset V(sram[2226]->outb) vsp
Xsram[2227] sram->in sram[2227]->out sram[2227]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2227]->out) 0
.nodeset V(sram[2227]->outb) vsp
Xsram[2228] sram->in sram[2228]->out sram[2228]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2228]->out) 0
.nodeset V(sram[2228]->outb) vsp
Xsram[2229] sram->in sram[2229]->out sram[2229]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2229]->out) 0
.nodeset V(sram[2229]->outb) vsp
Xsram[2230] sram->in sram[2230]->out sram[2230]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2230]->out) 0
.nodeset V(sram[2230]->outb) vsp
Xsram[2231] sram->in sram[2231]->out sram[2231]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2231]->out) 0
.nodeset V(sram[2231]->outb) vsp
Xsram[2232] sram->in sram[2232]->out sram[2232]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2232]->out) 0
.nodeset V(sram[2232]->outb) vsp
Xsram[2233] sram->in sram[2233]->out sram[2233]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2233]->out) 0
.nodeset V(sram[2233]->outb) vsp
Xmux_2level_tapbuf_size16[19] chanx[1][1]_midout[0] chanx[1][1]_midout[1] chanx[1][1]_midout[12] chanx[1][1]_midout[13] chanx[1][1]_midout[24] chanx[1][1]_midout[25] chanx[1][1]_midout[36] chanx[1][1]_midout[37] chanx[1][1]_midout[54] chanx[1][1]_midout[55] chanx[1][1]_midout[66] chanx[1][1]_midout[67] chanx[1][1]_midout[76] chanx[1][1]_midout[77] chanx[1][1]_midout[88] chanx[1][1]_midout[89] grid[1][2]_pin[0][2][2] sram[2234]->outb sram[2234]->out sram[2235]->out sram[2235]->outb sram[2236]->out sram[2236]->outb sram[2237]->out sram[2237]->outb sram[2238]->outb sram[2238]->out sram[2239]->out sram[2239]->outb sram[2240]->out sram[2240]->outb sram[2241]->out sram[2241]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[19], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2234] sram->in sram[2234]->out sram[2234]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2234]->out) 0
.nodeset V(sram[2234]->outb) vsp
Xsram[2235] sram->in sram[2235]->out sram[2235]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2235]->out) 0
.nodeset V(sram[2235]->outb) vsp
Xsram[2236] sram->in sram[2236]->out sram[2236]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2236]->out) 0
.nodeset V(sram[2236]->outb) vsp
Xsram[2237] sram->in sram[2237]->out sram[2237]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2237]->out) 0
.nodeset V(sram[2237]->outb) vsp
Xsram[2238] sram->in sram[2238]->out sram[2238]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2238]->out) 0
.nodeset V(sram[2238]->outb) vsp
Xsram[2239] sram->in sram[2239]->out sram[2239]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2239]->out) 0
.nodeset V(sram[2239]->outb) vsp
Xsram[2240] sram->in sram[2240]->out sram[2240]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2240]->out) 0
.nodeset V(sram[2240]->outb) vsp
Xsram[2241] sram->in sram[2241]->out sram[2241]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2241]->out) 0
.nodeset V(sram[2241]->outb) vsp
Xmux_2level_tapbuf_size16[20] chanx[1][1]_midout[0] chanx[1][1]_midout[1] chanx[1][1]_midout[22] chanx[1][1]_midout[23] chanx[1][1]_midout[26] chanx[1][1]_midout[27] chanx[1][1]_midout[42] chanx[1][1]_midout[43] chanx[1][1]_midout[54] chanx[1][1]_midout[55] chanx[1][1]_midout[64] chanx[1][1]_midout[65] chanx[1][1]_midout[78] chanx[1][1]_midout[79] chanx[1][1]_midout[90] chanx[1][1]_midout[91] grid[1][2]_pin[0][2][4] sram[2242]->outb sram[2242]->out sram[2243]->out sram[2243]->outb sram[2244]->out sram[2244]->outb sram[2245]->out sram[2245]->outb sram[2246]->outb sram[2246]->out sram[2247]->out sram[2247]->outb sram[2248]->out sram[2248]->outb sram[2249]->out sram[2249]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[20], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2242] sram->in sram[2242]->out sram[2242]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2242]->out) 0
.nodeset V(sram[2242]->outb) vsp
Xsram[2243] sram->in sram[2243]->out sram[2243]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2243]->out) 0
.nodeset V(sram[2243]->outb) vsp
Xsram[2244] sram->in sram[2244]->out sram[2244]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2244]->out) 0
.nodeset V(sram[2244]->outb) vsp
Xsram[2245] sram->in sram[2245]->out sram[2245]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2245]->out) 0
.nodeset V(sram[2245]->outb) vsp
Xsram[2246] sram->in sram[2246]->out sram[2246]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2246]->out) 0
.nodeset V(sram[2246]->outb) vsp
Xsram[2247] sram->in sram[2247]->out sram[2247]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2247]->out) 0
.nodeset V(sram[2247]->outb) vsp
Xsram[2248] sram->in sram[2248]->out sram[2248]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2248]->out) 0
.nodeset V(sram[2248]->outb) vsp
Xsram[2249] sram->in sram[2249]->out sram[2249]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2249]->out) 0
.nodeset V(sram[2249]->outb) vsp
Xmux_2level_tapbuf_size16[21] chanx[1][1]_midout[2] chanx[1][1]_midout[3] chanx[1][1]_midout[22] chanx[1][1]_midout[23] chanx[1][1]_midout[28] chanx[1][1]_midout[29] chanx[1][1]_midout[40] chanx[1][1]_midout[41] chanx[1][1]_midout[52] chanx[1][1]_midout[53] chanx[1][1]_midout[64] chanx[1][1]_midout[65] chanx[1][1]_midout[80] chanx[1][1]_midout[81] chanx[1][1]_midout[92] chanx[1][1]_midout[93] grid[1][2]_pin[0][2][6] sram[2250]->outb sram[2250]->out sram[2251]->out sram[2251]->outb sram[2252]->out sram[2252]->outb sram[2253]->out sram[2253]->outb sram[2254]->outb sram[2254]->out sram[2255]->out sram[2255]->outb sram[2256]->out sram[2256]->outb sram[2257]->out sram[2257]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[21], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2250] sram->in sram[2250]->out sram[2250]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2250]->out) 0
.nodeset V(sram[2250]->outb) vsp
Xsram[2251] sram->in sram[2251]->out sram[2251]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2251]->out) 0
.nodeset V(sram[2251]->outb) vsp
Xsram[2252] sram->in sram[2252]->out sram[2252]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2252]->out) 0
.nodeset V(sram[2252]->outb) vsp
Xsram[2253] sram->in sram[2253]->out sram[2253]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2253]->out) 0
.nodeset V(sram[2253]->outb) vsp
Xsram[2254] sram->in sram[2254]->out sram[2254]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2254]->out) 0
.nodeset V(sram[2254]->outb) vsp
Xsram[2255] sram->in sram[2255]->out sram[2255]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2255]->out) 0
.nodeset V(sram[2255]->outb) vsp
Xsram[2256] sram->in sram[2256]->out sram[2256]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2256]->out) 0
.nodeset V(sram[2256]->outb) vsp
Xsram[2257] sram->in sram[2257]->out sram[2257]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2257]->out) 0
.nodeset V(sram[2257]->outb) vsp
Xmux_2level_tapbuf_size16[22] chanx[1][1]_midout[4] chanx[1][1]_midout[5] chanx[1][1]_midout[16] chanx[1][1]_midout[17] chanx[1][1]_midout[38] chanx[1][1]_midout[39] chanx[1][1]_midout[46] chanx[1][1]_midout[47] chanx[1][1]_midout[58] chanx[1][1]_midout[59] chanx[1][1]_midout[68] chanx[1][1]_midout[69] chanx[1][1]_midout[82] chanx[1][1]_midout[83] chanx[1][1]_midout[94] chanx[1][1]_midout[95] grid[1][2]_pin[0][2][8] sram[2258]->outb sram[2258]->out sram[2259]->out sram[2259]->outb sram[2260]->out sram[2260]->outb sram[2261]->out sram[2261]->outb sram[2262]->outb sram[2262]->out sram[2263]->out sram[2263]->outb sram[2264]->out sram[2264]->outb sram[2265]->out sram[2265]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[22], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2258] sram->in sram[2258]->out sram[2258]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2258]->out) 0
.nodeset V(sram[2258]->outb) vsp
Xsram[2259] sram->in sram[2259]->out sram[2259]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2259]->out) 0
.nodeset V(sram[2259]->outb) vsp
Xsram[2260] sram->in sram[2260]->out sram[2260]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2260]->out) 0
.nodeset V(sram[2260]->outb) vsp
Xsram[2261] sram->in sram[2261]->out sram[2261]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2261]->out) 0
.nodeset V(sram[2261]->outb) vsp
Xsram[2262] sram->in sram[2262]->out sram[2262]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2262]->out) 0
.nodeset V(sram[2262]->outb) vsp
Xsram[2263] sram->in sram[2263]->out sram[2263]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2263]->out) 0
.nodeset V(sram[2263]->outb) vsp
Xsram[2264] sram->in sram[2264]->out sram[2264]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2264]->out) 0
.nodeset V(sram[2264]->outb) vsp
Xsram[2265] sram->in sram[2265]->out sram[2265]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2265]->out) 0
.nodeset V(sram[2265]->outb) vsp
Xmux_2level_tapbuf_size16[23] chanx[1][1]_midout[14] chanx[1][1]_midout[15] chanx[1][1]_midout[18] chanx[1][1]_midout[19] chanx[1][1]_midout[38] chanx[1][1]_midout[39] chanx[1][1]_midout[44] chanx[1][1]_midout[45] chanx[1][1]_midout[56] chanx[1][1]_midout[57] chanx[1][1]_midout[70] chanx[1][1]_midout[71] chanx[1][1]_midout[82] chanx[1][1]_midout[83] chanx[1][1]_midout[96] chanx[1][1]_midout[97] grid[1][2]_pin[0][2][10] sram[2266]->outb sram[2266]->out sram[2267]->out sram[2267]->outb sram[2268]->out sram[2268]->outb sram[2269]->out sram[2269]->outb sram[2270]->outb sram[2270]->out sram[2271]->out sram[2271]->outb sram[2272]->out sram[2272]->outb sram[2273]->out sram[2273]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[23], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2266] sram->in sram[2266]->out sram[2266]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2266]->out) 0
.nodeset V(sram[2266]->outb) vsp
Xsram[2267] sram->in sram[2267]->out sram[2267]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2267]->out) 0
.nodeset V(sram[2267]->outb) vsp
Xsram[2268] sram->in sram[2268]->out sram[2268]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2268]->out) 0
.nodeset V(sram[2268]->outb) vsp
Xsram[2269] sram->in sram[2269]->out sram[2269]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2269]->out) 0
.nodeset V(sram[2269]->outb) vsp
Xsram[2270] sram->in sram[2270]->out sram[2270]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2270]->out) 0
.nodeset V(sram[2270]->outb) vsp
Xsram[2271] sram->in sram[2271]->out sram[2271]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2271]->out) 0
.nodeset V(sram[2271]->outb) vsp
Xsram[2272] sram->in sram[2272]->out sram[2272]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2272]->out) 0
.nodeset V(sram[2272]->outb) vsp
Xsram[2273] sram->in sram[2273]->out sram[2273]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2273]->out) 0
.nodeset V(sram[2273]->outb) vsp
Xmux_2level_tapbuf_size16[24] chanx[1][1]_midout[8] chanx[1][1]_midout[9] chanx[1][1]_midout[20] chanx[1][1]_midout[21] chanx[1][1]_midout[32] chanx[1][1]_midout[33] chanx[1][1]_midout[44] chanx[1][1]_midout[45] chanx[1][1]_midout[62] chanx[1][1]_midout[63] chanx[1][1]_midout[72] chanx[1][1]_midout[73] chanx[1][1]_midout[84] chanx[1][1]_midout[85] chanx[1][1]_midout[96] chanx[1][1]_midout[97] grid[1][2]_pin[0][2][12] sram[2274]->outb sram[2274]->out sram[2275]->out sram[2275]->outb sram[2276]->out sram[2276]->outb sram[2277]->out sram[2277]->outb sram[2278]->out sram[2278]->outb sram[2279]->out sram[2279]->outb sram[2280]->outb sram[2280]->out sram[2281]->out sram[2281]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[24], level=2, select_path_id=2. *****
*****10000010*****
Xsram[2274] sram->in sram[2274]->out sram[2274]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2274]->out) 0
.nodeset V(sram[2274]->outb) vsp
Xsram[2275] sram->in sram[2275]->out sram[2275]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2275]->out) 0
.nodeset V(sram[2275]->outb) vsp
Xsram[2276] sram->in sram[2276]->out sram[2276]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2276]->out) 0
.nodeset V(sram[2276]->outb) vsp
Xsram[2277] sram->in sram[2277]->out sram[2277]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2277]->out) 0
.nodeset V(sram[2277]->outb) vsp
Xsram[2278] sram->in sram[2278]->out sram[2278]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2278]->out) 0
.nodeset V(sram[2278]->outb) vsp
Xsram[2279] sram->in sram[2279]->out sram[2279]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2279]->out) 0
.nodeset V(sram[2279]->outb) vsp
Xsram[2280] sram->in sram[2280]->out sram[2280]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2280]->out) 0
.nodeset V(sram[2280]->outb) vsp
Xsram[2281] sram->in sram[2281]->out sram[2281]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2281]->out) 0
.nodeset V(sram[2281]->outb) vsp
Xmux_2level_tapbuf_size16[25] chanx[1][1]_midout[8] chanx[1][1]_midout[9] chanx[1][1]_midout[30] chanx[1][1]_midout[31] chanx[1][1]_midout[34] chanx[1][1]_midout[35] chanx[1][1]_midout[50] chanx[1][1]_midout[51] chanx[1][1]_midout[62] chanx[1][1]_midout[63] chanx[1][1]_midout[74] chanx[1][1]_midout[75] chanx[1][1]_midout[86] chanx[1][1]_midout[87] chanx[1][1]_midout[98] chanx[1][1]_midout[99] grid[1][2]_pin[0][2][14] sram[2282]->outb sram[2282]->out sram[2283]->out sram[2283]->outb sram[2284]->out sram[2284]->outb sram[2285]->out sram[2285]->outb sram[2286]->outb sram[2286]->out sram[2287]->out sram[2287]->outb sram[2288]->out sram[2288]->outb sram[2289]->out sram[2289]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[25], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2282] sram->in sram[2282]->out sram[2282]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2282]->out) 0
.nodeset V(sram[2282]->outb) vsp
Xsram[2283] sram->in sram[2283]->out sram[2283]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2283]->out) 0
.nodeset V(sram[2283]->outb) vsp
Xsram[2284] sram->in sram[2284]->out sram[2284]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2284]->out) 0
.nodeset V(sram[2284]->outb) vsp
Xsram[2285] sram->in sram[2285]->out sram[2285]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2285]->out) 0
.nodeset V(sram[2285]->outb) vsp
Xsram[2286] sram->in sram[2286]->out sram[2286]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2286]->out) 0
.nodeset V(sram[2286]->outb) vsp
Xsram[2287] sram->in sram[2287]->out sram[2287]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2287]->out) 0
.nodeset V(sram[2287]->outb) vsp
Xsram[2288] sram->in sram[2288]->out sram[2288]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2288]->out) 0
.nodeset V(sram[2288]->outb) vsp
Xsram[2289] sram->in sram[2289]->out sram[2289]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2289]->out) 0
.nodeset V(sram[2289]->outb) vsp
Xmux_2level_tapbuf_size16[26] chanx[1][1]_midout[6] chanx[1][1]_midout[7] chanx[1][1]_midout[10] chanx[1][1]_midout[11] chanx[1][1]_midout[30] chanx[1][1]_midout[31] chanx[1][1]_midout[34] chanx[1][1]_midout[35] chanx[1][1]_midout[48] chanx[1][1]_midout[49] chanx[1][1]_midout[60] chanx[1][1]_midout[61] chanx[1][1]_midout[74] chanx[1][1]_midout[75] chanx[1][1]_midout[86] chanx[1][1]_midout[87] grid[1][1]_pin[0][0][0] sram[2290]->outb sram[2290]->out sram[2291]->out sram[2291]->outb sram[2292]->out sram[2292]->outb sram[2293]->out sram[2293]->outb sram[2294]->outb sram[2294]->out sram[2295]->out sram[2295]->outb sram[2296]->out sram[2296]->outb sram[2297]->out sram[2297]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[26], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2290] sram->in sram[2290]->out sram[2290]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2290]->out) 0
.nodeset V(sram[2290]->outb) vsp
Xsram[2291] sram->in sram[2291]->out sram[2291]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2291]->out) 0
.nodeset V(sram[2291]->outb) vsp
Xsram[2292] sram->in sram[2292]->out sram[2292]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2292]->out) 0
.nodeset V(sram[2292]->outb) vsp
Xsram[2293] sram->in sram[2293]->out sram[2293]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2293]->out) 0
.nodeset V(sram[2293]->outb) vsp
Xsram[2294] sram->in sram[2294]->out sram[2294]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2294]->out) 0
.nodeset V(sram[2294]->outb) vsp
Xsram[2295] sram->in sram[2295]->out sram[2295]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2295]->out) 0
.nodeset V(sram[2295]->outb) vsp
Xsram[2296] sram->in sram[2296]->out sram[2296]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2296]->out) 0
.nodeset V(sram[2296]->outb) vsp
Xsram[2297] sram->in sram[2297]->out sram[2297]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2297]->out) 0
.nodeset V(sram[2297]->outb) vsp
Xmux_2level_tapbuf_size16[27] chanx[1][1]_midout[6] chanx[1][1]_midout[7] chanx[1][1]_midout[10] chanx[1][1]_midout[11] chanx[1][1]_midout[24] chanx[1][1]_midout[25] chanx[1][1]_midout[36] chanx[1][1]_midout[37] chanx[1][1]_midout[48] chanx[1][1]_midout[49] chanx[1][1]_midout[60] chanx[1][1]_midout[61] chanx[1][1]_midout[76] chanx[1][1]_midout[77] chanx[1][1]_midout[88] chanx[1][1]_midout[89] grid[1][1]_pin[0][0][4] sram[2298]->outb sram[2298]->out sram[2299]->out sram[2299]->outb sram[2300]->out sram[2300]->outb sram[2301]->out sram[2301]->outb sram[2302]->outb sram[2302]->out sram[2303]->out sram[2303]->outb sram[2304]->out sram[2304]->outb sram[2305]->out sram[2305]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[27], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2298] sram->in sram[2298]->out sram[2298]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2298]->out) 0
.nodeset V(sram[2298]->outb) vsp
Xsram[2299] sram->in sram[2299]->out sram[2299]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2299]->out) 0
.nodeset V(sram[2299]->outb) vsp
Xsram[2300] sram->in sram[2300]->out sram[2300]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2300]->out) 0
.nodeset V(sram[2300]->outb) vsp
Xsram[2301] sram->in sram[2301]->out sram[2301]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2301]->out) 0
.nodeset V(sram[2301]->outb) vsp
Xsram[2302] sram->in sram[2302]->out sram[2302]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2302]->out) 0
.nodeset V(sram[2302]->outb) vsp
Xsram[2303] sram->in sram[2303]->out sram[2303]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2303]->out) 0
.nodeset V(sram[2303]->outb) vsp
Xsram[2304] sram->in sram[2304]->out sram[2304]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2304]->out) 0
.nodeset V(sram[2304]->outb) vsp
Xsram[2305] sram->in sram[2305]->out sram[2305]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2305]->out) 0
.nodeset V(sram[2305]->outb) vsp
Xmux_2level_tapbuf_size16[28] chanx[1][1]_midout[0] chanx[1][1]_midout[1] chanx[1][1]_midout[12] chanx[1][1]_midout[13] chanx[1][1]_midout[24] chanx[1][1]_midout[25] chanx[1][1]_midout[42] chanx[1][1]_midout[43] chanx[1][1]_midout[54] chanx[1][1]_midout[55] chanx[1][1]_midout[66] chanx[1][1]_midout[67] chanx[1][1]_midout[76] chanx[1][1]_midout[77] chanx[1][1]_midout[90] chanx[1][1]_midout[91] grid[1][1]_pin[0][0][8] sram[2306]->outb sram[2306]->out sram[2307]->out sram[2307]->outb sram[2308]->out sram[2308]->outb sram[2309]->out sram[2309]->outb sram[2310]->outb sram[2310]->out sram[2311]->out sram[2311]->outb sram[2312]->out sram[2312]->outb sram[2313]->out sram[2313]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[28], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2306] sram->in sram[2306]->out sram[2306]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2306]->out) 0
.nodeset V(sram[2306]->outb) vsp
Xsram[2307] sram->in sram[2307]->out sram[2307]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2307]->out) 0
.nodeset V(sram[2307]->outb) vsp
Xsram[2308] sram->in sram[2308]->out sram[2308]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2308]->out) 0
.nodeset V(sram[2308]->outb) vsp
Xsram[2309] sram->in sram[2309]->out sram[2309]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2309]->out) 0
.nodeset V(sram[2309]->outb) vsp
Xsram[2310] sram->in sram[2310]->out sram[2310]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2310]->out) 0
.nodeset V(sram[2310]->outb) vsp
Xsram[2311] sram->in sram[2311]->out sram[2311]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2311]->out) 0
.nodeset V(sram[2311]->outb) vsp
Xsram[2312] sram->in sram[2312]->out sram[2312]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2312]->out) 0
.nodeset V(sram[2312]->outb) vsp
Xsram[2313] sram->in sram[2313]->out sram[2313]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2313]->out) 0
.nodeset V(sram[2313]->outb) vsp
Xmux_2level_tapbuf_size16[29] chanx[1][1]_midout[0] chanx[1][1]_midout[1] chanx[1][1]_midout[22] chanx[1][1]_midout[23] chanx[1][1]_midout[26] chanx[1][1]_midout[27] chanx[1][1]_midout[42] chanx[1][1]_midout[43] chanx[1][1]_midout[54] chanx[1][1]_midout[55] chanx[1][1]_midout[64] chanx[1][1]_midout[65] chanx[1][1]_midout[78] chanx[1][1]_midout[79] chanx[1][1]_midout[90] chanx[1][1]_midout[91] grid[1][1]_pin[0][0][12] sram[2314]->outb sram[2314]->out sram[2315]->out sram[2315]->outb sram[2316]->out sram[2316]->outb sram[2317]->out sram[2317]->outb sram[2318]->outb sram[2318]->out sram[2319]->out sram[2319]->outb sram[2320]->out sram[2320]->outb sram[2321]->out sram[2321]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[29], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2314] sram->in sram[2314]->out sram[2314]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2314]->out) 0
.nodeset V(sram[2314]->outb) vsp
Xsram[2315] sram->in sram[2315]->out sram[2315]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2315]->out) 0
.nodeset V(sram[2315]->outb) vsp
Xsram[2316] sram->in sram[2316]->out sram[2316]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2316]->out) 0
.nodeset V(sram[2316]->outb) vsp
Xsram[2317] sram->in sram[2317]->out sram[2317]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2317]->out) 0
.nodeset V(sram[2317]->outb) vsp
Xsram[2318] sram->in sram[2318]->out sram[2318]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2318]->out) 0
.nodeset V(sram[2318]->outb) vsp
Xsram[2319] sram->in sram[2319]->out sram[2319]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2319]->out) 0
.nodeset V(sram[2319]->outb) vsp
Xsram[2320] sram->in sram[2320]->out sram[2320]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2320]->out) 0
.nodeset V(sram[2320]->outb) vsp
Xsram[2321] sram->in sram[2321]->out sram[2321]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2321]->out) 0
.nodeset V(sram[2321]->outb) vsp
Xmux_2level_tapbuf_size16[30] chanx[1][1]_midout[2] chanx[1][1]_midout[3] chanx[1][1]_midout[22] chanx[1][1]_midout[23] chanx[1][1]_midout[28] chanx[1][1]_midout[29] chanx[1][1]_midout[40] chanx[1][1]_midout[41] chanx[1][1]_midout[52] chanx[1][1]_midout[53] chanx[1][1]_midout[64] chanx[1][1]_midout[65] chanx[1][1]_midout[80] chanx[1][1]_midout[81] chanx[1][1]_midout[92] chanx[1][1]_midout[93] grid[1][1]_pin[0][0][16] sram[2322]->outb sram[2322]->out sram[2323]->out sram[2323]->outb sram[2324]->out sram[2324]->outb sram[2325]->out sram[2325]->outb sram[2326]->outb sram[2326]->out sram[2327]->out sram[2327]->outb sram[2328]->out sram[2328]->outb sram[2329]->out sram[2329]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[30], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2322] sram->in sram[2322]->out sram[2322]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2322]->out) 0
.nodeset V(sram[2322]->outb) vsp
Xsram[2323] sram->in sram[2323]->out sram[2323]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2323]->out) 0
.nodeset V(sram[2323]->outb) vsp
Xsram[2324] sram->in sram[2324]->out sram[2324]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2324]->out) 0
.nodeset V(sram[2324]->outb) vsp
Xsram[2325] sram->in sram[2325]->out sram[2325]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2325]->out) 0
.nodeset V(sram[2325]->outb) vsp
Xsram[2326] sram->in sram[2326]->out sram[2326]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2326]->out) 0
.nodeset V(sram[2326]->outb) vsp
Xsram[2327] sram->in sram[2327]->out sram[2327]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2327]->out) 0
.nodeset V(sram[2327]->outb) vsp
Xsram[2328] sram->in sram[2328]->out sram[2328]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2328]->out) 0
.nodeset V(sram[2328]->outb) vsp
Xsram[2329] sram->in sram[2329]->out sram[2329]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2329]->out) 0
.nodeset V(sram[2329]->outb) vsp
Xmux_2level_tapbuf_size16[31] chanx[1][1]_midout[4] chanx[1][1]_midout[5] chanx[1][1]_midout[16] chanx[1][1]_midout[17] chanx[1][1]_midout[28] chanx[1][1]_midout[29] chanx[1][1]_midout[40] chanx[1][1]_midout[41] chanx[1][1]_midout[58] chanx[1][1]_midout[59] chanx[1][1]_midout[68] chanx[1][1]_midout[69] chanx[1][1]_midout[80] chanx[1][1]_midout[81] chanx[1][1]_midout[92] chanx[1][1]_midout[93] grid[1][1]_pin[0][0][20] sram[2330]->outb sram[2330]->out sram[2331]->out sram[2331]->outb sram[2332]->out sram[2332]->outb sram[2333]->out sram[2333]->outb sram[2334]->outb sram[2334]->out sram[2335]->out sram[2335]->outb sram[2336]->out sram[2336]->outb sram[2337]->out sram[2337]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[31], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2330] sram->in sram[2330]->out sram[2330]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2330]->out) 0
.nodeset V(sram[2330]->outb) vsp
Xsram[2331] sram->in sram[2331]->out sram[2331]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2331]->out) 0
.nodeset V(sram[2331]->outb) vsp
Xsram[2332] sram->in sram[2332]->out sram[2332]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2332]->out) 0
.nodeset V(sram[2332]->outb) vsp
Xsram[2333] sram->in sram[2333]->out sram[2333]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2333]->out) 0
.nodeset V(sram[2333]->outb) vsp
Xsram[2334] sram->in sram[2334]->out sram[2334]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2334]->out) 0
.nodeset V(sram[2334]->outb) vsp
Xsram[2335] sram->in sram[2335]->out sram[2335]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2335]->out) 0
.nodeset V(sram[2335]->outb) vsp
Xsram[2336] sram->in sram[2336]->out sram[2336]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2336]->out) 0
.nodeset V(sram[2336]->outb) vsp
Xsram[2337] sram->in sram[2337]->out sram[2337]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2337]->out) 0
.nodeset V(sram[2337]->outb) vsp
Xmux_2level_tapbuf_size16[32] chanx[1][1]_midout[4] chanx[1][1]_midout[5] chanx[1][1]_midout[18] chanx[1][1]_midout[19] chanx[1][1]_midout[38] chanx[1][1]_midout[39] chanx[1][1]_midout[46] chanx[1][1]_midout[47] chanx[1][1]_midout[58] chanx[1][1]_midout[59] chanx[1][1]_midout[70] chanx[1][1]_midout[71] chanx[1][1]_midout[82] chanx[1][1]_midout[83] chanx[1][1]_midout[94] chanx[1][1]_midout[95] grid[1][1]_pin[0][0][24] sram[2338]->outb sram[2338]->out sram[2339]->out sram[2339]->outb sram[2340]->out sram[2340]->outb sram[2341]->out sram[2341]->outb sram[2342]->outb sram[2342]->out sram[2343]->out sram[2343]->outb sram[2344]->out sram[2344]->outb sram[2345]->out sram[2345]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[32], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2338] sram->in sram[2338]->out sram[2338]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2338]->out) 0
.nodeset V(sram[2338]->outb) vsp
Xsram[2339] sram->in sram[2339]->out sram[2339]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2339]->out) 0
.nodeset V(sram[2339]->outb) vsp
Xsram[2340] sram->in sram[2340]->out sram[2340]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2340]->out) 0
.nodeset V(sram[2340]->outb) vsp
Xsram[2341] sram->in sram[2341]->out sram[2341]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2341]->out) 0
.nodeset V(sram[2341]->outb) vsp
Xsram[2342] sram->in sram[2342]->out sram[2342]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2342]->out) 0
.nodeset V(sram[2342]->outb) vsp
Xsram[2343] sram->in sram[2343]->out sram[2343]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2343]->out) 0
.nodeset V(sram[2343]->outb) vsp
Xsram[2344] sram->in sram[2344]->out sram[2344]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2344]->out) 0
.nodeset V(sram[2344]->outb) vsp
Xsram[2345] sram->in sram[2345]->out sram[2345]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2345]->out) 0
.nodeset V(sram[2345]->outb) vsp
Xmux_2level_tapbuf_size16[33] chanx[1][1]_midout[14] chanx[1][1]_midout[15] chanx[1][1]_midout[18] chanx[1][1]_midout[19] chanx[1][1]_midout[38] chanx[1][1]_midout[39] chanx[1][1]_midout[44] chanx[1][1]_midout[45] chanx[1][1]_midout[56] chanx[1][1]_midout[57] chanx[1][1]_midout[70] chanx[1][1]_midout[71] chanx[1][1]_midout[82] chanx[1][1]_midout[83] chanx[1][1]_midout[96] chanx[1][1]_midout[97] grid[1][1]_pin[0][0][28] sram[2346]->outb sram[2346]->out sram[2347]->out sram[2347]->outb sram[2348]->out sram[2348]->outb sram[2349]->out sram[2349]->outb sram[2350]->outb sram[2350]->out sram[2351]->out sram[2351]->outb sram[2352]->out sram[2352]->outb sram[2353]->out sram[2353]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[33], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2346] sram->in sram[2346]->out sram[2346]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2346]->out) 0
.nodeset V(sram[2346]->outb) vsp
Xsram[2347] sram->in sram[2347]->out sram[2347]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2347]->out) 0
.nodeset V(sram[2347]->outb) vsp
Xsram[2348] sram->in sram[2348]->out sram[2348]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2348]->out) 0
.nodeset V(sram[2348]->outb) vsp
Xsram[2349] sram->in sram[2349]->out sram[2349]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2349]->out) 0
.nodeset V(sram[2349]->outb) vsp
Xsram[2350] sram->in sram[2350]->out sram[2350]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2350]->out) 0
.nodeset V(sram[2350]->outb) vsp
Xsram[2351] sram->in sram[2351]->out sram[2351]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2351]->out) 0
.nodeset V(sram[2351]->outb) vsp
Xsram[2352] sram->in sram[2352]->out sram[2352]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2352]->out) 0
.nodeset V(sram[2352]->outb) vsp
Xsram[2353] sram->in sram[2353]->out sram[2353]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2353]->out) 0
.nodeset V(sram[2353]->outb) vsp
Xmux_2level_tapbuf_size16[34] chanx[1][1]_midout[8] chanx[1][1]_midout[9] chanx[1][1]_midout[20] chanx[1][1]_midout[21] chanx[1][1]_midout[32] chanx[1][1]_midout[33] chanx[1][1]_midout[44] chanx[1][1]_midout[45] chanx[1][1]_midout[62] chanx[1][1]_midout[63] chanx[1][1]_midout[72] chanx[1][1]_midout[73] chanx[1][1]_midout[84] chanx[1][1]_midout[85] chanx[1][1]_midout[96] chanx[1][1]_midout[97] grid[1][1]_pin[0][0][32] sram[2354]->outb sram[2354]->out sram[2355]->out sram[2355]->outb sram[2356]->out sram[2356]->outb sram[2357]->out sram[2357]->outb sram[2358]->outb sram[2358]->out sram[2359]->out sram[2359]->outb sram[2360]->out sram[2360]->outb sram[2361]->out sram[2361]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[34], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2354] sram->in sram[2354]->out sram[2354]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2354]->out) 0
.nodeset V(sram[2354]->outb) vsp
Xsram[2355] sram->in sram[2355]->out sram[2355]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2355]->out) 0
.nodeset V(sram[2355]->outb) vsp
Xsram[2356] sram->in sram[2356]->out sram[2356]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2356]->out) 0
.nodeset V(sram[2356]->outb) vsp
Xsram[2357] sram->in sram[2357]->out sram[2357]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2357]->out) 0
.nodeset V(sram[2357]->outb) vsp
Xsram[2358] sram->in sram[2358]->out sram[2358]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2358]->out) 0
.nodeset V(sram[2358]->outb) vsp
Xsram[2359] sram->in sram[2359]->out sram[2359]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2359]->out) 0
.nodeset V(sram[2359]->outb) vsp
Xsram[2360] sram->in sram[2360]->out sram[2360]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2360]->out) 0
.nodeset V(sram[2360]->outb) vsp
Xsram[2361] sram->in sram[2361]->out sram[2361]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2361]->out) 0
.nodeset V(sram[2361]->outb) vsp
Xmux_2level_tapbuf_size16[35] chanx[1][1]_midout[8] chanx[1][1]_midout[9] chanx[1][1]_midout[20] chanx[1][1]_midout[21] chanx[1][1]_midout[34] chanx[1][1]_midout[35] chanx[1][1]_midout[50] chanx[1][1]_midout[51] chanx[1][1]_midout[62] chanx[1][1]_midout[63] chanx[1][1]_midout[72] chanx[1][1]_midout[73] chanx[1][1]_midout[86] chanx[1][1]_midout[87] chanx[1][1]_midout[98] chanx[1][1]_midout[99] grid[1][1]_pin[0][0][36] sram[2362]->outb sram[2362]->out sram[2363]->out sram[2363]->outb sram[2364]->out sram[2364]->outb sram[2365]->out sram[2365]->outb sram[2366]->outb sram[2366]->out sram[2367]->out sram[2367]->outb sram[2368]->out sram[2368]->outb sram[2369]->out sram[2369]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[35], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2362] sram->in sram[2362]->out sram[2362]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2362]->out) 0
.nodeset V(sram[2362]->outb) vsp
Xsram[2363] sram->in sram[2363]->out sram[2363]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2363]->out) 0
.nodeset V(sram[2363]->outb) vsp
Xsram[2364] sram->in sram[2364]->out sram[2364]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2364]->out) 0
.nodeset V(sram[2364]->outb) vsp
Xsram[2365] sram->in sram[2365]->out sram[2365]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2365]->out) 0
.nodeset V(sram[2365]->outb) vsp
Xsram[2366] sram->in sram[2366]->out sram[2366]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2366]->out) 0
.nodeset V(sram[2366]->outb) vsp
Xsram[2367] sram->in sram[2367]->out sram[2367]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2367]->out) 0
.nodeset V(sram[2367]->outb) vsp
Xsram[2368] sram->in sram[2368]->out sram[2368]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2368]->out) 0
.nodeset V(sram[2368]->outb) vsp
Xsram[2369] sram->in sram[2369]->out sram[2369]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2369]->out) 0
.nodeset V(sram[2369]->outb) vsp
.eom
