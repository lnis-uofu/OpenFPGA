


module bindfile;
	bind ADD_SUB sva_checker sva_checker_inst(.*);
endmodule
