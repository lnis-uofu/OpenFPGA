*****************************
*     FPGA SPICE Netlist    *
* Description: Logic Block [1][1] in FPGA *
*    Author: Xifan TANG     *
* Organization: EPFL/IC/LSI *
* Date: Thu Nov 15 14:26:08 2018
 *
*****************************
***** Grid[1][1] type_descriptor: clb[0] *****
.subckt grid[1][1]_clb[0]_mode[clb]_fle[0]_mode[n1_lut6]_ble6[0]_mode[ble6]_lut6[0] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] svdd sgnd
***** Truth Table for LUT[0], size=6. *****
***** SRAM bits for LUT[0], size=6, num_sram=64. *****
*****0000000000000000000000000000000000000000000000000000000000000000*****
Xsram[0] sram->in sram[0]->out sram[0]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[0]->out) 0
.nodeset V(sram[0]->outb) vsp
Xsram[1] sram->in sram[1]->out sram[1]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[1]->out) 0
.nodeset V(sram[1]->outb) vsp
Xsram[2] sram->in sram[2]->out sram[2]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[2]->out) 0
.nodeset V(sram[2]->outb) vsp
Xsram[3] sram->in sram[3]->out sram[3]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[3]->out) 0
.nodeset V(sram[3]->outb) vsp
Xsram[4] sram->in sram[4]->out sram[4]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[4]->out) 0
.nodeset V(sram[4]->outb) vsp
Xsram[5] sram->in sram[5]->out sram[5]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[5]->out) 0
.nodeset V(sram[5]->outb) vsp
Xsram[6] sram->in sram[6]->out sram[6]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[6]->out) 0
.nodeset V(sram[6]->outb) vsp
Xsram[7] sram->in sram[7]->out sram[7]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[7]->out) 0
.nodeset V(sram[7]->outb) vsp
Xsram[8] sram->in sram[8]->out sram[8]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[8]->out) 0
.nodeset V(sram[8]->outb) vsp
Xsram[9] sram->in sram[9]->out sram[9]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[9]->out) 0
.nodeset V(sram[9]->outb) vsp
Xsram[10] sram->in sram[10]->out sram[10]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[10]->out) 0
.nodeset V(sram[10]->outb) vsp
Xsram[11] sram->in sram[11]->out sram[11]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[11]->out) 0
.nodeset V(sram[11]->outb) vsp
Xsram[12] sram->in sram[12]->out sram[12]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[12]->out) 0
.nodeset V(sram[12]->outb) vsp
Xsram[13] sram->in sram[13]->out sram[13]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[13]->out) 0
.nodeset V(sram[13]->outb) vsp
Xsram[14] sram->in sram[14]->out sram[14]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[14]->out) 0
.nodeset V(sram[14]->outb) vsp
Xsram[15] sram->in sram[15]->out sram[15]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[15]->out) 0
.nodeset V(sram[15]->outb) vsp
Xsram[16] sram->in sram[16]->out sram[16]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[16]->out) 0
.nodeset V(sram[16]->outb) vsp
Xsram[17] sram->in sram[17]->out sram[17]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[17]->out) 0
.nodeset V(sram[17]->outb) vsp
Xsram[18] sram->in sram[18]->out sram[18]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[18]->out) 0
.nodeset V(sram[18]->outb) vsp
Xsram[19] sram->in sram[19]->out sram[19]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[19]->out) 0
.nodeset V(sram[19]->outb) vsp
Xsram[20] sram->in sram[20]->out sram[20]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[20]->out) 0
.nodeset V(sram[20]->outb) vsp
Xsram[21] sram->in sram[21]->out sram[21]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[21]->out) 0
.nodeset V(sram[21]->outb) vsp
Xsram[22] sram->in sram[22]->out sram[22]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[22]->out) 0
.nodeset V(sram[22]->outb) vsp
Xsram[23] sram->in sram[23]->out sram[23]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[23]->out) 0
.nodeset V(sram[23]->outb) vsp
Xsram[24] sram->in sram[24]->out sram[24]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[24]->out) 0
.nodeset V(sram[24]->outb) vsp
Xsram[25] sram->in sram[25]->out sram[25]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[25]->out) 0
.nodeset V(sram[25]->outb) vsp
Xsram[26] sram->in sram[26]->out sram[26]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[26]->out) 0
.nodeset V(sram[26]->outb) vsp
Xsram[27] sram->in sram[27]->out sram[27]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[27]->out) 0
.nodeset V(sram[27]->outb) vsp
Xsram[28] sram->in sram[28]->out sram[28]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[28]->out) 0
.nodeset V(sram[28]->outb) vsp
Xsram[29] sram->in sram[29]->out sram[29]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[29]->out) 0
.nodeset V(sram[29]->outb) vsp
Xsram[30] sram->in sram[30]->out sram[30]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[30]->out) 0
.nodeset V(sram[30]->outb) vsp
Xsram[31] sram->in sram[31]->out sram[31]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[31]->out) 0
.nodeset V(sram[31]->outb) vsp
Xsram[32] sram->in sram[32]->out sram[32]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[32]->out) 0
.nodeset V(sram[32]->outb) vsp
Xsram[33] sram->in sram[33]->out sram[33]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[33]->out) 0
.nodeset V(sram[33]->outb) vsp
Xsram[34] sram->in sram[34]->out sram[34]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[34]->out) 0
.nodeset V(sram[34]->outb) vsp
Xsram[35] sram->in sram[35]->out sram[35]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[35]->out) 0
.nodeset V(sram[35]->outb) vsp
Xsram[36] sram->in sram[36]->out sram[36]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[36]->out) 0
.nodeset V(sram[36]->outb) vsp
Xsram[37] sram->in sram[37]->out sram[37]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[37]->out) 0
.nodeset V(sram[37]->outb) vsp
Xsram[38] sram->in sram[38]->out sram[38]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[38]->out) 0
.nodeset V(sram[38]->outb) vsp
Xsram[39] sram->in sram[39]->out sram[39]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[39]->out) 0
.nodeset V(sram[39]->outb) vsp
Xsram[40] sram->in sram[40]->out sram[40]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[40]->out) 0
.nodeset V(sram[40]->outb) vsp
Xsram[41] sram->in sram[41]->out sram[41]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[41]->out) 0
.nodeset V(sram[41]->outb) vsp
Xsram[42] sram->in sram[42]->out sram[42]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[42]->out) 0
.nodeset V(sram[42]->outb) vsp
Xsram[43] sram->in sram[43]->out sram[43]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[43]->out) 0
.nodeset V(sram[43]->outb) vsp
Xsram[44] sram->in sram[44]->out sram[44]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[44]->out) 0
.nodeset V(sram[44]->outb) vsp
Xsram[45] sram->in sram[45]->out sram[45]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[45]->out) 0
.nodeset V(sram[45]->outb) vsp
Xsram[46] sram->in sram[46]->out sram[46]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[46]->out) 0
.nodeset V(sram[46]->outb) vsp
Xsram[47] sram->in sram[47]->out sram[47]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[47]->out) 0
.nodeset V(sram[47]->outb) vsp
Xsram[48] sram->in sram[48]->out sram[48]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[48]->out) 0
.nodeset V(sram[48]->outb) vsp
Xsram[49] sram->in sram[49]->out sram[49]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[49]->out) 0
.nodeset V(sram[49]->outb) vsp
Xsram[50] sram->in sram[50]->out sram[50]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[50]->out) 0
.nodeset V(sram[50]->outb) vsp
Xsram[51] sram->in sram[51]->out sram[51]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[51]->out) 0
.nodeset V(sram[51]->outb) vsp
Xsram[52] sram->in sram[52]->out sram[52]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[52]->out) 0
.nodeset V(sram[52]->outb) vsp
Xsram[53] sram->in sram[53]->out sram[53]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[53]->out) 0
.nodeset V(sram[53]->outb) vsp
Xsram[54] sram->in sram[54]->out sram[54]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[54]->out) 0
.nodeset V(sram[54]->outb) vsp
Xsram[55] sram->in sram[55]->out sram[55]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[55]->out) 0
.nodeset V(sram[55]->outb) vsp
Xsram[56] sram->in sram[56]->out sram[56]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[56]->out) 0
.nodeset V(sram[56]->outb) vsp
Xsram[57] sram->in sram[57]->out sram[57]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[57]->out) 0
.nodeset V(sram[57]->outb) vsp
Xsram[58] sram->in sram[58]->out sram[58]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[58]->out) 0
.nodeset V(sram[58]->outb) vsp
Xsram[59] sram->in sram[59]->out sram[59]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[59]->out) 0
.nodeset V(sram[59]->outb) vsp
Xsram[60] sram->in sram[60]->out sram[60]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[60]->out) 0
.nodeset V(sram[60]->outb) vsp
Xsram[61] sram->in sram[61]->out sram[61]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[61]->out) 0
.nodeset V(sram[61]->outb) vsp
Xsram[62] sram->in sram[62]->out sram[62]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[62]->out) 0
.nodeset V(sram[62]->outb) vsp
Xsram[63] sram->in sram[63]->out sram[63]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[63]->out) 0
.nodeset V(sram[63]->outb) vsp
Xlut6[0] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] sram[0]->out sram[1]->out sram[2]->out sram[3]->out sram[4]->out sram[5]->out sram[6]->out sram[7]->out sram[8]->out sram[9]->out sram[10]->out sram[11]->out sram[12]->out sram[13]->out sram[14]->out sram[15]->out sram[16]->out sram[17]->out sram[18]->out sram[19]->out sram[20]->out sram[21]->out sram[22]->out sram[23]->out sram[24]->out sram[25]->out sram[26]->out sram[27]->out sram[28]->out sram[29]->out sram[30]->out sram[31]->out sram[32]->out sram[33]->out sram[34]->out sram[35]->out sram[36]->out sram[37]->out sram[38]->out sram[39]->out sram[40]->out sram[41]->out sram[42]->out sram[43]->out sram[44]->out sram[45]->out sram[46]->out sram[47]->out sram[48]->out sram[49]->out sram[50]->out sram[51]->out sram[52]->out sram[53]->out sram[54]->out sram[55]->out sram[56]->out sram[57]->out sram[58]->out sram[59]->out sram[60]->out sram[61]->out sram[62]->out sram[63]->out gvdd_lut6[0] sgnd lut6
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[0]_mode[n1_lut6]_ble6[0]_mode[ble6]_ff[0] ff[0]->D[0] ff[0]->Q[0] svdd sgnd
Xdff[0] 
***** BEGIN Global ports of SPICE_MODEL(static_dff) *****
+  Set[0]  Reset[0]  clk[0] 
***** END Global ports of SPICE_MODEL(static_dff) *****
+ ff[0]->D[0] ff[0]->Q[0] gvdd_dff[0] sgnd static_dff
.nodeset V(ff[0]->Q[0]) 0
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[0]_mode[n1_lut6]_ble6[0]_mode[ble6] mode[ble6]->in[0] mode[ble6]->in[1] mode[ble6]->in[2] mode[ble6]->in[3] mode[ble6]->in[4] mode[ble6]->in[5] mode[ble6]->out[0] mode[ble6]->clk[0] svdd sgnd
Xlut6[0] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[0]_mode[n1_lut6]_ble6[0]_mode[ble6]_lut6[0]
Xff[0] ff[0]->D[0] ff[0]->Q[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[0]_mode[n1_lut6]_ble6[0]_mode[ble6]_ff[0]
Xmux_1level_tapbuf_size2[0] ff[0]->Q[0] lut6[0]->out[0] mode[ble6]->out[0] sram[64]->outb sram[64]->out gvdd_local_interc sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[0], level=1, select_path_id=0. *****
*****1*****
Xsram[64] sram->in sram[64]->out sram[64]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[64]->out) 0
.nodeset V(sram[64]->outb) vsp
Xdirect_interc[0] mode[ble6]->in[0] lut6[0]->in[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[1] mode[ble6]->in[1] lut6[0]->in[1] gvdd_local_interc sgnd direct_interc
Xdirect_interc[2] mode[ble6]->in[2] lut6[0]->in[2] gvdd_local_interc sgnd direct_interc
Xdirect_interc[3] mode[ble6]->in[3] lut6[0]->in[3] gvdd_local_interc sgnd direct_interc
Xdirect_interc[4] mode[ble6]->in[4] lut6[0]->in[4] gvdd_local_interc sgnd direct_interc
Xdirect_interc[5] mode[ble6]->in[5] lut6[0]->in[5] gvdd_local_interc sgnd direct_interc
Xdirect_interc[6] lut6[0]->out[0] ff[0]->D[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[7] mode[ble6]->clk[0] ff[0]->clk[0] gvdd_local_interc sgnd direct_interc
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[0]_mode[n1_lut6] mode[n1_lut6]->in[0] mode[n1_lut6]->in[1] mode[n1_lut6]->in[2] mode[n1_lut6]->in[3] mode[n1_lut6]->in[4] mode[n1_lut6]->in[5] mode[n1_lut6]->out[0] mode[n1_lut6]->clk[0] svdd sgnd
Xble6[0] ble6[0]->in[0] ble6[0]->in[1] ble6[0]->in[2] ble6[0]->in[3] ble6[0]->in[4] ble6[0]->in[5] ble6[0]->out[0] ble6[0]->clk[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[0]_mode[n1_lut6]_ble6[0]_mode[ble6]
Xdirect_interc[8] ble6[0]->out[0] mode[n1_lut6]->out[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[9] mode[n1_lut6]->in[0] ble6[0]->in[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[10] mode[n1_lut6]->in[1] ble6[0]->in[1] gvdd_local_interc sgnd direct_interc
Xdirect_interc[11] mode[n1_lut6]->in[2] ble6[0]->in[2] gvdd_local_interc sgnd direct_interc
Xdirect_interc[12] mode[n1_lut6]->in[3] ble6[0]->in[3] gvdd_local_interc sgnd direct_interc
Xdirect_interc[13] mode[n1_lut6]->in[4] ble6[0]->in[4] gvdd_local_interc sgnd direct_interc
Xdirect_interc[14] mode[n1_lut6]->in[5] ble6[0]->in[5] gvdd_local_interc sgnd direct_interc
Xdirect_interc[15] mode[n1_lut6]->clk[0] ble6[0]->clk[0] gvdd_local_interc sgnd direct_interc
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[1]_mode[n1_lut6]_ble6[0]_mode[ble6]_lut6[0] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] svdd sgnd
***** Truth Table for LUT[1], size=6. *****
***** SRAM bits for LUT[1], size=6, num_sram=64. *****
*****0000000000000000000000000000000000000000000000000000000000000000*****
Xsram[65] sram->in sram[65]->out sram[65]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[65]->out) 0
.nodeset V(sram[65]->outb) vsp
Xsram[66] sram->in sram[66]->out sram[66]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[66]->out) 0
.nodeset V(sram[66]->outb) vsp
Xsram[67] sram->in sram[67]->out sram[67]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[67]->out) 0
.nodeset V(sram[67]->outb) vsp
Xsram[68] sram->in sram[68]->out sram[68]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[68]->out) 0
.nodeset V(sram[68]->outb) vsp
Xsram[69] sram->in sram[69]->out sram[69]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[69]->out) 0
.nodeset V(sram[69]->outb) vsp
Xsram[70] sram->in sram[70]->out sram[70]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[70]->out) 0
.nodeset V(sram[70]->outb) vsp
Xsram[71] sram->in sram[71]->out sram[71]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[71]->out) 0
.nodeset V(sram[71]->outb) vsp
Xsram[72] sram->in sram[72]->out sram[72]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[72]->out) 0
.nodeset V(sram[72]->outb) vsp
Xsram[73] sram->in sram[73]->out sram[73]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[73]->out) 0
.nodeset V(sram[73]->outb) vsp
Xsram[74] sram->in sram[74]->out sram[74]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[74]->out) 0
.nodeset V(sram[74]->outb) vsp
Xsram[75] sram->in sram[75]->out sram[75]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[75]->out) 0
.nodeset V(sram[75]->outb) vsp
Xsram[76] sram->in sram[76]->out sram[76]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[76]->out) 0
.nodeset V(sram[76]->outb) vsp
Xsram[77] sram->in sram[77]->out sram[77]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[77]->out) 0
.nodeset V(sram[77]->outb) vsp
Xsram[78] sram->in sram[78]->out sram[78]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[78]->out) 0
.nodeset V(sram[78]->outb) vsp
Xsram[79] sram->in sram[79]->out sram[79]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[79]->out) 0
.nodeset V(sram[79]->outb) vsp
Xsram[80] sram->in sram[80]->out sram[80]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[80]->out) 0
.nodeset V(sram[80]->outb) vsp
Xsram[81] sram->in sram[81]->out sram[81]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[81]->out) 0
.nodeset V(sram[81]->outb) vsp
Xsram[82] sram->in sram[82]->out sram[82]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[82]->out) 0
.nodeset V(sram[82]->outb) vsp
Xsram[83] sram->in sram[83]->out sram[83]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[83]->out) 0
.nodeset V(sram[83]->outb) vsp
Xsram[84] sram->in sram[84]->out sram[84]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[84]->out) 0
.nodeset V(sram[84]->outb) vsp
Xsram[85] sram->in sram[85]->out sram[85]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[85]->out) 0
.nodeset V(sram[85]->outb) vsp
Xsram[86] sram->in sram[86]->out sram[86]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[86]->out) 0
.nodeset V(sram[86]->outb) vsp
Xsram[87] sram->in sram[87]->out sram[87]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[87]->out) 0
.nodeset V(sram[87]->outb) vsp
Xsram[88] sram->in sram[88]->out sram[88]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[88]->out) 0
.nodeset V(sram[88]->outb) vsp
Xsram[89] sram->in sram[89]->out sram[89]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[89]->out) 0
.nodeset V(sram[89]->outb) vsp
Xsram[90] sram->in sram[90]->out sram[90]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[90]->out) 0
.nodeset V(sram[90]->outb) vsp
Xsram[91] sram->in sram[91]->out sram[91]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[91]->out) 0
.nodeset V(sram[91]->outb) vsp
Xsram[92] sram->in sram[92]->out sram[92]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[92]->out) 0
.nodeset V(sram[92]->outb) vsp
Xsram[93] sram->in sram[93]->out sram[93]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[93]->out) 0
.nodeset V(sram[93]->outb) vsp
Xsram[94] sram->in sram[94]->out sram[94]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[94]->out) 0
.nodeset V(sram[94]->outb) vsp
Xsram[95] sram->in sram[95]->out sram[95]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[95]->out) 0
.nodeset V(sram[95]->outb) vsp
Xsram[96] sram->in sram[96]->out sram[96]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[96]->out) 0
.nodeset V(sram[96]->outb) vsp
Xsram[97] sram->in sram[97]->out sram[97]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[97]->out) 0
.nodeset V(sram[97]->outb) vsp
Xsram[98] sram->in sram[98]->out sram[98]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[98]->out) 0
.nodeset V(sram[98]->outb) vsp
Xsram[99] sram->in sram[99]->out sram[99]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[99]->out) 0
.nodeset V(sram[99]->outb) vsp
Xsram[100] sram->in sram[100]->out sram[100]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[100]->out) 0
.nodeset V(sram[100]->outb) vsp
Xsram[101] sram->in sram[101]->out sram[101]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[101]->out) 0
.nodeset V(sram[101]->outb) vsp
Xsram[102] sram->in sram[102]->out sram[102]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[102]->out) 0
.nodeset V(sram[102]->outb) vsp
Xsram[103] sram->in sram[103]->out sram[103]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[103]->out) 0
.nodeset V(sram[103]->outb) vsp
Xsram[104] sram->in sram[104]->out sram[104]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[104]->out) 0
.nodeset V(sram[104]->outb) vsp
Xsram[105] sram->in sram[105]->out sram[105]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[105]->out) 0
.nodeset V(sram[105]->outb) vsp
Xsram[106] sram->in sram[106]->out sram[106]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[106]->out) 0
.nodeset V(sram[106]->outb) vsp
Xsram[107] sram->in sram[107]->out sram[107]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[107]->out) 0
.nodeset V(sram[107]->outb) vsp
Xsram[108] sram->in sram[108]->out sram[108]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[108]->out) 0
.nodeset V(sram[108]->outb) vsp
Xsram[109] sram->in sram[109]->out sram[109]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[109]->out) 0
.nodeset V(sram[109]->outb) vsp
Xsram[110] sram->in sram[110]->out sram[110]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[110]->out) 0
.nodeset V(sram[110]->outb) vsp
Xsram[111] sram->in sram[111]->out sram[111]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[111]->out) 0
.nodeset V(sram[111]->outb) vsp
Xsram[112] sram->in sram[112]->out sram[112]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[112]->out) 0
.nodeset V(sram[112]->outb) vsp
Xsram[113] sram->in sram[113]->out sram[113]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[113]->out) 0
.nodeset V(sram[113]->outb) vsp
Xsram[114] sram->in sram[114]->out sram[114]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[114]->out) 0
.nodeset V(sram[114]->outb) vsp
Xsram[115] sram->in sram[115]->out sram[115]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[115]->out) 0
.nodeset V(sram[115]->outb) vsp
Xsram[116] sram->in sram[116]->out sram[116]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[116]->out) 0
.nodeset V(sram[116]->outb) vsp
Xsram[117] sram->in sram[117]->out sram[117]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[117]->out) 0
.nodeset V(sram[117]->outb) vsp
Xsram[118] sram->in sram[118]->out sram[118]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[118]->out) 0
.nodeset V(sram[118]->outb) vsp
Xsram[119] sram->in sram[119]->out sram[119]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[119]->out) 0
.nodeset V(sram[119]->outb) vsp
Xsram[120] sram->in sram[120]->out sram[120]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[120]->out) 0
.nodeset V(sram[120]->outb) vsp
Xsram[121] sram->in sram[121]->out sram[121]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[121]->out) 0
.nodeset V(sram[121]->outb) vsp
Xsram[122] sram->in sram[122]->out sram[122]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[122]->out) 0
.nodeset V(sram[122]->outb) vsp
Xsram[123] sram->in sram[123]->out sram[123]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[123]->out) 0
.nodeset V(sram[123]->outb) vsp
Xsram[124] sram->in sram[124]->out sram[124]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[124]->out) 0
.nodeset V(sram[124]->outb) vsp
Xsram[125] sram->in sram[125]->out sram[125]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[125]->out) 0
.nodeset V(sram[125]->outb) vsp
Xsram[126] sram->in sram[126]->out sram[126]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[126]->out) 0
.nodeset V(sram[126]->outb) vsp
Xsram[127] sram->in sram[127]->out sram[127]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[127]->out) 0
.nodeset V(sram[127]->outb) vsp
Xsram[128] sram->in sram[128]->out sram[128]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[128]->out) 0
.nodeset V(sram[128]->outb) vsp
Xlut6[1] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] sram[65]->out sram[66]->out sram[67]->out sram[68]->out sram[69]->out sram[70]->out sram[71]->out sram[72]->out sram[73]->out sram[74]->out sram[75]->out sram[76]->out sram[77]->out sram[78]->out sram[79]->out sram[80]->out sram[81]->out sram[82]->out sram[83]->out sram[84]->out sram[85]->out sram[86]->out sram[87]->out sram[88]->out sram[89]->out sram[90]->out sram[91]->out sram[92]->out sram[93]->out sram[94]->out sram[95]->out sram[96]->out sram[97]->out sram[98]->out sram[99]->out sram[100]->out sram[101]->out sram[102]->out sram[103]->out sram[104]->out sram[105]->out sram[106]->out sram[107]->out sram[108]->out sram[109]->out sram[110]->out sram[111]->out sram[112]->out sram[113]->out sram[114]->out sram[115]->out sram[116]->out sram[117]->out sram[118]->out sram[119]->out sram[120]->out sram[121]->out sram[122]->out sram[123]->out sram[124]->out sram[125]->out sram[126]->out sram[127]->out sram[128]->out gvdd_lut6[1] sgnd lut6
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[1]_mode[n1_lut6]_ble6[0]_mode[ble6]_ff[0] ff[0]->D[0] ff[0]->Q[0] svdd sgnd
Xdff[1] 
***** BEGIN Global ports of SPICE_MODEL(static_dff) *****
+  Set[0]  Reset[0]  clk[0] 
***** END Global ports of SPICE_MODEL(static_dff) *****
+ ff[0]->D[0] ff[0]->Q[0] gvdd_dff[1] sgnd static_dff
.nodeset V(ff[0]->Q[0]) 0
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[1]_mode[n1_lut6]_ble6[0]_mode[ble6] mode[ble6]->in[0] mode[ble6]->in[1] mode[ble6]->in[2] mode[ble6]->in[3] mode[ble6]->in[4] mode[ble6]->in[5] mode[ble6]->out[0] mode[ble6]->clk[0] svdd sgnd
Xlut6[0] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[1]_mode[n1_lut6]_ble6[0]_mode[ble6]_lut6[0]
Xff[0] ff[0]->D[0] ff[0]->Q[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[1]_mode[n1_lut6]_ble6[0]_mode[ble6]_ff[0]
Xmux_1level_tapbuf_size2[1] ff[0]->Q[0] lut6[0]->out[0] mode[ble6]->out[0] sram[129]->outb sram[129]->out gvdd_local_interc sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[1], level=1, select_path_id=0. *****
*****1*****
Xsram[129] sram->in sram[129]->out sram[129]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[129]->out) 0
.nodeset V(sram[129]->outb) vsp
Xdirect_interc[16] mode[ble6]->in[0] lut6[0]->in[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[17] mode[ble6]->in[1] lut6[0]->in[1] gvdd_local_interc sgnd direct_interc
Xdirect_interc[18] mode[ble6]->in[2] lut6[0]->in[2] gvdd_local_interc sgnd direct_interc
Xdirect_interc[19] mode[ble6]->in[3] lut6[0]->in[3] gvdd_local_interc sgnd direct_interc
Xdirect_interc[20] mode[ble6]->in[4] lut6[0]->in[4] gvdd_local_interc sgnd direct_interc
Xdirect_interc[21] mode[ble6]->in[5] lut6[0]->in[5] gvdd_local_interc sgnd direct_interc
Xdirect_interc[22] lut6[0]->out[0] ff[0]->D[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[23] mode[ble6]->clk[0] ff[0]->clk[0] gvdd_local_interc sgnd direct_interc
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[1]_mode[n1_lut6] mode[n1_lut6]->in[0] mode[n1_lut6]->in[1] mode[n1_lut6]->in[2] mode[n1_lut6]->in[3] mode[n1_lut6]->in[4] mode[n1_lut6]->in[5] mode[n1_lut6]->out[0] mode[n1_lut6]->clk[0] svdd sgnd
Xble6[0] ble6[0]->in[0] ble6[0]->in[1] ble6[0]->in[2] ble6[0]->in[3] ble6[0]->in[4] ble6[0]->in[5] ble6[0]->out[0] ble6[0]->clk[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[1]_mode[n1_lut6]_ble6[0]_mode[ble6]
Xdirect_interc[24] ble6[0]->out[0] mode[n1_lut6]->out[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[25] mode[n1_lut6]->in[0] ble6[0]->in[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[26] mode[n1_lut6]->in[1] ble6[0]->in[1] gvdd_local_interc sgnd direct_interc
Xdirect_interc[27] mode[n1_lut6]->in[2] ble6[0]->in[2] gvdd_local_interc sgnd direct_interc
Xdirect_interc[28] mode[n1_lut6]->in[3] ble6[0]->in[3] gvdd_local_interc sgnd direct_interc
Xdirect_interc[29] mode[n1_lut6]->in[4] ble6[0]->in[4] gvdd_local_interc sgnd direct_interc
Xdirect_interc[30] mode[n1_lut6]->in[5] ble6[0]->in[5] gvdd_local_interc sgnd direct_interc
Xdirect_interc[31] mode[n1_lut6]->clk[0] ble6[0]->clk[0] gvdd_local_interc sgnd direct_interc
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[2]_mode[n1_lut6]_ble6[0]_mode[ble6]_lut6[0] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] svdd sgnd
***** Truth Table for LUT[2], size=6. *****
***** SRAM bits for LUT[2], size=6, num_sram=64. *****
*****0000000000000000000000000000000000000000000000000000000000000000*****
Xsram[130] sram->in sram[130]->out sram[130]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[130]->out) 0
.nodeset V(sram[130]->outb) vsp
Xsram[131] sram->in sram[131]->out sram[131]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[131]->out) 0
.nodeset V(sram[131]->outb) vsp
Xsram[132] sram->in sram[132]->out sram[132]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[132]->out) 0
.nodeset V(sram[132]->outb) vsp
Xsram[133] sram->in sram[133]->out sram[133]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[133]->out) 0
.nodeset V(sram[133]->outb) vsp
Xsram[134] sram->in sram[134]->out sram[134]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[134]->out) 0
.nodeset V(sram[134]->outb) vsp
Xsram[135] sram->in sram[135]->out sram[135]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[135]->out) 0
.nodeset V(sram[135]->outb) vsp
Xsram[136] sram->in sram[136]->out sram[136]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[136]->out) 0
.nodeset V(sram[136]->outb) vsp
Xsram[137] sram->in sram[137]->out sram[137]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[137]->out) 0
.nodeset V(sram[137]->outb) vsp
Xsram[138] sram->in sram[138]->out sram[138]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[138]->out) 0
.nodeset V(sram[138]->outb) vsp
Xsram[139] sram->in sram[139]->out sram[139]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[139]->out) 0
.nodeset V(sram[139]->outb) vsp
Xsram[140] sram->in sram[140]->out sram[140]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[140]->out) 0
.nodeset V(sram[140]->outb) vsp
Xsram[141] sram->in sram[141]->out sram[141]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[141]->out) 0
.nodeset V(sram[141]->outb) vsp
Xsram[142] sram->in sram[142]->out sram[142]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[142]->out) 0
.nodeset V(sram[142]->outb) vsp
Xsram[143] sram->in sram[143]->out sram[143]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[143]->out) 0
.nodeset V(sram[143]->outb) vsp
Xsram[144] sram->in sram[144]->out sram[144]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[144]->out) 0
.nodeset V(sram[144]->outb) vsp
Xsram[145] sram->in sram[145]->out sram[145]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[145]->out) 0
.nodeset V(sram[145]->outb) vsp
Xsram[146] sram->in sram[146]->out sram[146]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[146]->out) 0
.nodeset V(sram[146]->outb) vsp
Xsram[147] sram->in sram[147]->out sram[147]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[147]->out) 0
.nodeset V(sram[147]->outb) vsp
Xsram[148] sram->in sram[148]->out sram[148]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[148]->out) 0
.nodeset V(sram[148]->outb) vsp
Xsram[149] sram->in sram[149]->out sram[149]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[149]->out) 0
.nodeset V(sram[149]->outb) vsp
Xsram[150] sram->in sram[150]->out sram[150]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[150]->out) 0
.nodeset V(sram[150]->outb) vsp
Xsram[151] sram->in sram[151]->out sram[151]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[151]->out) 0
.nodeset V(sram[151]->outb) vsp
Xsram[152] sram->in sram[152]->out sram[152]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[152]->out) 0
.nodeset V(sram[152]->outb) vsp
Xsram[153] sram->in sram[153]->out sram[153]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[153]->out) 0
.nodeset V(sram[153]->outb) vsp
Xsram[154] sram->in sram[154]->out sram[154]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[154]->out) 0
.nodeset V(sram[154]->outb) vsp
Xsram[155] sram->in sram[155]->out sram[155]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[155]->out) 0
.nodeset V(sram[155]->outb) vsp
Xsram[156] sram->in sram[156]->out sram[156]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[156]->out) 0
.nodeset V(sram[156]->outb) vsp
Xsram[157] sram->in sram[157]->out sram[157]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[157]->out) 0
.nodeset V(sram[157]->outb) vsp
Xsram[158] sram->in sram[158]->out sram[158]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[158]->out) 0
.nodeset V(sram[158]->outb) vsp
Xsram[159] sram->in sram[159]->out sram[159]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[159]->out) 0
.nodeset V(sram[159]->outb) vsp
Xsram[160] sram->in sram[160]->out sram[160]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[160]->out) 0
.nodeset V(sram[160]->outb) vsp
Xsram[161] sram->in sram[161]->out sram[161]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[161]->out) 0
.nodeset V(sram[161]->outb) vsp
Xsram[162] sram->in sram[162]->out sram[162]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[162]->out) 0
.nodeset V(sram[162]->outb) vsp
Xsram[163] sram->in sram[163]->out sram[163]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[163]->out) 0
.nodeset V(sram[163]->outb) vsp
Xsram[164] sram->in sram[164]->out sram[164]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[164]->out) 0
.nodeset V(sram[164]->outb) vsp
Xsram[165] sram->in sram[165]->out sram[165]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[165]->out) 0
.nodeset V(sram[165]->outb) vsp
Xsram[166] sram->in sram[166]->out sram[166]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[166]->out) 0
.nodeset V(sram[166]->outb) vsp
Xsram[167] sram->in sram[167]->out sram[167]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[167]->out) 0
.nodeset V(sram[167]->outb) vsp
Xsram[168] sram->in sram[168]->out sram[168]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[168]->out) 0
.nodeset V(sram[168]->outb) vsp
Xsram[169] sram->in sram[169]->out sram[169]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[169]->out) 0
.nodeset V(sram[169]->outb) vsp
Xsram[170] sram->in sram[170]->out sram[170]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[170]->out) 0
.nodeset V(sram[170]->outb) vsp
Xsram[171] sram->in sram[171]->out sram[171]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[171]->out) 0
.nodeset V(sram[171]->outb) vsp
Xsram[172] sram->in sram[172]->out sram[172]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[172]->out) 0
.nodeset V(sram[172]->outb) vsp
Xsram[173] sram->in sram[173]->out sram[173]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[173]->out) 0
.nodeset V(sram[173]->outb) vsp
Xsram[174] sram->in sram[174]->out sram[174]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[174]->out) 0
.nodeset V(sram[174]->outb) vsp
Xsram[175] sram->in sram[175]->out sram[175]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[175]->out) 0
.nodeset V(sram[175]->outb) vsp
Xsram[176] sram->in sram[176]->out sram[176]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[176]->out) 0
.nodeset V(sram[176]->outb) vsp
Xsram[177] sram->in sram[177]->out sram[177]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[177]->out) 0
.nodeset V(sram[177]->outb) vsp
Xsram[178] sram->in sram[178]->out sram[178]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[178]->out) 0
.nodeset V(sram[178]->outb) vsp
Xsram[179] sram->in sram[179]->out sram[179]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[179]->out) 0
.nodeset V(sram[179]->outb) vsp
Xsram[180] sram->in sram[180]->out sram[180]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[180]->out) 0
.nodeset V(sram[180]->outb) vsp
Xsram[181] sram->in sram[181]->out sram[181]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[181]->out) 0
.nodeset V(sram[181]->outb) vsp
Xsram[182] sram->in sram[182]->out sram[182]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[182]->out) 0
.nodeset V(sram[182]->outb) vsp
Xsram[183] sram->in sram[183]->out sram[183]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[183]->out) 0
.nodeset V(sram[183]->outb) vsp
Xsram[184] sram->in sram[184]->out sram[184]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[184]->out) 0
.nodeset V(sram[184]->outb) vsp
Xsram[185] sram->in sram[185]->out sram[185]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[185]->out) 0
.nodeset V(sram[185]->outb) vsp
Xsram[186] sram->in sram[186]->out sram[186]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[186]->out) 0
.nodeset V(sram[186]->outb) vsp
Xsram[187] sram->in sram[187]->out sram[187]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[187]->out) 0
.nodeset V(sram[187]->outb) vsp
Xsram[188] sram->in sram[188]->out sram[188]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[188]->out) 0
.nodeset V(sram[188]->outb) vsp
Xsram[189] sram->in sram[189]->out sram[189]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[189]->out) 0
.nodeset V(sram[189]->outb) vsp
Xsram[190] sram->in sram[190]->out sram[190]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[190]->out) 0
.nodeset V(sram[190]->outb) vsp
Xsram[191] sram->in sram[191]->out sram[191]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[191]->out) 0
.nodeset V(sram[191]->outb) vsp
Xsram[192] sram->in sram[192]->out sram[192]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[192]->out) 0
.nodeset V(sram[192]->outb) vsp
Xsram[193] sram->in sram[193]->out sram[193]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[193]->out) 0
.nodeset V(sram[193]->outb) vsp
Xlut6[2] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] sram[130]->out sram[131]->out sram[132]->out sram[133]->out sram[134]->out sram[135]->out sram[136]->out sram[137]->out sram[138]->out sram[139]->out sram[140]->out sram[141]->out sram[142]->out sram[143]->out sram[144]->out sram[145]->out sram[146]->out sram[147]->out sram[148]->out sram[149]->out sram[150]->out sram[151]->out sram[152]->out sram[153]->out sram[154]->out sram[155]->out sram[156]->out sram[157]->out sram[158]->out sram[159]->out sram[160]->out sram[161]->out sram[162]->out sram[163]->out sram[164]->out sram[165]->out sram[166]->out sram[167]->out sram[168]->out sram[169]->out sram[170]->out sram[171]->out sram[172]->out sram[173]->out sram[174]->out sram[175]->out sram[176]->out sram[177]->out sram[178]->out sram[179]->out sram[180]->out sram[181]->out sram[182]->out sram[183]->out sram[184]->out sram[185]->out sram[186]->out sram[187]->out sram[188]->out sram[189]->out sram[190]->out sram[191]->out sram[192]->out sram[193]->out gvdd_lut6[2] sgnd lut6
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[2]_mode[n1_lut6]_ble6[0]_mode[ble6]_ff[0] ff[0]->D[0] ff[0]->Q[0] svdd sgnd
Xdff[2] 
***** BEGIN Global ports of SPICE_MODEL(static_dff) *****
+  Set[0]  Reset[0]  clk[0] 
***** END Global ports of SPICE_MODEL(static_dff) *****
+ ff[0]->D[0] ff[0]->Q[0] gvdd_dff[2] sgnd static_dff
.nodeset V(ff[0]->Q[0]) 0
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[2]_mode[n1_lut6]_ble6[0]_mode[ble6] mode[ble6]->in[0] mode[ble6]->in[1] mode[ble6]->in[2] mode[ble6]->in[3] mode[ble6]->in[4] mode[ble6]->in[5] mode[ble6]->out[0] mode[ble6]->clk[0] svdd sgnd
Xlut6[0] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[2]_mode[n1_lut6]_ble6[0]_mode[ble6]_lut6[0]
Xff[0] ff[0]->D[0] ff[0]->Q[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[2]_mode[n1_lut6]_ble6[0]_mode[ble6]_ff[0]
Xmux_1level_tapbuf_size2[2] ff[0]->Q[0] lut6[0]->out[0] mode[ble6]->out[0] sram[194]->outb sram[194]->out gvdd_local_interc sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[2], level=1, select_path_id=0. *****
*****1*****
Xsram[194] sram->in sram[194]->out sram[194]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[194]->out) 0
.nodeset V(sram[194]->outb) vsp
Xdirect_interc[32] mode[ble6]->in[0] lut6[0]->in[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[33] mode[ble6]->in[1] lut6[0]->in[1] gvdd_local_interc sgnd direct_interc
Xdirect_interc[34] mode[ble6]->in[2] lut6[0]->in[2] gvdd_local_interc sgnd direct_interc
Xdirect_interc[35] mode[ble6]->in[3] lut6[0]->in[3] gvdd_local_interc sgnd direct_interc
Xdirect_interc[36] mode[ble6]->in[4] lut6[0]->in[4] gvdd_local_interc sgnd direct_interc
Xdirect_interc[37] mode[ble6]->in[5] lut6[0]->in[5] gvdd_local_interc sgnd direct_interc
Xdirect_interc[38] lut6[0]->out[0] ff[0]->D[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[39] mode[ble6]->clk[0] ff[0]->clk[0] gvdd_local_interc sgnd direct_interc
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[2]_mode[n1_lut6] mode[n1_lut6]->in[0] mode[n1_lut6]->in[1] mode[n1_lut6]->in[2] mode[n1_lut6]->in[3] mode[n1_lut6]->in[4] mode[n1_lut6]->in[5] mode[n1_lut6]->out[0] mode[n1_lut6]->clk[0] svdd sgnd
Xble6[0] ble6[0]->in[0] ble6[0]->in[1] ble6[0]->in[2] ble6[0]->in[3] ble6[0]->in[4] ble6[0]->in[5] ble6[0]->out[0] ble6[0]->clk[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[2]_mode[n1_lut6]_ble6[0]_mode[ble6]
Xdirect_interc[40] ble6[0]->out[0] mode[n1_lut6]->out[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[41] mode[n1_lut6]->in[0] ble6[0]->in[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[42] mode[n1_lut6]->in[1] ble6[0]->in[1] gvdd_local_interc sgnd direct_interc
Xdirect_interc[43] mode[n1_lut6]->in[2] ble6[0]->in[2] gvdd_local_interc sgnd direct_interc
Xdirect_interc[44] mode[n1_lut6]->in[3] ble6[0]->in[3] gvdd_local_interc sgnd direct_interc
Xdirect_interc[45] mode[n1_lut6]->in[4] ble6[0]->in[4] gvdd_local_interc sgnd direct_interc
Xdirect_interc[46] mode[n1_lut6]->in[5] ble6[0]->in[5] gvdd_local_interc sgnd direct_interc
Xdirect_interc[47] mode[n1_lut6]->clk[0] ble6[0]->clk[0] gvdd_local_interc sgnd direct_interc
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[3]_mode[n1_lut6]_ble6[0]_mode[ble6]_lut6[0] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] svdd sgnd
***** Truth Table for LUT[3], size=6. *****
***** SRAM bits for LUT[3], size=6, num_sram=64. *****
*****0000000000000000000000000000000000000000000000000000000000000000*****
Xsram[195] sram->in sram[195]->out sram[195]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[195]->out) 0
.nodeset V(sram[195]->outb) vsp
Xsram[196] sram->in sram[196]->out sram[196]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[196]->out) 0
.nodeset V(sram[196]->outb) vsp
Xsram[197] sram->in sram[197]->out sram[197]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[197]->out) 0
.nodeset V(sram[197]->outb) vsp
Xsram[198] sram->in sram[198]->out sram[198]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[198]->out) 0
.nodeset V(sram[198]->outb) vsp
Xsram[199] sram->in sram[199]->out sram[199]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[199]->out) 0
.nodeset V(sram[199]->outb) vsp
Xsram[200] sram->in sram[200]->out sram[200]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[200]->out) 0
.nodeset V(sram[200]->outb) vsp
Xsram[201] sram->in sram[201]->out sram[201]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[201]->out) 0
.nodeset V(sram[201]->outb) vsp
Xsram[202] sram->in sram[202]->out sram[202]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[202]->out) 0
.nodeset V(sram[202]->outb) vsp
Xsram[203] sram->in sram[203]->out sram[203]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[203]->out) 0
.nodeset V(sram[203]->outb) vsp
Xsram[204] sram->in sram[204]->out sram[204]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[204]->out) 0
.nodeset V(sram[204]->outb) vsp
Xsram[205] sram->in sram[205]->out sram[205]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[205]->out) 0
.nodeset V(sram[205]->outb) vsp
Xsram[206] sram->in sram[206]->out sram[206]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[206]->out) 0
.nodeset V(sram[206]->outb) vsp
Xsram[207] sram->in sram[207]->out sram[207]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[207]->out) 0
.nodeset V(sram[207]->outb) vsp
Xsram[208] sram->in sram[208]->out sram[208]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[208]->out) 0
.nodeset V(sram[208]->outb) vsp
Xsram[209] sram->in sram[209]->out sram[209]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[209]->out) 0
.nodeset V(sram[209]->outb) vsp
Xsram[210] sram->in sram[210]->out sram[210]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[210]->out) 0
.nodeset V(sram[210]->outb) vsp
Xsram[211] sram->in sram[211]->out sram[211]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[211]->out) 0
.nodeset V(sram[211]->outb) vsp
Xsram[212] sram->in sram[212]->out sram[212]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[212]->out) 0
.nodeset V(sram[212]->outb) vsp
Xsram[213] sram->in sram[213]->out sram[213]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[213]->out) 0
.nodeset V(sram[213]->outb) vsp
Xsram[214] sram->in sram[214]->out sram[214]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[214]->out) 0
.nodeset V(sram[214]->outb) vsp
Xsram[215] sram->in sram[215]->out sram[215]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[215]->out) 0
.nodeset V(sram[215]->outb) vsp
Xsram[216] sram->in sram[216]->out sram[216]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[216]->out) 0
.nodeset V(sram[216]->outb) vsp
Xsram[217] sram->in sram[217]->out sram[217]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[217]->out) 0
.nodeset V(sram[217]->outb) vsp
Xsram[218] sram->in sram[218]->out sram[218]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[218]->out) 0
.nodeset V(sram[218]->outb) vsp
Xsram[219] sram->in sram[219]->out sram[219]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[219]->out) 0
.nodeset V(sram[219]->outb) vsp
Xsram[220] sram->in sram[220]->out sram[220]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[220]->out) 0
.nodeset V(sram[220]->outb) vsp
Xsram[221] sram->in sram[221]->out sram[221]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[221]->out) 0
.nodeset V(sram[221]->outb) vsp
Xsram[222] sram->in sram[222]->out sram[222]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[222]->out) 0
.nodeset V(sram[222]->outb) vsp
Xsram[223] sram->in sram[223]->out sram[223]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[223]->out) 0
.nodeset V(sram[223]->outb) vsp
Xsram[224] sram->in sram[224]->out sram[224]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[224]->out) 0
.nodeset V(sram[224]->outb) vsp
Xsram[225] sram->in sram[225]->out sram[225]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[225]->out) 0
.nodeset V(sram[225]->outb) vsp
Xsram[226] sram->in sram[226]->out sram[226]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[226]->out) 0
.nodeset V(sram[226]->outb) vsp
Xsram[227] sram->in sram[227]->out sram[227]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[227]->out) 0
.nodeset V(sram[227]->outb) vsp
Xsram[228] sram->in sram[228]->out sram[228]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[228]->out) 0
.nodeset V(sram[228]->outb) vsp
Xsram[229] sram->in sram[229]->out sram[229]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[229]->out) 0
.nodeset V(sram[229]->outb) vsp
Xsram[230] sram->in sram[230]->out sram[230]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[230]->out) 0
.nodeset V(sram[230]->outb) vsp
Xsram[231] sram->in sram[231]->out sram[231]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[231]->out) 0
.nodeset V(sram[231]->outb) vsp
Xsram[232] sram->in sram[232]->out sram[232]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[232]->out) 0
.nodeset V(sram[232]->outb) vsp
Xsram[233] sram->in sram[233]->out sram[233]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[233]->out) 0
.nodeset V(sram[233]->outb) vsp
Xsram[234] sram->in sram[234]->out sram[234]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[234]->out) 0
.nodeset V(sram[234]->outb) vsp
Xsram[235] sram->in sram[235]->out sram[235]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[235]->out) 0
.nodeset V(sram[235]->outb) vsp
Xsram[236] sram->in sram[236]->out sram[236]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[236]->out) 0
.nodeset V(sram[236]->outb) vsp
Xsram[237] sram->in sram[237]->out sram[237]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[237]->out) 0
.nodeset V(sram[237]->outb) vsp
Xsram[238] sram->in sram[238]->out sram[238]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[238]->out) 0
.nodeset V(sram[238]->outb) vsp
Xsram[239] sram->in sram[239]->out sram[239]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[239]->out) 0
.nodeset V(sram[239]->outb) vsp
Xsram[240] sram->in sram[240]->out sram[240]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[240]->out) 0
.nodeset V(sram[240]->outb) vsp
Xsram[241] sram->in sram[241]->out sram[241]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[241]->out) 0
.nodeset V(sram[241]->outb) vsp
Xsram[242] sram->in sram[242]->out sram[242]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[242]->out) 0
.nodeset V(sram[242]->outb) vsp
Xsram[243] sram->in sram[243]->out sram[243]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[243]->out) 0
.nodeset V(sram[243]->outb) vsp
Xsram[244] sram->in sram[244]->out sram[244]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[244]->out) 0
.nodeset V(sram[244]->outb) vsp
Xsram[245] sram->in sram[245]->out sram[245]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[245]->out) 0
.nodeset V(sram[245]->outb) vsp
Xsram[246] sram->in sram[246]->out sram[246]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[246]->out) 0
.nodeset V(sram[246]->outb) vsp
Xsram[247] sram->in sram[247]->out sram[247]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[247]->out) 0
.nodeset V(sram[247]->outb) vsp
Xsram[248] sram->in sram[248]->out sram[248]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[248]->out) 0
.nodeset V(sram[248]->outb) vsp
Xsram[249] sram->in sram[249]->out sram[249]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[249]->out) 0
.nodeset V(sram[249]->outb) vsp
Xsram[250] sram->in sram[250]->out sram[250]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[250]->out) 0
.nodeset V(sram[250]->outb) vsp
Xsram[251] sram->in sram[251]->out sram[251]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[251]->out) 0
.nodeset V(sram[251]->outb) vsp
Xsram[252] sram->in sram[252]->out sram[252]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[252]->out) 0
.nodeset V(sram[252]->outb) vsp
Xsram[253] sram->in sram[253]->out sram[253]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[253]->out) 0
.nodeset V(sram[253]->outb) vsp
Xsram[254] sram->in sram[254]->out sram[254]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[254]->out) 0
.nodeset V(sram[254]->outb) vsp
Xsram[255] sram->in sram[255]->out sram[255]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[255]->out) 0
.nodeset V(sram[255]->outb) vsp
Xsram[256] sram->in sram[256]->out sram[256]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[256]->out) 0
.nodeset V(sram[256]->outb) vsp
Xsram[257] sram->in sram[257]->out sram[257]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[257]->out) 0
.nodeset V(sram[257]->outb) vsp
Xsram[258] sram->in sram[258]->out sram[258]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[258]->out) 0
.nodeset V(sram[258]->outb) vsp
Xlut6[3] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] sram[195]->out sram[196]->out sram[197]->out sram[198]->out sram[199]->out sram[200]->out sram[201]->out sram[202]->out sram[203]->out sram[204]->out sram[205]->out sram[206]->out sram[207]->out sram[208]->out sram[209]->out sram[210]->out sram[211]->out sram[212]->out sram[213]->out sram[214]->out sram[215]->out sram[216]->out sram[217]->out sram[218]->out sram[219]->out sram[220]->out sram[221]->out sram[222]->out sram[223]->out sram[224]->out sram[225]->out sram[226]->out sram[227]->out sram[228]->out sram[229]->out sram[230]->out sram[231]->out sram[232]->out sram[233]->out sram[234]->out sram[235]->out sram[236]->out sram[237]->out sram[238]->out sram[239]->out sram[240]->out sram[241]->out sram[242]->out sram[243]->out sram[244]->out sram[245]->out sram[246]->out sram[247]->out sram[248]->out sram[249]->out sram[250]->out sram[251]->out sram[252]->out sram[253]->out sram[254]->out sram[255]->out sram[256]->out sram[257]->out sram[258]->out gvdd_lut6[3] sgnd lut6
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[3]_mode[n1_lut6]_ble6[0]_mode[ble6]_ff[0] ff[0]->D[0] ff[0]->Q[0] svdd sgnd
Xdff[3] 
***** BEGIN Global ports of SPICE_MODEL(static_dff) *****
+  Set[0]  Reset[0]  clk[0] 
***** END Global ports of SPICE_MODEL(static_dff) *****
+ ff[0]->D[0] ff[0]->Q[0] gvdd_dff[3] sgnd static_dff
.nodeset V(ff[0]->Q[0]) 0
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[3]_mode[n1_lut6]_ble6[0]_mode[ble6] mode[ble6]->in[0] mode[ble6]->in[1] mode[ble6]->in[2] mode[ble6]->in[3] mode[ble6]->in[4] mode[ble6]->in[5] mode[ble6]->out[0] mode[ble6]->clk[0] svdd sgnd
Xlut6[0] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[3]_mode[n1_lut6]_ble6[0]_mode[ble6]_lut6[0]
Xff[0] ff[0]->D[0] ff[0]->Q[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[3]_mode[n1_lut6]_ble6[0]_mode[ble6]_ff[0]
Xmux_1level_tapbuf_size2[3] ff[0]->Q[0] lut6[0]->out[0] mode[ble6]->out[0] sram[259]->outb sram[259]->out gvdd_local_interc sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[3], level=1, select_path_id=0. *****
*****1*****
Xsram[259] sram->in sram[259]->out sram[259]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[259]->out) 0
.nodeset V(sram[259]->outb) vsp
Xdirect_interc[48] mode[ble6]->in[0] lut6[0]->in[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[49] mode[ble6]->in[1] lut6[0]->in[1] gvdd_local_interc sgnd direct_interc
Xdirect_interc[50] mode[ble6]->in[2] lut6[0]->in[2] gvdd_local_interc sgnd direct_interc
Xdirect_interc[51] mode[ble6]->in[3] lut6[0]->in[3] gvdd_local_interc sgnd direct_interc
Xdirect_interc[52] mode[ble6]->in[4] lut6[0]->in[4] gvdd_local_interc sgnd direct_interc
Xdirect_interc[53] mode[ble6]->in[5] lut6[0]->in[5] gvdd_local_interc sgnd direct_interc
Xdirect_interc[54] lut6[0]->out[0] ff[0]->D[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[55] mode[ble6]->clk[0] ff[0]->clk[0] gvdd_local_interc sgnd direct_interc
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[3]_mode[n1_lut6] mode[n1_lut6]->in[0] mode[n1_lut6]->in[1] mode[n1_lut6]->in[2] mode[n1_lut6]->in[3] mode[n1_lut6]->in[4] mode[n1_lut6]->in[5] mode[n1_lut6]->out[0] mode[n1_lut6]->clk[0] svdd sgnd
Xble6[0] ble6[0]->in[0] ble6[0]->in[1] ble6[0]->in[2] ble6[0]->in[3] ble6[0]->in[4] ble6[0]->in[5] ble6[0]->out[0] ble6[0]->clk[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[3]_mode[n1_lut6]_ble6[0]_mode[ble6]
Xdirect_interc[56] ble6[0]->out[0] mode[n1_lut6]->out[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[57] mode[n1_lut6]->in[0] ble6[0]->in[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[58] mode[n1_lut6]->in[1] ble6[0]->in[1] gvdd_local_interc sgnd direct_interc
Xdirect_interc[59] mode[n1_lut6]->in[2] ble6[0]->in[2] gvdd_local_interc sgnd direct_interc
Xdirect_interc[60] mode[n1_lut6]->in[3] ble6[0]->in[3] gvdd_local_interc sgnd direct_interc
Xdirect_interc[61] mode[n1_lut6]->in[4] ble6[0]->in[4] gvdd_local_interc sgnd direct_interc
Xdirect_interc[62] mode[n1_lut6]->in[5] ble6[0]->in[5] gvdd_local_interc sgnd direct_interc
Xdirect_interc[63] mode[n1_lut6]->clk[0] ble6[0]->clk[0] gvdd_local_interc sgnd direct_interc
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[4]_mode[n1_lut6]_ble6[0]_mode[ble6]_lut6[0] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] svdd sgnd
***** Truth Table for LUT[4], size=6. *****
***** SRAM bits for LUT[4], size=6, num_sram=64. *****
*****0000000000000000000000000000000000000000000000000000000000000000*****
Xsram[260] sram->in sram[260]->out sram[260]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[260]->out) 0
.nodeset V(sram[260]->outb) vsp
Xsram[261] sram->in sram[261]->out sram[261]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[261]->out) 0
.nodeset V(sram[261]->outb) vsp
Xsram[262] sram->in sram[262]->out sram[262]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[262]->out) 0
.nodeset V(sram[262]->outb) vsp
Xsram[263] sram->in sram[263]->out sram[263]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[263]->out) 0
.nodeset V(sram[263]->outb) vsp
Xsram[264] sram->in sram[264]->out sram[264]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[264]->out) 0
.nodeset V(sram[264]->outb) vsp
Xsram[265] sram->in sram[265]->out sram[265]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[265]->out) 0
.nodeset V(sram[265]->outb) vsp
Xsram[266] sram->in sram[266]->out sram[266]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[266]->out) 0
.nodeset V(sram[266]->outb) vsp
Xsram[267] sram->in sram[267]->out sram[267]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[267]->out) 0
.nodeset V(sram[267]->outb) vsp
Xsram[268] sram->in sram[268]->out sram[268]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[268]->out) 0
.nodeset V(sram[268]->outb) vsp
Xsram[269] sram->in sram[269]->out sram[269]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[269]->out) 0
.nodeset V(sram[269]->outb) vsp
Xsram[270] sram->in sram[270]->out sram[270]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[270]->out) 0
.nodeset V(sram[270]->outb) vsp
Xsram[271] sram->in sram[271]->out sram[271]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[271]->out) 0
.nodeset V(sram[271]->outb) vsp
Xsram[272] sram->in sram[272]->out sram[272]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[272]->out) 0
.nodeset V(sram[272]->outb) vsp
Xsram[273] sram->in sram[273]->out sram[273]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[273]->out) 0
.nodeset V(sram[273]->outb) vsp
Xsram[274] sram->in sram[274]->out sram[274]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[274]->out) 0
.nodeset V(sram[274]->outb) vsp
Xsram[275] sram->in sram[275]->out sram[275]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[275]->out) 0
.nodeset V(sram[275]->outb) vsp
Xsram[276] sram->in sram[276]->out sram[276]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[276]->out) 0
.nodeset V(sram[276]->outb) vsp
Xsram[277] sram->in sram[277]->out sram[277]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[277]->out) 0
.nodeset V(sram[277]->outb) vsp
Xsram[278] sram->in sram[278]->out sram[278]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[278]->out) 0
.nodeset V(sram[278]->outb) vsp
Xsram[279] sram->in sram[279]->out sram[279]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[279]->out) 0
.nodeset V(sram[279]->outb) vsp
Xsram[280] sram->in sram[280]->out sram[280]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[280]->out) 0
.nodeset V(sram[280]->outb) vsp
Xsram[281] sram->in sram[281]->out sram[281]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[281]->out) 0
.nodeset V(sram[281]->outb) vsp
Xsram[282] sram->in sram[282]->out sram[282]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[282]->out) 0
.nodeset V(sram[282]->outb) vsp
Xsram[283] sram->in sram[283]->out sram[283]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[283]->out) 0
.nodeset V(sram[283]->outb) vsp
Xsram[284] sram->in sram[284]->out sram[284]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[284]->out) 0
.nodeset V(sram[284]->outb) vsp
Xsram[285] sram->in sram[285]->out sram[285]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[285]->out) 0
.nodeset V(sram[285]->outb) vsp
Xsram[286] sram->in sram[286]->out sram[286]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[286]->out) 0
.nodeset V(sram[286]->outb) vsp
Xsram[287] sram->in sram[287]->out sram[287]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[287]->out) 0
.nodeset V(sram[287]->outb) vsp
Xsram[288] sram->in sram[288]->out sram[288]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[288]->out) 0
.nodeset V(sram[288]->outb) vsp
Xsram[289] sram->in sram[289]->out sram[289]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[289]->out) 0
.nodeset V(sram[289]->outb) vsp
Xsram[290] sram->in sram[290]->out sram[290]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[290]->out) 0
.nodeset V(sram[290]->outb) vsp
Xsram[291] sram->in sram[291]->out sram[291]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[291]->out) 0
.nodeset V(sram[291]->outb) vsp
Xsram[292] sram->in sram[292]->out sram[292]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[292]->out) 0
.nodeset V(sram[292]->outb) vsp
Xsram[293] sram->in sram[293]->out sram[293]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[293]->out) 0
.nodeset V(sram[293]->outb) vsp
Xsram[294] sram->in sram[294]->out sram[294]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[294]->out) 0
.nodeset V(sram[294]->outb) vsp
Xsram[295] sram->in sram[295]->out sram[295]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[295]->out) 0
.nodeset V(sram[295]->outb) vsp
Xsram[296] sram->in sram[296]->out sram[296]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[296]->out) 0
.nodeset V(sram[296]->outb) vsp
Xsram[297] sram->in sram[297]->out sram[297]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[297]->out) 0
.nodeset V(sram[297]->outb) vsp
Xsram[298] sram->in sram[298]->out sram[298]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[298]->out) 0
.nodeset V(sram[298]->outb) vsp
Xsram[299] sram->in sram[299]->out sram[299]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[299]->out) 0
.nodeset V(sram[299]->outb) vsp
Xsram[300] sram->in sram[300]->out sram[300]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[300]->out) 0
.nodeset V(sram[300]->outb) vsp
Xsram[301] sram->in sram[301]->out sram[301]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[301]->out) 0
.nodeset V(sram[301]->outb) vsp
Xsram[302] sram->in sram[302]->out sram[302]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[302]->out) 0
.nodeset V(sram[302]->outb) vsp
Xsram[303] sram->in sram[303]->out sram[303]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[303]->out) 0
.nodeset V(sram[303]->outb) vsp
Xsram[304] sram->in sram[304]->out sram[304]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[304]->out) 0
.nodeset V(sram[304]->outb) vsp
Xsram[305] sram->in sram[305]->out sram[305]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[305]->out) 0
.nodeset V(sram[305]->outb) vsp
Xsram[306] sram->in sram[306]->out sram[306]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[306]->out) 0
.nodeset V(sram[306]->outb) vsp
Xsram[307] sram->in sram[307]->out sram[307]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[307]->out) 0
.nodeset V(sram[307]->outb) vsp
Xsram[308] sram->in sram[308]->out sram[308]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[308]->out) 0
.nodeset V(sram[308]->outb) vsp
Xsram[309] sram->in sram[309]->out sram[309]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[309]->out) 0
.nodeset V(sram[309]->outb) vsp
Xsram[310] sram->in sram[310]->out sram[310]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[310]->out) 0
.nodeset V(sram[310]->outb) vsp
Xsram[311] sram->in sram[311]->out sram[311]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[311]->out) 0
.nodeset V(sram[311]->outb) vsp
Xsram[312] sram->in sram[312]->out sram[312]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[312]->out) 0
.nodeset V(sram[312]->outb) vsp
Xsram[313] sram->in sram[313]->out sram[313]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[313]->out) 0
.nodeset V(sram[313]->outb) vsp
Xsram[314] sram->in sram[314]->out sram[314]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[314]->out) 0
.nodeset V(sram[314]->outb) vsp
Xsram[315] sram->in sram[315]->out sram[315]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[315]->out) 0
.nodeset V(sram[315]->outb) vsp
Xsram[316] sram->in sram[316]->out sram[316]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[316]->out) 0
.nodeset V(sram[316]->outb) vsp
Xsram[317] sram->in sram[317]->out sram[317]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[317]->out) 0
.nodeset V(sram[317]->outb) vsp
Xsram[318] sram->in sram[318]->out sram[318]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[318]->out) 0
.nodeset V(sram[318]->outb) vsp
Xsram[319] sram->in sram[319]->out sram[319]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[319]->out) 0
.nodeset V(sram[319]->outb) vsp
Xsram[320] sram->in sram[320]->out sram[320]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[320]->out) 0
.nodeset V(sram[320]->outb) vsp
Xsram[321] sram->in sram[321]->out sram[321]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[321]->out) 0
.nodeset V(sram[321]->outb) vsp
Xsram[322] sram->in sram[322]->out sram[322]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[322]->out) 0
.nodeset V(sram[322]->outb) vsp
Xsram[323] sram->in sram[323]->out sram[323]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[323]->out) 0
.nodeset V(sram[323]->outb) vsp
Xlut6[4] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] sram[260]->out sram[261]->out sram[262]->out sram[263]->out sram[264]->out sram[265]->out sram[266]->out sram[267]->out sram[268]->out sram[269]->out sram[270]->out sram[271]->out sram[272]->out sram[273]->out sram[274]->out sram[275]->out sram[276]->out sram[277]->out sram[278]->out sram[279]->out sram[280]->out sram[281]->out sram[282]->out sram[283]->out sram[284]->out sram[285]->out sram[286]->out sram[287]->out sram[288]->out sram[289]->out sram[290]->out sram[291]->out sram[292]->out sram[293]->out sram[294]->out sram[295]->out sram[296]->out sram[297]->out sram[298]->out sram[299]->out sram[300]->out sram[301]->out sram[302]->out sram[303]->out sram[304]->out sram[305]->out sram[306]->out sram[307]->out sram[308]->out sram[309]->out sram[310]->out sram[311]->out sram[312]->out sram[313]->out sram[314]->out sram[315]->out sram[316]->out sram[317]->out sram[318]->out sram[319]->out sram[320]->out sram[321]->out sram[322]->out sram[323]->out gvdd_lut6[4] sgnd lut6
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[4]_mode[n1_lut6]_ble6[0]_mode[ble6]_ff[0] ff[0]->D[0] ff[0]->Q[0] svdd sgnd
Xdff[4] 
***** BEGIN Global ports of SPICE_MODEL(static_dff) *****
+  Set[0]  Reset[0]  clk[0] 
***** END Global ports of SPICE_MODEL(static_dff) *****
+ ff[0]->D[0] ff[0]->Q[0] gvdd_dff[4] sgnd static_dff
.nodeset V(ff[0]->Q[0]) 0
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[4]_mode[n1_lut6]_ble6[0]_mode[ble6] mode[ble6]->in[0] mode[ble6]->in[1] mode[ble6]->in[2] mode[ble6]->in[3] mode[ble6]->in[4] mode[ble6]->in[5] mode[ble6]->out[0] mode[ble6]->clk[0] svdd sgnd
Xlut6[0] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[4]_mode[n1_lut6]_ble6[0]_mode[ble6]_lut6[0]
Xff[0] ff[0]->D[0] ff[0]->Q[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[4]_mode[n1_lut6]_ble6[0]_mode[ble6]_ff[0]
Xmux_1level_tapbuf_size2[4] ff[0]->Q[0] lut6[0]->out[0] mode[ble6]->out[0] sram[324]->outb sram[324]->out gvdd_local_interc sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[4], level=1, select_path_id=0. *****
*****1*****
Xsram[324] sram->in sram[324]->out sram[324]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[324]->out) 0
.nodeset V(sram[324]->outb) vsp
Xdirect_interc[64] mode[ble6]->in[0] lut6[0]->in[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[65] mode[ble6]->in[1] lut6[0]->in[1] gvdd_local_interc sgnd direct_interc
Xdirect_interc[66] mode[ble6]->in[2] lut6[0]->in[2] gvdd_local_interc sgnd direct_interc
Xdirect_interc[67] mode[ble6]->in[3] lut6[0]->in[3] gvdd_local_interc sgnd direct_interc
Xdirect_interc[68] mode[ble6]->in[4] lut6[0]->in[4] gvdd_local_interc sgnd direct_interc
Xdirect_interc[69] mode[ble6]->in[5] lut6[0]->in[5] gvdd_local_interc sgnd direct_interc
Xdirect_interc[70] lut6[0]->out[0] ff[0]->D[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[71] mode[ble6]->clk[0] ff[0]->clk[0] gvdd_local_interc sgnd direct_interc
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[4]_mode[n1_lut6] mode[n1_lut6]->in[0] mode[n1_lut6]->in[1] mode[n1_lut6]->in[2] mode[n1_lut6]->in[3] mode[n1_lut6]->in[4] mode[n1_lut6]->in[5] mode[n1_lut6]->out[0] mode[n1_lut6]->clk[0] svdd sgnd
Xble6[0] ble6[0]->in[0] ble6[0]->in[1] ble6[0]->in[2] ble6[0]->in[3] ble6[0]->in[4] ble6[0]->in[5] ble6[0]->out[0] ble6[0]->clk[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[4]_mode[n1_lut6]_ble6[0]_mode[ble6]
Xdirect_interc[72] ble6[0]->out[0] mode[n1_lut6]->out[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[73] mode[n1_lut6]->in[0] ble6[0]->in[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[74] mode[n1_lut6]->in[1] ble6[0]->in[1] gvdd_local_interc sgnd direct_interc
Xdirect_interc[75] mode[n1_lut6]->in[2] ble6[0]->in[2] gvdd_local_interc sgnd direct_interc
Xdirect_interc[76] mode[n1_lut6]->in[3] ble6[0]->in[3] gvdd_local_interc sgnd direct_interc
Xdirect_interc[77] mode[n1_lut6]->in[4] ble6[0]->in[4] gvdd_local_interc sgnd direct_interc
Xdirect_interc[78] mode[n1_lut6]->in[5] ble6[0]->in[5] gvdd_local_interc sgnd direct_interc
Xdirect_interc[79] mode[n1_lut6]->clk[0] ble6[0]->clk[0] gvdd_local_interc sgnd direct_interc
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[5]_mode[n1_lut6]_ble6[0]_mode[ble6]_lut6[0] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] svdd sgnd
***** Truth Table for LUT[5], size=6. *****
***** SRAM bits for LUT[5], size=6, num_sram=64. *****
*****0000000000000000000000000000000000000000000000000000000000000000*****
Xsram[325] sram->in sram[325]->out sram[325]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[325]->out) 0
.nodeset V(sram[325]->outb) vsp
Xsram[326] sram->in sram[326]->out sram[326]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[326]->out) 0
.nodeset V(sram[326]->outb) vsp
Xsram[327] sram->in sram[327]->out sram[327]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[327]->out) 0
.nodeset V(sram[327]->outb) vsp
Xsram[328] sram->in sram[328]->out sram[328]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[328]->out) 0
.nodeset V(sram[328]->outb) vsp
Xsram[329] sram->in sram[329]->out sram[329]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[329]->out) 0
.nodeset V(sram[329]->outb) vsp
Xsram[330] sram->in sram[330]->out sram[330]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[330]->out) 0
.nodeset V(sram[330]->outb) vsp
Xsram[331] sram->in sram[331]->out sram[331]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[331]->out) 0
.nodeset V(sram[331]->outb) vsp
Xsram[332] sram->in sram[332]->out sram[332]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[332]->out) 0
.nodeset V(sram[332]->outb) vsp
Xsram[333] sram->in sram[333]->out sram[333]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[333]->out) 0
.nodeset V(sram[333]->outb) vsp
Xsram[334] sram->in sram[334]->out sram[334]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[334]->out) 0
.nodeset V(sram[334]->outb) vsp
Xsram[335] sram->in sram[335]->out sram[335]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[335]->out) 0
.nodeset V(sram[335]->outb) vsp
Xsram[336] sram->in sram[336]->out sram[336]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[336]->out) 0
.nodeset V(sram[336]->outb) vsp
Xsram[337] sram->in sram[337]->out sram[337]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[337]->out) 0
.nodeset V(sram[337]->outb) vsp
Xsram[338] sram->in sram[338]->out sram[338]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[338]->out) 0
.nodeset V(sram[338]->outb) vsp
Xsram[339] sram->in sram[339]->out sram[339]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[339]->out) 0
.nodeset V(sram[339]->outb) vsp
Xsram[340] sram->in sram[340]->out sram[340]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[340]->out) 0
.nodeset V(sram[340]->outb) vsp
Xsram[341] sram->in sram[341]->out sram[341]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[341]->out) 0
.nodeset V(sram[341]->outb) vsp
Xsram[342] sram->in sram[342]->out sram[342]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[342]->out) 0
.nodeset V(sram[342]->outb) vsp
Xsram[343] sram->in sram[343]->out sram[343]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[343]->out) 0
.nodeset V(sram[343]->outb) vsp
Xsram[344] sram->in sram[344]->out sram[344]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[344]->out) 0
.nodeset V(sram[344]->outb) vsp
Xsram[345] sram->in sram[345]->out sram[345]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[345]->out) 0
.nodeset V(sram[345]->outb) vsp
Xsram[346] sram->in sram[346]->out sram[346]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[346]->out) 0
.nodeset V(sram[346]->outb) vsp
Xsram[347] sram->in sram[347]->out sram[347]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[347]->out) 0
.nodeset V(sram[347]->outb) vsp
Xsram[348] sram->in sram[348]->out sram[348]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[348]->out) 0
.nodeset V(sram[348]->outb) vsp
Xsram[349] sram->in sram[349]->out sram[349]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[349]->out) 0
.nodeset V(sram[349]->outb) vsp
Xsram[350] sram->in sram[350]->out sram[350]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[350]->out) 0
.nodeset V(sram[350]->outb) vsp
Xsram[351] sram->in sram[351]->out sram[351]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[351]->out) 0
.nodeset V(sram[351]->outb) vsp
Xsram[352] sram->in sram[352]->out sram[352]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[352]->out) 0
.nodeset V(sram[352]->outb) vsp
Xsram[353] sram->in sram[353]->out sram[353]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[353]->out) 0
.nodeset V(sram[353]->outb) vsp
Xsram[354] sram->in sram[354]->out sram[354]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[354]->out) 0
.nodeset V(sram[354]->outb) vsp
Xsram[355] sram->in sram[355]->out sram[355]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[355]->out) 0
.nodeset V(sram[355]->outb) vsp
Xsram[356] sram->in sram[356]->out sram[356]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[356]->out) 0
.nodeset V(sram[356]->outb) vsp
Xsram[357] sram->in sram[357]->out sram[357]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[357]->out) 0
.nodeset V(sram[357]->outb) vsp
Xsram[358] sram->in sram[358]->out sram[358]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[358]->out) 0
.nodeset V(sram[358]->outb) vsp
Xsram[359] sram->in sram[359]->out sram[359]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[359]->out) 0
.nodeset V(sram[359]->outb) vsp
Xsram[360] sram->in sram[360]->out sram[360]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[360]->out) 0
.nodeset V(sram[360]->outb) vsp
Xsram[361] sram->in sram[361]->out sram[361]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[361]->out) 0
.nodeset V(sram[361]->outb) vsp
Xsram[362] sram->in sram[362]->out sram[362]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[362]->out) 0
.nodeset V(sram[362]->outb) vsp
Xsram[363] sram->in sram[363]->out sram[363]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[363]->out) 0
.nodeset V(sram[363]->outb) vsp
Xsram[364] sram->in sram[364]->out sram[364]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[364]->out) 0
.nodeset V(sram[364]->outb) vsp
Xsram[365] sram->in sram[365]->out sram[365]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[365]->out) 0
.nodeset V(sram[365]->outb) vsp
Xsram[366] sram->in sram[366]->out sram[366]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[366]->out) 0
.nodeset V(sram[366]->outb) vsp
Xsram[367] sram->in sram[367]->out sram[367]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[367]->out) 0
.nodeset V(sram[367]->outb) vsp
Xsram[368] sram->in sram[368]->out sram[368]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[368]->out) 0
.nodeset V(sram[368]->outb) vsp
Xsram[369] sram->in sram[369]->out sram[369]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[369]->out) 0
.nodeset V(sram[369]->outb) vsp
Xsram[370] sram->in sram[370]->out sram[370]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[370]->out) 0
.nodeset V(sram[370]->outb) vsp
Xsram[371] sram->in sram[371]->out sram[371]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[371]->out) 0
.nodeset V(sram[371]->outb) vsp
Xsram[372] sram->in sram[372]->out sram[372]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[372]->out) 0
.nodeset V(sram[372]->outb) vsp
Xsram[373] sram->in sram[373]->out sram[373]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[373]->out) 0
.nodeset V(sram[373]->outb) vsp
Xsram[374] sram->in sram[374]->out sram[374]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[374]->out) 0
.nodeset V(sram[374]->outb) vsp
Xsram[375] sram->in sram[375]->out sram[375]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[375]->out) 0
.nodeset V(sram[375]->outb) vsp
Xsram[376] sram->in sram[376]->out sram[376]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[376]->out) 0
.nodeset V(sram[376]->outb) vsp
Xsram[377] sram->in sram[377]->out sram[377]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[377]->out) 0
.nodeset V(sram[377]->outb) vsp
Xsram[378] sram->in sram[378]->out sram[378]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[378]->out) 0
.nodeset V(sram[378]->outb) vsp
Xsram[379] sram->in sram[379]->out sram[379]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[379]->out) 0
.nodeset V(sram[379]->outb) vsp
Xsram[380] sram->in sram[380]->out sram[380]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[380]->out) 0
.nodeset V(sram[380]->outb) vsp
Xsram[381] sram->in sram[381]->out sram[381]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[381]->out) 0
.nodeset V(sram[381]->outb) vsp
Xsram[382] sram->in sram[382]->out sram[382]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[382]->out) 0
.nodeset V(sram[382]->outb) vsp
Xsram[383] sram->in sram[383]->out sram[383]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[383]->out) 0
.nodeset V(sram[383]->outb) vsp
Xsram[384] sram->in sram[384]->out sram[384]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[384]->out) 0
.nodeset V(sram[384]->outb) vsp
Xsram[385] sram->in sram[385]->out sram[385]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[385]->out) 0
.nodeset V(sram[385]->outb) vsp
Xsram[386] sram->in sram[386]->out sram[386]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[386]->out) 0
.nodeset V(sram[386]->outb) vsp
Xsram[387] sram->in sram[387]->out sram[387]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[387]->out) 0
.nodeset V(sram[387]->outb) vsp
Xsram[388] sram->in sram[388]->out sram[388]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[388]->out) 0
.nodeset V(sram[388]->outb) vsp
Xlut6[5] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] sram[325]->out sram[326]->out sram[327]->out sram[328]->out sram[329]->out sram[330]->out sram[331]->out sram[332]->out sram[333]->out sram[334]->out sram[335]->out sram[336]->out sram[337]->out sram[338]->out sram[339]->out sram[340]->out sram[341]->out sram[342]->out sram[343]->out sram[344]->out sram[345]->out sram[346]->out sram[347]->out sram[348]->out sram[349]->out sram[350]->out sram[351]->out sram[352]->out sram[353]->out sram[354]->out sram[355]->out sram[356]->out sram[357]->out sram[358]->out sram[359]->out sram[360]->out sram[361]->out sram[362]->out sram[363]->out sram[364]->out sram[365]->out sram[366]->out sram[367]->out sram[368]->out sram[369]->out sram[370]->out sram[371]->out sram[372]->out sram[373]->out sram[374]->out sram[375]->out sram[376]->out sram[377]->out sram[378]->out sram[379]->out sram[380]->out sram[381]->out sram[382]->out sram[383]->out sram[384]->out sram[385]->out sram[386]->out sram[387]->out sram[388]->out gvdd_lut6[5] sgnd lut6
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[5]_mode[n1_lut6]_ble6[0]_mode[ble6]_ff[0] ff[0]->D[0] ff[0]->Q[0] svdd sgnd
Xdff[5] 
***** BEGIN Global ports of SPICE_MODEL(static_dff) *****
+  Set[0]  Reset[0]  clk[0] 
***** END Global ports of SPICE_MODEL(static_dff) *****
+ ff[0]->D[0] ff[0]->Q[0] gvdd_dff[5] sgnd static_dff
.nodeset V(ff[0]->Q[0]) 0
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[5]_mode[n1_lut6]_ble6[0]_mode[ble6] mode[ble6]->in[0] mode[ble6]->in[1] mode[ble6]->in[2] mode[ble6]->in[3] mode[ble6]->in[4] mode[ble6]->in[5] mode[ble6]->out[0] mode[ble6]->clk[0] svdd sgnd
Xlut6[0] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[5]_mode[n1_lut6]_ble6[0]_mode[ble6]_lut6[0]
Xff[0] ff[0]->D[0] ff[0]->Q[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[5]_mode[n1_lut6]_ble6[0]_mode[ble6]_ff[0]
Xmux_1level_tapbuf_size2[5] ff[0]->Q[0] lut6[0]->out[0] mode[ble6]->out[0] sram[389]->outb sram[389]->out gvdd_local_interc sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[5], level=1, select_path_id=0. *****
*****1*****
Xsram[389] sram->in sram[389]->out sram[389]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[389]->out) 0
.nodeset V(sram[389]->outb) vsp
Xdirect_interc[80] mode[ble6]->in[0] lut6[0]->in[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[81] mode[ble6]->in[1] lut6[0]->in[1] gvdd_local_interc sgnd direct_interc
Xdirect_interc[82] mode[ble6]->in[2] lut6[0]->in[2] gvdd_local_interc sgnd direct_interc
Xdirect_interc[83] mode[ble6]->in[3] lut6[0]->in[3] gvdd_local_interc sgnd direct_interc
Xdirect_interc[84] mode[ble6]->in[4] lut6[0]->in[4] gvdd_local_interc sgnd direct_interc
Xdirect_interc[85] mode[ble6]->in[5] lut6[0]->in[5] gvdd_local_interc sgnd direct_interc
Xdirect_interc[86] lut6[0]->out[0] ff[0]->D[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[87] mode[ble6]->clk[0] ff[0]->clk[0] gvdd_local_interc sgnd direct_interc
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[5]_mode[n1_lut6] mode[n1_lut6]->in[0] mode[n1_lut6]->in[1] mode[n1_lut6]->in[2] mode[n1_lut6]->in[3] mode[n1_lut6]->in[4] mode[n1_lut6]->in[5] mode[n1_lut6]->out[0] mode[n1_lut6]->clk[0] svdd sgnd
Xble6[0] ble6[0]->in[0] ble6[0]->in[1] ble6[0]->in[2] ble6[0]->in[3] ble6[0]->in[4] ble6[0]->in[5] ble6[0]->out[0] ble6[0]->clk[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[5]_mode[n1_lut6]_ble6[0]_mode[ble6]
Xdirect_interc[88] ble6[0]->out[0] mode[n1_lut6]->out[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[89] mode[n1_lut6]->in[0] ble6[0]->in[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[90] mode[n1_lut6]->in[1] ble6[0]->in[1] gvdd_local_interc sgnd direct_interc
Xdirect_interc[91] mode[n1_lut6]->in[2] ble6[0]->in[2] gvdd_local_interc sgnd direct_interc
Xdirect_interc[92] mode[n1_lut6]->in[3] ble6[0]->in[3] gvdd_local_interc sgnd direct_interc
Xdirect_interc[93] mode[n1_lut6]->in[4] ble6[0]->in[4] gvdd_local_interc sgnd direct_interc
Xdirect_interc[94] mode[n1_lut6]->in[5] ble6[0]->in[5] gvdd_local_interc sgnd direct_interc
Xdirect_interc[95] mode[n1_lut6]->clk[0] ble6[0]->clk[0] gvdd_local_interc sgnd direct_interc
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[6]_mode[n1_lut6]_ble6[0]_mode[ble6]_lut6[0] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] svdd sgnd
***** Truth Table for LUT[6], size=6. *****
***** SRAM bits for LUT[6], size=6, num_sram=64. *****
*****0000000000000000000000000000000000000000000000000000000000000000*****
Xsram[390] sram->in sram[390]->out sram[390]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[390]->out) 0
.nodeset V(sram[390]->outb) vsp
Xsram[391] sram->in sram[391]->out sram[391]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[391]->out) 0
.nodeset V(sram[391]->outb) vsp
Xsram[392] sram->in sram[392]->out sram[392]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[392]->out) 0
.nodeset V(sram[392]->outb) vsp
Xsram[393] sram->in sram[393]->out sram[393]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[393]->out) 0
.nodeset V(sram[393]->outb) vsp
Xsram[394] sram->in sram[394]->out sram[394]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[394]->out) 0
.nodeset V(sram[394]->outb) vsp
Xsram[395] sram->in sram[395]->out sram[395]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[395]->out) 0
.nodeset V(sram[395]->outb) vsp
Xsram[396] sram->in sram[396]->out sram[396]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[396]->out) 0
.nodeset V(sram[396]->outb) vsp
Xsram[397] sram->in sram[397]->out sram[397]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[397]->out) 0
.nodeset V(sram[397]->outb) vsp
Xsram[398] sram->in sram[398]->out sram[398]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[398]->out) 0
.nodeset V(sram[398]->outb) vsp
Xsram[399] sram->in sram[399]->out sram[399]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[399]->out) 0
.nodeset V(sram[399]->outb) vsp
Xsram[400] sram->in sram[400]->out sram[400]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[400]->out) 0
.nodeset V(sram[400]->outb) vsp
Xsram[401] sram->in sram[401]->out sram[401]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[401]->out) 0
.nodeset V(sram[401]->outb) vsp
Xsram[402] sram->in sram[402]->out sram[402]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[402]->out) 0
.nodeset V(sram[402]->outb) vsp
Xsram[403] sram->in sram[403]->out sram[403]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[403]->out) 0
.nodeset V(sram[403]->outb) vsp
Xsram[404] sram->in sram[404]->out sram[404]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[404]->out) 0
.nodeset V(sram[404]->outb) vsp
Xsram[405] sram->in sram[405]->out sram[405]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[405]->out) 0
.nodeset V(sram[405]->outb) vsp
Xsram[406] sram->in sram[406]->out sram[406]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[406]->out) 0
.nodeset V(sram[406]->outb) vsp
Xsram[407] sram->in sram[407]->out sram[407]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[407]->out) 0
.nodeset V(sram[407]->outb) vsp
Xsram[408] sram->in sram[408]->out sram[408]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[408]->out) 0
.nodeset V(sram[408]->outb) vsp
Xsram[409] sram->in sram[409]->out sram[409]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[409]->out) 0
.nodeset V(sram[409]->outb) vsp
Xsram[410] sram->in sram[410]->out sram[410]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[410]->out) 0
.nodeset V(sram[410]->outb) vsp
Xsram[411] sram->in sram[411]->out sram[411]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[411]->out) 0
.nodeset V(sram[411]->outb) vsp
Xsram[412] sram->in sram[412]->out sram[412]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[412]->out) 0
.nodeset V(sram[412]->outb) vsp
Xsram[413] sram->in sram[413]->out sram[413]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[413]->out) 0
.nodeset V(sram[413]->outb) vsp
Xsram[414] sram->in sram[414]->out sram[414]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[414]->out) 0
.nodeset V(sram[414]->outb) vsp
Xsram[415] sram->in sram[415]->out sram[415]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[415]->out) 0
.nodeset V(sram[415]->outb) vsp
Xsram[416] sram->in sram[416]->out sram[416]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[416]->out) 0
.nodeset V(sram[416]->outb) vsp
Xsram[417] sram->in sram[417]->out sram[417]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[417]->out) 0
.nodeset V(sram[417]->outb) vsp
Xsram[418] sram->in sram[418]->out sram[418]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[418]->out) 0
.nodeset V(sram[418]->outb) vsp
Xsram[419] sram->in sram[419]->out sram[419]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[419]->out) 0
.nodeset V(sram[419]->outb) vsp
Xsram[420] sram->in sram[420]->out sram[420]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[420]->out) 0
.nodeset V(sram[420]->outb) vsp
Xsram[421] sram->in sram[421]->out sram[421]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[421]->out) 0
.nodeset V(sram[421]->outb) vsp
Xsram[422] sram->in sram[422]->out sram[422]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[422]->out) 0
.nodeset V(sram[422]->outb) vsp
Xsram[423] sram->in sram[423]->out sram[423]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[423]->out) 0
.nodeset V(sram[423]->outb) vsp
Xsram[424] sram->in sram[424]->out sram[424]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[424]->out) 0
.nodeset V(sram[424]->outb) vsp
Xsram[425] sram->in sram[425]->out sram[425]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[425]->out) 0
.nodeset V(sram[425]->outb) vsp
Xsram[426] sram->in sram[426]->out sram[426]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[426]->out) 0
.nodeset V(sram[426]->outb) vsp
Xsram[427] sram->in sram[427]->out sram[427]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[427]->out) 0
.nodeset V(sram[427]->outb) vsp
Xsram[428] sram->in sram[428]->out sram[428]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[428]->out) 0
.nodeset V(sram[428]->outb) vsp
Xsram[429] sram->in sram[429]->out sram[429]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[429]->out) 0
.nodeset V(sram[429]->outb) vsp
Xsram[430] sram->in sram[430]->out sram[430]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[430]->out) 0
.nodeset V(sram[430]->outb) vsp
Xsram[431] sram->in sram[431]->out sram[431]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[431]->out) 0
.nodeset V(sram[431]->outb) vsp
Xsram[432] sram->in sram[432]->out sram[432]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[432]->out) 0
.nodeset V(sram[432]->outb) vsp
Xsram[433] sram->in sram[433]->out sram[433]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[433]->out) 0
.nodeset V(sram[433]->outb) vsp
Xsram[434] sram->in sram[434]->out sram[434]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[434]->out) 0
.nodeset V(sram[434]->outb) vsp
Xsram[435] sram->in sram[435]->out sram[435]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[435]->out) 0
.nodeset V(sram[435]->outb) vsp
Xsram[436] sram->in sram[436]->out sram[436]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[436]->out) 0
.nodeset V(sram[436]->outb) vsp
Xsram[437] sram->in sram[437]->out sram[437]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[437]->out) 0
.nodeset V(sram[437]->outb) vsp
Xsram[438] sram->in sram[438]->out sram[438]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[438]->out) 0
.nodeset V(sram[438]->outb) vsp
Xsram[439] sram->in sram[439]->out sram[439]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[439]->out) 0
.nodeset V(sram[439]->outb) vsp
Xsram[440] sram->in sram[440]->out sram[440]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[440]->out) 0
.nodeset V(sram[440]->outb) vsp
Xsram[441] sram->in sram[441]->out sram[441]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[441]->out) 0
.nodeset V(sram[441]->outb) vsp
Xsram[442] sram->in sram[442]->out sram[442]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[442]->out) 0
.nodeset V(sram[442]->outb) vsp
Xsram[443] sram->in sram[443]->out sram[443]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[443]->out) 0
.nodeset V(sram[443]->outb) vsp
Xsram[444] sram->in sram[444]->out sram[444]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[444]->out) 0
.nodeset V(sram[444]->outb) vsp
Xsram[445] sram->in sram[445]->out sram[445]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[445]->out) 0
.nodeset V(sram[445]->outb) vsp
Xsram[446] sram->in sram[446]->out sram[446]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[446]->out) 0
.nodeset V(sram[446]->outb) vsp
Xsram[447] sram->in sram[447]->out sram[447]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[447]->out) 0
.nodeset V(sram[447]->outb) vsp
Xsram[448] sram->in sram[448]->out sram[448]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[448]->out) 0
.nodeset V(sram[448]->outb) vsp
Xsram[449] sram->in sram[449]->out sram[449]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[449]->out) 0
.nodeset V(sram[449]->outb) vsp
Xsram[450] sram->in sram[450]->out sram[450]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[450]->out) 0
.nodeset V(sram[450]->outb) vsp
Xsram[451] sram->in sram[451]->out sram[451]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[451]->out) 0
.nodeset V(sram[451]->outb) vsp
Xsram[452] sram->in sram[452]->out sram[452]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[452]->out) 0
.nodeset V(sram[452]->outb) vsp
Xsram[453] sram->in sram[453]->out sram[453]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[453]->out) 0
.nodeset V(sram[453]->outb) vsp
Xlut6[6] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] sram[390]->out sram[391]->out sram[392]->out sram[393]->out sram[394]->out sram[395]->out sram[396]->out sram[397]->out sram[398]->out sram[399]->out sram[400]->out sram[401]->out sram[402]->out sram[403]->out sram[404]->out sram[405]->out sram[406]->out sram[407]->out sram[408]->out sram[409]->out sram[410]->out sram[411]->out sram[412]->out sram[413]->out sram[414]->out sram[415]->out sram[416]->out sram[417]->out sram[418]->out sram[419]->out sram[420]->out sram[421]->out sram[422]->out sram[423]->out sram[424]->out sram[425]->out sram[426]->out sram[427]->out sram[428]->out sram[429]->out sram[430]->out sram[431]->out sram[432]->out sram[433]->out sram[434]->out sram[435]->out sram[436]->out sram[437]->out sram[438]->out sram[439]->out sram[440]->out sram[441]->out sram[442]->out sram[443]->out sram[444]->out sram[445]->out sram[446]->out sram[447]->out sram[448]->out sram[449]->out sram[450]->out sram[451]->out sram[452]->out sram[453]->out gvdd_lut6[6] sgnd lut6
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[6]_mode[n1_lut6]_ble6[0]_mode[ble6]_ff[0] ff[0]->D[0] ff[0]->Q[0] svdd sgnd
Xdff[6] 
***** BEGIN Global ports of SPICE_MODEL(static_dff) *****
+  Set[0]  Reset[0]  clk[0] 
***** END Global ports of SPICE_MODEL(static_dff) *****
+ ff[0]->D[0] ff[0]->Q[0] gvdd_dff[6] sgnd static_dff
.nodeset V(ff[0]->Q[0]) 0
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[6]_mode[n1_lut6]_ble6[0]_mode[ble6] mode[ble6]->in[0] mode[ble6]->in[1] mode[ble6]->in[2] mode[ble6]->in[3] mode[ble6]->in[4] mode[ble6]->in[5] mode[ble6]->out[0] mode[ble6]->clk[0] svdd sgnd
Xlut6[0] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[6]_mode[n1_lut6]_ble6[0]_mode[ble6]_lut6[0]
Xff[0] ff[0]->D[0] ff[0]->Q[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[6]_mode[n1_lut6]_ble6[0]_mode[ble6]_ff[0]
Xmux_1level_tapbuf_size2[6] ff[0]->Q[0] lut6[0]->out[0] mode[ble6]->out[0] sram[454]->outb sram[454]->out gvdd_local_interc sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[6], level=1, select_path_id=0. *****
*****1*****
Xsram[454] sram->in sram[454]->out sram[454]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[454]->out) 0
.nodeset V(sram[454]->outb) vsp
Xdirect_interc[96] mode[ble6]->in[0] lut6[0]->in[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[97] mode[ble6]->in[1] lut6[0]->in[1] gvdd_local_interc sgnd direct_interc
Xdirect_interc[98] mode[ble6]->in[2] lut6[0]->in[2] gvdd_local_interc sgnd direct_interc
Xdirect_interc[99] mode[ble6]->in[3] lut6[0]->in[3] gvdd_local_interc sgnd direct_interc
Xdirect_interc[100] mode[ble6]->in[4] lut6[0]->in[4] gvdd_local_interc sgnd direct_interc
Xdirect_interc[101] mode[ble6]->in[5] lut6[0]->in[5] gvdd_local_interc sgnd direct_interc
Xdirect_interc[102] lut6[0]->out[0] ff[0]->D[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[103] mode[ble6]->clk[0] ff[0]->clk[0] gvdd_local_interc sgnd direct_interc
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[6]_mode[n1_lut6] mode[n1_lut6]->in[0] mode[n1_lut6]->in[1] mode[n1_lut6]->in[2] mode[n1_lut6]->in[3] mode[n1_lut6]->in[4] mode[n1_lut6]->in[5] mode[n1_lut6]->out[0] mode[n1_lut6]->clk[0] svdd sgnd
Xble6[0] ble6[0]->in[0] ble6[0]->in[1] ble6[0]->in[2] ble6[0]->in[3] ble6[0]->in[4] ble6[0]->in[5] ble6[0]->out[0] ble6[0]->clk[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[6]_mode[n1_lut6]_ble6[0]_mode[ble6]
Xdirect_interc[104] ble6[0]->out[0] mode[n1_lut6]->out[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[105] mode[n1_lut6]->in[0] ble6[0]->in[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[106] mode[n1_lut6]->in[1] ble6[0]->in[1] gvdd_local_interc sgnd direct_interc
Xdirect_interc[107] mode[n1_lut6]->in[2] ble6[0]->in[2] gvdd_local_interc sgnd direct_interc
Xdirect_interc[108] mode[n1_lut6]->in[3] ble6[0]->in[3] gvdd_local_interc sgnd direct_interc
Xdirect_interc[109] mode[n1_lut6]->in[4] ble6[0]->in[4] gvdd_local_interc sgnd direct_interc
Xdirect_interc[110] mode[n1_lut6]->in[5] ble6[0]->in[5] gvdd_local_interc sgnd direct_interc
Xdirect_interc[111] mode[n1_lut6]->clk[0] ble6[0]->clk[0] gvdd_local_interc sgnd direct_interc
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[7]_mode[n1_lut6]_ble6[0]_mode[ble6]_lut6[0] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] svdd sgnd
***** Truth Table for LUT[7], size=6. *****
***** SRAM bits for LUT[7], size=6, num_sram=64. *****
*****0000000000000000000000000000000000000000000000000000000000000000*****
Xsram[455] sram->in sram[455]->out sram[455]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[455]->out) 0
.nodeset V(sram[455]->outb) vsp
Xsram[456] sram->in sram[456]->out sram[456]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[456]->out) 0
.nodeset V(sram[456]->outb) vsp
Xsram[457] sram->in sram[457]->out sram[457]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[457]->out) 0
.nodeset V(sram[457]->outb) vsp
Xsram[458] sram->in sram[458]->out sram[458]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[458]->out) 0
.nodeset V(sram[458]->outb) vsp
Xsram[459] sram->in sram[459]->out sram[459]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[459]->out) 0
.nodeset V(sram[459]->outb) vsp
Xsram[460] sram->in sram[460]->out sram[460]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[460]->out) 0
.nodeset V(sram[460]->outb) vsp
Xsram[461] sram->in sram[461]->out sram[461]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[461]->out) 0
.nodeset V(sram[461]->outb) vsp
Xsram[462] sram->in sram[462]->out sram[462]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[462]->out) 0
.nodeset V(sram[462]->outb) vsp
Xsram[463] sram->in sram[463]->out sram[463]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[463]->out) 0
.nodeset V(sram[463]->outb) vsp
Xsram[464] sram->in sram[464]->out sram[464]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[464]->out) 0
.nodeset V(sram[464]->outb) vsp
Xsram[465] sram->in sram[465]->out sram[465]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[465]->out) 0
.nodeset V(sram[465]->outb) vsp
Xsram[466] sram->in sram[466]->out sram[466]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[466]->out) 0
.nodeset V(sram[466]->outb) vsp
Xsram[467] sram->in sram[467]->out sram[467]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[467]->out) 0
.nodeset V(sram[467]->outb) vsp
Xsram[468] sram->in sram[468]->out sram[468]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[468]->out) 0
.nodeset V(sram[468]->outb) vsp
Xsram[469] sram->in sram[469]->out sram[469]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[469]->out) 0
.nodeset V(sram[469]->outb) vsp
Xsram[470] sram->in sram[470]->out sram[470]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[470]->out) 0
.nodeset V(sram[470]->outb) vsp
Xsram[471] sram->in sram[471]->out sram[471]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[471]->out) 0
.nodeset V(sram[471]->outb) vsp
Xsram[472] sram->in sram[472]->out sram[472]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[472]->out) 0
.nodeset V(sram[472]->outb) vsp
Xsram[473] sram->in sram[473]->out sram[473]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[473]->out) 0
.nodeset V(sram[473]->outb) vsp
Xsram[474] sram->in sram[474]->out sram[474]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[474]->out) 0
.nodeset V(sram[474]->outb) vsp
Xsram[475] sram->in sram[475]->out sram[475]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[475]->out) 0
.nodeset V(sram[475]->outb) vsp
Xsram[476] sram->in sram[476]->out sram[476]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[476]->out) 0
.nodeset V(sram[476]->outb) vsp
Xsram[477] sram->in sram[477]->out sram[477]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[477]->out) 0
.nodeset V(sram[477]->outb) vsp
Xsram[478] sram->in sram[478]->out sram[478]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[478]->out) 0
.nodeset V(sram[478]->outb) vsp
Xsram[479] sram->in sram[479]->out sram[479]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[479]->out) 0
.nodeset V(sram[479]->outb) vsp
Xsram[480] sram->in sram[480]->out sram[480]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[480]->out) 0
.nodeset V(sram[480]->outb) vsp
Xsram[481] sram->in sram[481]->out sram[481]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[481]->out) 0
.nodeset V(sram[481]->outb) vsp
Xsram[482] sram->in sram[482]->out sram[482]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[482]->out) 0
.nodeset V(sram[482]->outb) vsp
Xsram[483] sram->in sram[483]->out sram[483]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[483]->out) 0
.nodeset V(sram[483]->outb) vsp
Xsram[484] sram->in sram[484]->out sram[484]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[484]->out) 0
.nodeset V(sram[484]->outb) vsp
Xsram[485] sram->in sram[485]->out sram[485]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[485]->out) 0
.nodeset V(sram[485]->outb) vsp
Xsram[486] sram->in sram[486]->out sram[486]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[486]->out) 0
.nodeset V(sram[486]->outb) vsp
Xsram[487] sram->in sram[487]->out sram[487]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[487]->out) 0
.nodeset V(sram[487]->outb) vsp
Xsram[488] sram->in sram[488]->out sram[488]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[488]->out) 0
.nodeset V(sram[488]->outb) vsp
Xsram[489] sram->in sram[489]->out sram[489]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[489]->out) 0
.nodeset V(sram[489]->outb) vsp
Xsram[490] sram->in sram[490]->out sram[490]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[490]->out) 0
.nodeset V(sram[490]->outb) vsp
Xsram[491] sram->in sram[491]->out sram[491]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[491]->out) 0
.nodeset V(sram[491]->outb) vsp
Xsram[492] sram->in sram[492]->out sram[492]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[492]->out) 0
.nodeset V(sram[492]->outb) vsp
Xsram[493] sram->in sram[493]->out sram[493]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[493]->out) 0
.nodeset V(sram[493]->outb) vsp
Xsram[494] sram->in sram[494]->out sram[494]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[494]->out) 0
.nodeset V(sram[494]->outb) vsp
Xsram[495] sram->in sram[495]->out sram[495]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[495]->out) 0
.nodeset V(sram[495]->outb) vsp
Xsram[496] sram->in sram[496]->out sram[496]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[496]->out) 0
.nodeset V(sram[496]->outb) vsp
Xsram[497] sram->in sram[497]->out sram[497]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[497]->out) 0
.nodeset V(sram[497]->outb) vsp
Xsram[498] sram->in sram[498]->out sram[498]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[498]->out) 0
.nodeset V(sram[498]->outb) vsp
Xsram[499] sram->in sram[499]->out sram[499]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[499]->out) 0
.nodeset V(sram[499]->outb) vsp
Xsram[500] sram->in sram[500]->out sram[500]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[500]->out) 0
.nodeset V(sram[500]->outb) vsp
Xsram[501] sram->in sram[501]->out sram[501]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[501]->out) 0
.nodeset V(sram[501]->outb) vsp
Xsram[502] sram->in sram[502]->out sram[502]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[502]->out) 0
.nodeset V(sram[502]->outb) vsp
Xsram[503] sram->in sram[503]->out sram[503]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[503]->out) 0
.nodeset V(sram[503]->outb) vsp
Xsram[504] sram->in sram[504]->out sram[504]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[504]->out) 0
.nodeset V(sram[504]->outb) vsp
Xsram[505] sram->in sram[505]->out sram[505]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[505]->out) 0
.nodeset V(sram[505]->outb) vsp
Xsram[506] sram->in sram[506]->out sram[506]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[506]->out) 0
.nodeset V(sram[506]->outb) vsp
Xsram[507] sram->in sram[507]->out sram[507]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[507]->out) 0
.nodeset V(sram[507]->outb) vsp
Xsram[508] sram->in sram[508]->out sram[508]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[508]->out) 0
.nodeset V(sram[508]->outb) vsp
Xsram[509] sram->in sram[509]->out sram[509]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[509]->out) 0
.nodeset V(sram[509]->outb) vsp
Xsram[510] sram->in sram[510]->out sram[510]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[510]->out) 0
.nodeset V(sram[510]->outb) vsp
Xsram[511] sram->in sram[511]->out sram[511]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[511]->out) 0
.nodeset V(sram[511]->outb) vsp
Xsram[512] sram->in sram[512]->out sram[512]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[512]->out) 0
.nodeset V(sram[512]->outb) vsp
Xsram[513] sram->in sram[513]->out sram[513]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[513]->out) 0
.nodeset V(sram[513]->outb) vsp
Xsram[514] sram->in sram[514]->out sram[514]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[514]->out) 0
.nodeset V(sram[514]->outb) vsp
Xsram[515] sram->in sram[515]->out sram[515]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[515]->out) 0
.nodeset V(sram[515]->outb) vsp
Xsram[516] sram->in sram[516]->out sram[516]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[516]->out) 0
.nodeset V(sram[516]->outb) vsp
Xsram[517] sram->in sram[517]->out sram[517]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[517]->out) 0
.nodeset V(sram[517]->outb) vsp
Xsram[518] sram->in sram[518]->out sram[518]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[518]->out) 0
.nodeset V(sram[518]->outb) vsp
Xlut6[7] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] sram[455]->out sram[456]->out sram[457]->out sram[458]->out sram[459]->out sram[460]->out sram[461]->out sram[462]->out sram[463]->out sram[464]->out sram[465]->out sram[466]->out sram[467]->out sram[468]->out sram[469]->out sram[470]->out sram[471]->out sram[472]->out sram[473]->out sram[474]->out sram[475]->out sram[476]->out sram[477]->out sram[478]->out sram[479]->out sram[480]->out sram[481]->out sram[482]->out sram[483]->out sram[484]->out sram[485]->out sram[486]->out sram[487]->out sram[488]->out sram[489]->out sram[490]->out sram[491]->out sram[492]->out sram[493]->out sram[494]->out sram[495]->out sram[496]->out sram[497]->out sram[498]->out sram[499]->out sram[500]->out sram[501]->out sram[502]->out sram[503]->out sram[504]->out sram[505]->out sram[506]->out sram[507]->out sram[508]->out sram[509]->out sram[510]->out sram[511]->out sram[512]->out sram[513]->out sram[514]->out sram[515]->out sram[516]->out sram[517]->out sram[518]->out gvdd_lut6[7] sgnd lut6
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[7]_mode[n1_lut6]_ble6[0]_mode[ble6]_ff[0] ff[0]->D[0] ff[0]->Q[0] svdd sgnd
Xdff[7] 
***** BEGIN Global ports of SPICE_MODEL(static_dff) *****
+  Set[0]  Reset[0]  clk[0] 
***** END Global ports of SPICE_MODEL(static_dff) *****
+ ff[0]->D[0] ff[0]->Q[0] gvdd_dff[7] sgnd static_dff
.nodeset V(ff[0]->Q[0]) 0
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[7]_mode[n1_lut6]_ble6[0]_mode[ble6] mode[ble6]->in[0] mode[ble6]->in[1] mode[ble6]->in[2] mode[ble6]->in[3] mode[ble6]->in[4] mode[ble6]->in[5] mode[ble6]->out[0] mode[ble6]->clk[0] svdd sgnd
Xlut6[0] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[7]_mode[n1_lut6]_ble6[0]_mode[ble6]_lut6[0]
Xff[0] ff[0]->D[0] ff[0]->Q[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[7]_mode[n1_lut6]_ble6[0]_mode[ble6]_ff[0]
Xmux_1level_tapbuf_size2[7] ff[0]->Q[0] lut6[0]->out[0] mode[ble6]->out[0] sram[519]->outb sram[519]->out gvdd_local_interc sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[7], level=1, select_path_id=0. *****
*****1*****
Xsram[519] sram->in sram[519]->out sram[519]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[519]->out) 0
.nodeset V(sram[519]->outb) vsp
Xdirect_interc[112] mode[ble6]->in[0] lut6[0]->in[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[113] mode[ble6]->in[1] lut6[0]->in[1] gvdd_local_interc sgnd direct_interc
Xdirect_interc[114] mode[ble6]->in[2] lut6[0]->in[2] gvdd_local_interc sgnd direct_interc
Xdirect_interc[115] mode[ble6]->in[3] lut6[0]->in[3] gvdd_local_interc sgnd direct_interc
Xdirect_interc[116] mode[ble6]->in[4] lut6[0]->in[4] gvdd_local_interc sgnd direct_interc
Xdirect_interc[117] mode[ble6]->in[5] lut6[0]->in[5] gvdd_local_interc sgnd direct_interc
Xdirect_interc[118] lut6[0]->out[0] ff[0]->D[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[119] mode[ble6]->clk[0] ff[0]->clk[0] gvdd_local_interc sgnd direct_interc
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[7]_mode[n1_lut6] mode[n1_lut6]->in[0] mode[n1_lut6]->in[1] mode[n1_lut6]->in[2] mode[n1_lut6]->in[3] mode[n1_lut6]->in[4] mode[n1_lut6]->in[5] mode[n1_lut6]->out[0] mode[n1_lut6]->clk[0] svdd sgnd
Xble6[0] ble6[0]->in[0] ble6[0]->in[1] ble6[0]->in[2] ble6[0]->in[3] ble6[0]->in[4] ble6[0]->in[5] ble6[0]->out[0] ble6[0]->clk[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[7]_mode[n1_lut6]_ble6[0]_mode[ble6]
Xdirect_interc[120] ble6[0]->out[0] mode[n1_lut6]->out[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[121] mode[n1_lut6]->in[0] ble6[0]->in[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[122] mode[n1_lut6]->in[1] ble6[0]->in[1] gvdd_local_interc sgnd direct_interc
Xdirect_interc[123] mode[n1_lut6]->in[2] ble6[0]->in[2] gvdd_local_interc sgnd direct_interc
Xdirect_interc[124] mode[n1_lut6]->in[3] ble6[0]->in[3] gvdd_local_interc sgnd direct_interc
Xdirect_interc[125] mode[n1_lut6]->in[4] ble6[0]->in[4] gvdd_local_interc sgnd direct_interc
Xdirect_interc[126] mode[n1_lut6]->in[5] ble6[0]->in[5] gvdd_local_interc sgnd direct_interc
Xdirect_interc[127] mode[n1_lut6]->clk[0] ble6[0]->clk[0] gvdd_local_interc sgnd direct_interc
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[8]_mode[n1_lut6]_ble6[0]_mode[ble6]_lut6[0] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] svdd sgnd
***** Truth Table for LUT[8], size=6. *****
***** SRAM bits for LUT[8], size=6, num_sram=64. *****
*****0000000000000000000000000000000000000000000000000000000000000000*****
Xsram[520] sram->in sram[520]->out sram[520]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[520]->out) 0
.nodeset V(sram[520]->outb) vsp
Xsram[521] sram->in sram[521]->out sram[521]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[521]->out) 0
.nodeset V(sram[521]->outb) vsp
Xsram[522] sram->in sram[522]->out sram[522]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[522]->out) 0
.nodeset V(sram[522]->outb) vsp
Xsram[523] sram->in sram[523]->out sram[523]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[523]->out) 0
.nodeset V(sram[523]->outb) vsp
Xsram[524] sram->in sram[524]->out sram[524]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[524]->out) 0
.nodeset V(sram[524]->outb) vsp
Xsram[525] sram->in sram[525]->out sram[525]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[525]->out) 0
.nodeset V(sram[525]->outb) vsp
Xsram[526] sram->in sram[526]->out sram[526]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[526]->out) 0
.nodeset V(sram[526]->outb) vsp
Xsram[527] sram->in sram[527]->out sram[527]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[527]->out) 0
.nodeset V(sram[527]->outb) vsp
Xsram[528] sram->in sram[528]->out sram[528]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[528]->out) 0
.nodeset V(sram[528]->outb) vsp
Xsram[529] sram->in sram[529]->out sram[529]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[529]->out) 0
.nodeset V(sram[529]->outb) vsp
Xsram[530] sram->in sram[530]->out sram[530]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[530]->out) 0
.nodeset V(sram[530]->outb) vsp
Xsram[531] sram->in sram[531]->out sram[531]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[531]->out) 0
.nodeset V(sram[531]->outb) vsp
Xsram[532] sram->in sram[532]->out sram[532]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[532]->out) 0
.nodeset V(sram[532]->outb) vsp
Xsram[533] sram->in sram[533]->out sram[533]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[533]->out) 0
.nodeset V(sram[533]->outb) vsp
Xsram[534] sram->in sram[534]->out sram[534]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[534]->out) 0
.nodeset V(sram[534]->outb) vsp
Xsram[535] sram->in sram[535]->out sram[535]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[535]->out) 0
.nodeset V(sram[535]->outb) vsp
Xsram[536] sram->in sram[536]->out sram[536]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[536]->out) 0
.nodeset V(sram[536]->outb) vsp
Xsram[537] sram->in sram[537]->out sram[537]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[537]->out) 0
.nodeset V(sram[537]->outb) vsp
Xsram[538] sram->in sram[538]->out sram[538]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[538]->out) 0
.nodeset V(sram[538]->outb) vsp
Xsram[539] sram->in sram[539]->out sram[539]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[539]->out) 0
.nodeset V(sram[539]->outb) vsp
Xsram[540] sram->in sram[540]->out sram[540]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[540]->out) 0
.nodeset V(sram[540]->outb) vsp
Xsram[541] sram->in sram[541]->out sram[541]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[541]->out) 0
.nodeset V(sram[541]->outb) vsp
Xsram[542] sram->in sram[542]->out sram[542]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[542]->out) 0
.nodeset V(sram[542]->outb) vsp
Xsram[543] sram->in sram[543]->out sram[543]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[543]->out) 0
.nodeset V(sram[543]->outb) vsp
Xsram[544] sram->in sram[544]->out sram[544]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[544]->out) 0
.nodeset V(sram[544]->outb) vsp
Xsram[545] sram->in sram[545]->out sram[545]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[545]->out) 0
.nodeset V(sram[545]->outb) vsp
Xsram[546] sram->in sram[546]->out sram[546]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[546]->out) 0
.nodeset V(sram[546]->outb) vsp
Xsram[547] sram->in sram[547]->out sram[547]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[547]->out) 0
.nodeset V(sram[547]->outb) vsp
Xsram[548] sram->in sram[548]->out sram[548]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[548]->out) 0
.nodeset V(sram[548]->outb) vsp
Xsram[549] sram->in sram[549]->out sram[549]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[549]->out) 0
.nodeset V(sram[549]->outb) vsp
Xsram[550] sram->in sram[550]->out sram[550]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[550]->out) 0
.nodeset V(sram[550]->outb) vsp
Xsram[551] sram->in sram[551]->out sram[551]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[551]->out) 0
.nodeset V(sram[551]->outb) vsp
Xsram[552] sram->in sram[552]->out sram[552]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[552]->out) 0
.nodeset V(sram[552]->outb) vsp
Xsram[553] sram->in sram[553]->out sram[553]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[553]->out) 0
.nodeset V(sram[553]->outb) vsp
Xsram[554] sram->in sram[554]->out sram[554]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[554]->out) 0
.nodeset V(sram[554]->outb) vsp
Xsram[555] sram->in sram[555]->out sram[555]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[555]->out) 0
.nodeset V(sram[555]->outb) vsp
Xsram[556] sram->in sram[556]->out sram[556]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[556]->out) 0
.nodeset V(sram[556]->outb) vsp
Xsram[557] sram->in sram[557]->out sram[557]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[557]->out) 0
.nodeset V(sram[557]->outb) vsp
Xsram[558] sram->in sram[558]->out sram[558]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[558]->out) 0
.nodeset V(sram[558]->outb) vsp
Xsram[559] sram->in sram[559]->out sram[559]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[559]->out) 0
.nodeset V(sram[559]->outb) vsp
Xsram[560] sram->in sram[560]->out sram[560]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[560]->out) 0
.nodeset V(sram[560]->outb) vsp
Xsram[561] sram->in sram[561]->out sram[561]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[561]->out) 0
.nodeset V(sram[561]->outb) vsp
Xsram[562] sram->in sram[562]->out sram[562]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[562]->out) 0
.nodeset V(sram[562]->outb) vsp
Xsram[563] sram->in sram[563]->out sram[563]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[563]->out) 0
.nodeset V(sram[563]->outb) vsp
Xsram[564] sram->in sram[564]->out sram[564]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[564]->out) 0
.nodeset V(sram[564]->outb) vsp
Xsram[565] sram->in sram[565]->out sram[565]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[565]->out) 0
.nodeset V(sram[565]->outb) vsp
Xsram[566] sram->in sram[566]->out sram[566]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[566]->out) 0
.nodeset V(sram[566]->outb) vsp
Xsram[567] sram->in sram[567]->out sram[567]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[567]->out) 0
.nodeset V(sram[567]->outb) vsp
Xsram[568] sram->in sram[568]->out sram[568]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[568]->out) 0
.nodeset V(sram[568]->outb) vsp
Xsram[569] sram->in sram[569]->out sram[569]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[569]->out) 0
.nodeset V(sram[569]->outb) vsp
Xsram[570] sram->in sram[570]->out sram[570]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[570]->out) 0
.nodeset V(sram[570]->outb) vsp
Xsram[571] sram->in sram[571]->out sram[571]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[571]->out) 0
.nodeset V(sram[571]->outb) vsp
Xsram[572] sram->in sram[572]->out sram[572]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[572]->out) 0
.nodeset V(sram[572]->outb) vsp
Xsram[573] sram->in sram[573]->out sram[573]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[573]->out) 0
.nodeset V(sram[573]->outb) vsp
Xsram[574] sram->in sram[574]->out sram[574]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[574]->out) 0
.nodeset V(sram[574]->outb) vsp
Xsram[575] sram->in sram[575]->out sram[575]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[575]->out) 0
.nodeset V(sram[575]->outb) vsp
Xsram[576] sram->in sram[576]->out sram[576]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[576]->out) 0
.nodeset V(sram[576]->outb) vsp
Xsram[577] sram->in sram[577]->out sram[577]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[577]->out) 0
.nodeset V(sram[577]->outb) vsp
Xsram[578] sram->in sram[578]->out sram[578]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[578]->out) 0
.nodeset V(sram[578]->outb) vsp
Xsram[579] sram->in sram[579]->out sram[579]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[579]->out) 0
.nodeset V(sram[579]->outb) vsp
Xsram[580] sram->in sram[580]->out sram[580]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[580]->out) 0
.nodeset V(sram[580]->outb) vsp
Xsram[581] sram->in sram[581]->out sram[581]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[581]->out) 0
.nodeset V(sram[581]->outb) vsp
Xsram[582] sram->in sram[582]->out sram[582]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[582]->out) 0
.nodeset V(sram[582]->outb) vsp
Xsram[583] sram->in sram[583]->out sram[583]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[583]->out) 0
.nodeset V(sram[583]->outb) vsp
Xlut6[8] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] sram[520]->out sram[521]->out sram[522]->out sram[523]->out sram[524]->out sram[525]->out sram[526]->out sram[527]->out sram[528]->out sram[529]->out sram[530]->out sram[531]->out sram[532]->out sram[533]->out sram[534]->out sram[535]->out sram[536]->out sram[537]->out sram[538]->out sram[539]->out sram[540]->out sram[541]->out sram[542]->out sram[543]->out sram[544]->out sram[545]->out sram[546]->out sram[547]->out sram[548]->out sram[549]->out sram[550]->out sram[551]->out sram[552]->out sram[553]->out sram[554]->out sram[555]->out sram[556]->out sram[557]->out sram[558]->out sram[559]->out sram[560]->out sram[561]->out sram[562]->out sram[563]->out sram[564]->out sram[565]->out sram[566]->out sram[567]->out sram[568]->out sram[569]->out sram[570]->out sram[571]->out sram[572]->out sram[573]->out sram[574]->out sram[575]->out sram[576]->out sram[577]->out sram[578]->out sram[579]->out sram[580]->out sram[581]->out sram[582]->out sram[583]->out gvdd_lut6[8] sgnd lut6
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[8]_mode[n1_lut6]_ble6[0]_mode[ble6]_ff[0] ff[0]->D[0] ff[0]->Q[0] svdd sgnd
Xdff[8] 
***** BEGIN Global ports of SPICE_MODEL(static_dff) *****
+  Set[0]  Reset[0]  clk[0] 
***** END Global ports of SPICE_MODEL(static_dff) *****
+ ff[0]->D[0] ff[0]->Q[0] gvdd_dff[8] sgnd static_dff
.nodeset V(ff[0]->Q[0]) 0
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[8]_mode[n1_lut6]_ble6[0]_mode[ble6] mode[ble6]->in[0] mode[ble6]->in[1] mode[ble6]->in[2] mode[ble6]->in[3] mode[ble6]->in[4] mode[ble6]->in[5] mode[ble6]->out[0] mode[ble6]->clk[0] svdd sgnd
Xlut6[0] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[8]_mode[n1_lut6]_ble6[0]_mode[ble6]_lut6[0]
Xff[0] ff[0]->D[0] ff[0]->Q[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[8]_mode[n1_lut6]_ble6[0]_mode[ble6]_ff[0]
Xmux_1level_tapbuf_size2[8] ff[0]->Q[0] lut6[0]->out[0] mode[ble6]->out[0] sram[584]->outb sram[584]->out gvdd_local_interc sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[8], level=1, select_path_id=0. *****
*****1*****
Xsram[584] sram->in sram[584]->out sram[584]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[584]->out) 0
.nodeset V(sram[584]->outb) vsp
Xdirect_interc[128] mode[ble6]->in[0] lut6[0]->in[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[129] mode[ble6]->in[1] lut6[0]->in[1] gvdd_local_interc sgnd direct_interc
Xdirect_interc[130] mode[ble6]->in[2] lut6[0]->in[2] gvdd_local_interc sgnd direct_interc
Xdirect_interc[131] mode[ble6]->in[3] lut6[0]->in[3] gvdd_local_interc sgnd direct_interc
Xdirect_interc[132] mode[ble6]->in[4] lut6[0]->in[4] gvdd_local_interc sgnd direct_interc
Xdirect_interc[133] mode[ble6]->in[5] lut6[0]->in[5] gvdd_local_interc sgnd direct_interc
Xdirect_interc[134] lut6[0]->out[0] ff[0]->D[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[135] mode[ble6]->clk[0] ff[0]->clk[0] gvdd_local_interc sgnd direct_interc
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[8]_mode[n1_lut6] mode[n1_lut6]->in[0] mode[n1_lut6]->in[1] mode[n1_lut6]->in[2] mode[n1_lut6]->in[3] mode[n1_lut6]->in[4] mode[n1_lut6]->in[5] mode[n1_lut6]->out[0] mode[n1_lut6]->clk[0] svdd sgnd
Xble6[0] ble6[0]->in[0] ble6[0]->in[1] ble6[0]->in[2] ble6[0]->in[3] ble6[0]->in[4] ble6[0]->in[5] ble6[0]->out[0] ble6[0]->clk[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[8]_mode[n1_lut6]_ble6[0]_mode[ble6]
Xdirect_interc[136] ble6[0]->out[0] mode[n1_lut6]->out[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[137] mode[n1_lut6]->in[0] ble6[0]->in[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[138] mode[n1_lut6]->in[1] ble6[0]->in[1] gvdd_local_interc sgnd direct_interc
Xdirect_interc[139] mode[n1_lut6]->in[2] ble6[0]->in[2] gvdd_local_interc sgnd direct_interc
Xdirect_interc[140] mode[n1_lut6]->in[3] ble6[0]->in[3] gvdd_local_interc sgnd direct_interc
Xdirect_interc[141] mode[n1_lut6]->in[4] ble6[0]->in[4] gvdd_local_interc sgnd direct_interc
Xdirect_interc[142] mode[n1_lut6]->in[5] ble6[0]->in[5] gvdd_local_interc sgnd direct_interc
Xdirect_interc[143] mode[n1_lut6]->clk[0] ble6[0]->clk[0] gvdd_local_interc sgnd direct_interc
.eom
***** Logical block mapped to this LUT: n7 *****
.subckt grid[1][1]_clb[0]_mode[clb]_fle[9]_mode[n1_lut6]_ble6[0]_mode[ble6]_lut6[0] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] svdd sgnd
***** Truth Table for LUT[9], size=6. *****
* 0----- 1 *
***** SRAM bits for LUT[9], size=6, num_sram=64. *****
*****0101010101010101010101010101010101010101010101010101010101010101*****
Xsram[585] sram->in sram[585]->out sram[585]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[585]->out) 0
.nodeset V(sram[585]->outb) vsp
Xsram[586] sram->in sram[586]->out sram[586]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[586]->out) 0
.nodeset V(sram[586]->outb) vsp
Xsram[587] sram->in sram[587]->out sram[587]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[587]->out) 0
.nodeset V(sram[587]->outb) vsp
Xsram[588] sram->in sram[588]->out sram[588]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[588]->out) 0
.nodeset V(sram[588]->outb) vsp
Xsram[589] sram->in sram[589]->out sram[589]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[589]->out) 0
.nodeset V(sram[589]->outb) vsp
Xsram[590] sram->in sram[590]->out sram[590]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[590]->out) 0
.nodeset V(sram[590]->outb) vsp
Xsram[591] sram->in sram[591]->out sram[591]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[591]->out) 0
.nodeset V(sram[591]->outb) vsp
Xsram[592] sram->in sram[592]->out sram[592]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[592]->out) 0
.nodeset V(sram[592]->outb) vsp
Xsram[593] sram->in sram[593]->out sram[593]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[593]->out) 0
.nodeset V(sram[593]->outb) vsp
Xsram[594] sram->in sram[594]->out sram[594]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[594]->out) 0
.nodeset V(sram[594]->outb) vsp
Xsram[595] sram->in sram[595]->out sram[595]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[595]->out) 0
.nodeset V(sram[595]->outb) vsp
Xsram[596] sram->in sram[596]->out sram[596]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[596]->out) 0
.nodeset V(sram[596]->outb) vsp
Xsram[597] sram->in sram[597]->out sram[597]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[597]->out) 0
.nodeset V(sram[597]->outb) vsp
Xsram[598] sram->in sram[598]->out sram[598]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[598]->out) 0
.nodeset V(sram[598]->outb) vsp
Xsram[599] sram->in sram[599]->out sram[599]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[599]->out) 0
.nodeset V(sram[599]->outb) vsp
Xsram[600] sram->in sram[600]->out sram[600]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[600]->out) 0
.nodeset V(sram[600]->outb) vsp
Xsram[601] sram->in sram[601]->out sram[601]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[601]->out) 0
.nodeset V(sram[601]->outb) vsp
Xsram[602] sram->in sram[602]->out sram[602]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[602]->out) 0
.nodeset V(sram[602]->outb) vsp
Xsram[603] sram->in sram[603]->out sram[603]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[603]->out) 0
.nodeset V(sram[603]->outb) vsp
Xsram[604] sram->in sram[604]->out sram[604]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[604]->out) 0
.nodeset V(sram[604]->outb) vsp
Xsram[605] sram->in sram[605]->out sram[605]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[605]->out) 0
.nodeset V(sram[605]->outb) vsp
Xsram[606] sram->in sram[606]->out sram[606]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[606]->out) 0
.nodeset V(sram[606]->outb) vsp
Xsram[607] sram->in sram[607]->out sram[607]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[607]->out) 0
.nodeset V(sram[607]->outb) vsp
Xsram[608] sram->in sram[608]->out sram[608]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[608]->out) 0
.nodeset V(sram[608]->outb) vsp
Xsram[609] sram->in sram[609]->out sram[609]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[609]->out) 0
.nodeset V(sram[609]->outb) vsp
Xsram[610] sram->in sram[610]->out sram[610]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[610]->out) 0
.nodeset V(sram[610]->outb) vsp
Xsram[611] sram->in sram[611]->out sram[611]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[611]->out) 0
.nodeset V(sram[611]->outb) vsp
Xsram[612] sram->in sram[612]->out sram[612]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[612]->out) 0
.nodeset V(sram[612]->outb) vsp
Xsram[613] sram->in sram[613]->out sram[613]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[613]->out) 0
.nodeset V(sram[613]->outb) vsp
Xsram[614] sram->in sram[614]->out sram[614]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[614]->out) 0
.nodeset V(sram[614]->outb) vsp
Xsram[615] sram->in sram[615]->out sram[615]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[615]->out) 0
.nodeset V(sram[615]->outb) vsp
Xsram[616] sram->in sram[616]->out sram[616]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[616]->out) 0
.nodeset V(sram[616]->outb) vsp
Xsram[617] sram->in sram[617]->out sram[617]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[617]->out) 0
.nodeset V(sram[617]->outb) vsp
Xsram[618] sram->in sram[618]->out sram[618]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[618]->out) 0
.nodeset V(sram[618]->outb) vsp
Xsram[619] sram->in sram[619]->out sram[619]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[619]->out) 0
.nodeset V(sram[619]->outb) vsp
Xsram[620] sram->in sram[620]->out sram[620]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[620]->out) 0
.nodeset V(sram[620]->outb) vsp
Xsram[621] sram->in sram[621]->out sram[621]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[621]->out) 0
.nodeset V(sram[621]->outb) vsp
Xsram[622] sram->in sram[622]->out sram[622]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[622]->out) 0
.nodeset V(sram[622]->outb) vsp
Xsram[623] sram->in sram[623]->out sram[623]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[623]->out) 0
.nodeset V(sram[623]->outb) vsp
Xsram[624] sram->in sram[624]->out sram[624]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[624]->out) 0
.nodeset V(sram[624]->outb) vsp
Xsram[625] sram->in sram[625]->out sram[625]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[625]->out) 0
.nodeset V(sram[625]->outb) vsp
Xsram[626] sram->in sram[626]->out sram[626]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[626]->out) 0
.nodeset V(sram[626]->outb) vsp
Xsram[627] sram->in sram[627]->out sram[627]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[627]->out) 0
.nodeset V(sram[627]->outb) vsp
Xsram[628] sram->in sram[628]->out sram[628]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[628]->out) 0
.nodeset V(sram[628]->outb) vsp
Xsram[629] sram->in sram[629]->out sram[629]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[629]->out) 0
.nodeset V(sram[629]->outb) vsp
Xsram[630] sram->in sram[630]->out sram[630]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[630]->out) 0
.nodeset V(sram[630]->outb) vsp
Xsram[631] sram->in sram[631]->out sram[631]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[631]->out) 0
.nodeset V(sram[631]->outb) vsp
Xsram[632] sram->in sram[632]->out sram[632]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[632]->out) 0
.nodeset V(sram[632]->outb) vsp
Xsram[633] sram->in sram[633]->out sram[633]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[633]->out) 0
.nodeset V(sram[633]->outb) vsp
Xsram[634] sram->in sram[634]->out sram[634]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[634]->out) 0
.nodeset V(sram[634]->outb) vsp
Xsram[635] sram->in sram[635]->out sram[635]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[635]->out) 0
.nodeset V(sram[635]->outb) vsp
Xsram[636] sram->in sram[636]->out sram[636]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[636]->out) 0
.nodeset V(sram[636]->outb) vsp
Xsram[637] sram->in sram[637]->out sram[637]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[637]->out) 0
.nodeset V(sram[637]->outb) vsp
Xsram[638] sram->in sram[638]->out sram[638]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[638]->out) 0
.nodeset V(sram[638]->outb) vsp
Xsram[639] sram->in sram[639]->out sram[639]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[639]->out) 0
.nodeset V(sram[639]->outb) vsp
Xsram[640] sram->in sram[640]->out sram[640]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[640]->out) 0
.nodeset V(sram[640]->outb) vsp
Xsram[641] sram->in sram[641]->out sram[641]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[641]->out) 0
.nodeset V(sram[641]->outb) vsp
Xsram[642] sram->in sram[642]->out sram[642]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[642]->out) 0
.nodeset V(sram[642]->outb) vsp
Xsram[643] sram->in sram[643]->out sram[643]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[643]->out) 0
.nodeset V(sram[643]->outb) vsp
Xsram[644] sram->in sram[644]->out sram[644]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[644]->out) 0
.nodeset V(sram[644]->outb) vsp
Xsram[645] sram->in sram[645]->out sram[645]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[645]->out) 0
.nodeset V(sram[645]->outb) vsp
Xsram[646] sram->in sram[646]->out sram[646]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[646]->out) 0
.nodeset V(sram[646]->outb) vsp
Xsram[647] sram->in sram[647]->out sram[647]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[647]->out) 0
.nodeset V(sram[647]->outb) vsp
Xsram[648] sram->in sram[648]->out sram[648]->outb gvdd_sram_luts sgnd  sram6T
.nodeset V(sram[648]->out) 0
.nodeset V(sram[648]->outb) vsp
Xlut6[9] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] sram[585]->out sram[586]->outb sram[587]->out sram[588]->outb sram[589]->out sram[590]->outb sram[591]->out sram[592]->outb sram[593]->out sram[594]->outb sram[595]->out sram[596]->outb sram[597]->out sram[598]->outb sram[599]->out sram[600]->outb sram[601]->out sram[602]->outb sram[603]->out sram[604]->outb sram[605]->out sram[606]->outb sram[607]->out sram[608]->outb sram[609]->out sram[610]->outb sram[611]->out sram[612]->outb sram[613]->out sram[614]->outb sram[615]->out sram[616]->outb sram[617]->out sram[618]->outb sram[619]->out sram[620]->outb sram[621]->out sram[622]->outb sram[623]->out sram[624]->outb sram[625]->out sram[626]->outb sram[627]->out sram[628]->outb sram[629]->out sram[630]->outb sram[631]->out sram[632]->outb sram[633]->out sram[634]->outb sram[635]->out sram[636]->outb sram[637]->out sram[638]->outb sram[639]->out sram[640]->outb sram[641]->out sram[642]->outb sram[643]->out sram[644]->outb sram[645]->out sram[646]->outb sram[647]->out sram[648]->outb gvdd_lut6[9] sgnd lut6
.eom
***** Logical block mapped to this FF: Q0 *****
.subckt grid[1][1]_clb[0]_mode[clb]_fle[9]_mode[n1_lut6]_ble6[0]_mode[ble6]_ff[0] ff[0]->D[0] ff[0]->Q[0] svdd sgnd
Xdff[9] 
***** BEGIN Global ports of SPICE_MODEL(static_dff) *****
+  Set[0]  Reset[0]  clk[0] 
***** END Global ports of SPICE_MODEL(static_dff) *****
+ ff[0]->D[0] ff[0]->Q[0] gvdd_dff[9] sgnd static_dff
.nodeset V(ff[0]->Q[0]) 0
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[9]_mode[n1_lut6]_ble6[0]_mode[ble6] mode[ble6]->in[0] mode[ble6]->in[1] mode[ble6]->in[2] mode[ble6]->in[3] mode[ble6]->in[4] mode[ble6]->in[5] mode[ble6]->out[0] mode[ble6]->clk[0] svdd sgnd
Xlut6[0] lut6[0]->in[0] lut6[0]->in[1] lut6[0]->in[2] lut6[0]->in[3] lut6[0]->in[4] lut6[0]->in[5] lut6[0]->out[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[9]_mode[n1_lut6]_ble6[0]_mode[ble6]_lut6[0]
Xff[0] ff[0]->D[0] ff[0]->Q[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[9]_mode[n1_lut6]_ble6[0]_mode[ble6]_ff[0]
Xmux_1level_tapbuf_size2[9] ff[0]->Q[0] lut6[0]->out[0] mode[ble6]->out[0] sram[649]->outb sram[649]->out gvdd_local_interc sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[9], level=1, select_path_id=0. *****
*****1*****
Xsram[649] sram->in sram[649]->out sram[649]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[649]->out) 0
.nodeset V(sram[649]->outb) vsp
Xdirect_interc[144] mode[ble6]->in[0] lut6[0]->in[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[145] mode[ble6]->in[1] lut6[0]->in[1] gvdd_local_interc sgnd direct_interc
Xdirect_interc[146] mode[ble6]->in[2] lut6[0]->in[2] gvdd_local_interc sgnd direct_interc
Xdirect_interc[147] mode[ble6]->in[3] lut6[0]->in[3] gvdd_local_interc sgnd direct_interc
Xdirect_interc[148] mode[ble6]->in[4] lut6[0]->in[4] gvdd_local_interc sgnd direct_interc
Xdirect_interc[149] mode[ble6]->in[5] lut6[0]->in[5] gvdd_local_interc sgnd direct_interc
Xdirect_interc[150] lut6[0]->out[0] ff[0]->D[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[151] mode[ble6]->clk[0] ff[0]->clk[0] gvdd_local_interc sgnd direct_interc
.eom
.subckt grid[1][1]_clb[0]_mode[clb]_fle[9]_mode[n1_lut6] mode[n1_lut6]->in[0] mode[n1_lut6]->in[1] mode[n1_lut6]->in[2] mode[n1_lut6]->in[3] mode[n1_lut6]->in[4] mode[n1_lut6]->in[5] mode[n1_lut6]->out[0] mode[n1_lut6]->clk[0] svdd sgnd
Xble6[0] ble6[0]->in[0] ble6[0]->in[1] ble6[0]->in[2] ble6[0]->in[3] ble6[0]->in[4] ble6[0]->in[5] ble6[0]->out[0] ble6[0]->clk[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[9]_mode[n1_lut6]_ble6[0]_mode[ble6]
Xdirect_interc[152] ble6[0]->out[0] mode[n1_lut6]->out[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[153] mode[n1_lut6]->in[0] ble6[0]->in[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[154] mode[n1_lut6]->in[1] ble6[0]->in[1] gvdd_local_interc sgnd direct_interc
Xdirect_interc[155] mode[n1_lut6]->in[2] ble6[0]->in[2] gvdd_local_interc sgnd direct_interc
Xdirect_interc[156] mode[n1_lut6]->in[3] ble6[0]->in[3] gvdd_local_interc sgnd direct_interc
Xdirect_interc[157] mode[n1_lut6]->in[4] ble6[0]->in[4] gvdd_local_interc sgnd direct_interc
Xdirect_interc[158] mode[n1_lut6]->in[5] ble6[0]->in[5] gvdd_local_interc sgnd direct_interc
Xdirect_interc[159] mode[n1_lut6]->clk[0] ble6[0]->clk[0] gvdd_local_interc sgnd direct_interc
.eom
.subckt grid[1][1]_clb[0]_mode[clb] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] mode[clb]->O[0] mode[clb]->O[1] mode[clb]->O[2] mode[clb]->O[3] mode[clb]->O[4] mode[clb]->O[5] mode[clb]->O[6] mode[clb]->O[7] mode[clb]->O[8] mode[clb]->O[9] mode[clb]->clk[0] svdd sgnd
Xfle[0] fle[0]->in[0] fle[0]->in[1] fle[0]->in[2] fle[0]->in[3] fle[0]->in[4] fle[0]->in[5] fle[0]->out[0] fle[0]->clk[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[0]_mode[n1_lut6]
Xfle[1] fle[1]->in[0] fle[1]->in[1] fle[1]->in[2] fle[1]->in[3] fle[1]->in[4] fle[1]->in[5] fle[1]->out[0] fle[1]->clk[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[1]_mode[n1_lut6]
Xfle[2] fle[2]->in[0] fle[2]->in[1] fle[2]->in[2] fle[2]->in[3] fle[2]->in[4] fle[2]->in[5] fle[2]->out[0] fle[2]->clk[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[2]_mode[n1_lut6]
Xfle[3] fle[3]->in[0] fle[3]->in[1] fle[3]->in[2] fle[3]->in[3] fle[3]->in[4] fle[3]->in[5] fle[3]->out[0] fle[3]->clk[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[3]_mode[n1_lut6]
Xfle[4] fle[4]->in[0] fle[4]->in[1] fle[4]->in[2] fle[4]->in[3] fle[4]->in[4] fle[4]->in[5] fle[4]->out[0] fle[4]->clk[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[4]_mode[n1_lut6]
Xfle[5] fle[5]->in[0] fle[5]->in[1] fle[5]->in[2] fle[5]->in[3] fle[5]->in[4] fle[5]->in[5] fle[5]->out[0] fle[5]->clk[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[5]_mode[n1_lut6]
Xfle[6] fle[6]->in[0] fle[6]->in[1] fle[6]->in[2] fle[6]->in[3] fle[6]->in[4] fle[6]->in[5] fle[6]->out[0] fle[6]->clk[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[6]_mode[n1_lut6]
Xfle[7] fle[7]->in[0] fle[7]->in[1] fle[7]->in[2] fle[7]->in[3] fle[7]->in[4] fle[7]->in[5] fle[7]->out[0] fle[7]->clk[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[7]_mode[n1_lut6]
Xfle[8] fle[8]->in[0] fle[8]->in[1] fle[8]->in[2] fle[8]->in[3] fle[8]->in[4] fle[8]->in[5] fle[8]->out[0] fle[8]->clk[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[8]_mode[n1_lut6]
Xfle[9] fle[9]->in[0] fle[9]->in[1] fle[9]->in[2] fle[9]->in[3] fle[9]->in[4] fle[9]->in[5] fle[9]->out[0] fle[9]->clk[0] svdd sgnd grid[1][1]_clb[0]_mode[clb]_fle[9]_mode[n1_lut6]
Xdirect_interc[160] fle[0]->out[0] mode[clb]->O[0] gvdd_local_interc sgnd direct_interc
Xdirect_interc[161] fle[1]->out[0] mode[clb]->O[1] gvdd_local_interc sgnd direct_interc
Xdirect_interc[162] fle[2]->out[0] mode[clb]->O[2] gvdd_local_interc sgnd direct_interc
Xdirect_interc[163] fle[3]->out[0] mode[clb]->O[3] gvdd_local_interc sgnd direct_interc
Xdirect_interc[164] fle[4]->out[0] mode[clb]->O[4] gvdd_local_interc sgnd direct_interc
Xdirect_interc[165] fle[5]->out[0] mode[clb]->O[5] gvdd_local_interc sgnd direct_interc
Xdirect_interc[166] fle[6]->out[0] mode[clb]->O[6] gvdd_local_interc sgnd direct_interc
Xdirect_interc[167] fle[7]->out[0] mode[clb]->O[7] gvdd_local_interc sgnd direct_interc
Xdirect_interc[168] fle[8]->out[0] mode[clb]->O[8] gvdd_local_interc sgnd direct_interc
Xdirect_interc[169] fle[9]->out[0] mode[clb]->O[9] gvdd_local_interc sgnd direct_interc
Xmux_2level_size50[0] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[0]->in[0] sram[650]->outb sram[650]->out sram[651]->out sram[651]->outb sram[652]->out sram[652]->outb sram[653]->out sram[653]->outb sram[654]->out sram[654]->outb sram[655]->out sram[655]->outb sram[656]->out sram[656]->outb sram[657]->out sram[657]->outb sram[658]->outb sram[658]->out sram[659]->out sram[659]->outb sram[660]->out sram[660]->outb sram[661]->out sram[661]->outb sram[662]->out sram[662]->outb sram[663]->out sram[663]->outb sram[664]->out sram[664]->outb sram[665]->out sram[665]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[0], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[650] sram->in sram[650]->out sram[650]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[650]->out) 0
.nodeset V(sram[650]->outb) vsp
Xsram[651] sram->in sram[651]->out sram[651]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[651]->out) 0
.nodeset V(sram[651]->outb) vsp
Xsram[652] sram->in sram[652]->out sram[652]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[652]->out) 0
.nodeset V(sram[652]->outb) vsp
Xsram[653] sram->in sram[653]->out sram[653]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[653]->out) 0
.nodeset V(sram[653]->outb) vsp
Xsram[654] sram->in sram[654]->out sram[654]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[654]->out) 0
.nodeset V(sram[654]->outb) vsp
Xsram[655] sram->in sram[655]->out sram[655]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[655]->out) 0
.nodeset V(sram[655]->outb) vsp
Xsram[656] sram->in sram[656]->out sram[656]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[656]->out) 0
.nodeset V(sram[656]->outb) vsp
Xsram[657] sram->in sram[657]->out sram[657]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[657]->out) 0
.nodeset V(sram[657]->outb) vsp
Xsram[658] sram->in sram[658]->out sram[658]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[658]->out) 0
.nodeset V(sram[658]->outb) vsp
Xsram[659] sram->in sram[659]->out sram[659]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[659]->out) 0
.nodeset V(sram[659]->outb) vsp
Xsram[660] sram->in sram[660]->out sram[660]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[660]->out) 0
.nodeset V(sram[660]->outb) vsp
Xsram[661] sram->in sram[661]->out sram[661]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[661]->out) 0
.nodeset V(sram[661]->outb) vsp
Xsram[662] sram->in sram[662]->out sram[662]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[662]->out) 0
.nodeset V(sram[662]->outb) vsp
Xsram[663] sram->in sram[663]->out sram[663]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[663]->out) 0
.nodeset V(sram[663]->outb) vsp
Xsram[664] sram->in sram[664]->out sram[664]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[664]->out) 0
.nodeset V(sram[664]->outb) vsp
Xsram[665] sram->in sram[665]->out sram[665]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[665]->out) 0
.nodeset V(sram[665]->outb) vsp
Xmux_2level_size50[1] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[0]->in[1] sram[666]->outb sram[666]->out sram[667]->out sram[667]->outb sram[668]->out sram[668]->outb sram[669]->out sram[669]->outb sram[670]->out sram[670]->outb sram[671]->out sram[671]->outb sram[672]->out sram[672]->outb sram[673]->out sram[673]->outb sram[674]->outb sram[674]->out sram[675]->out sram[675]->outb sram[676]->out sram[676]->outb sram[677]->out sram[677]->outb sram[678]->out sram[678]->outb sram[679]->out sram[679]->outb sram[680]->out sram[680]->outb sram[681]->out sram[681]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[1], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[666] sram->in sram[666]->out sram[666]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[666]->out) 0
.nodeset V(sram[666]->outb) vsp
Xsram[667] sram->in sram[667]->out sram[667]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[667]->out) 0
.nodeset V(sram[667]->outb) vsp
Xsram[668] sram->in sram[668]->out sram[668]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[668]->out) 0
.nodeset V(sram[668]->outb) vsp
Xsram[669] sram->in sram[669]->out sram[669]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[669]->out) 0
.nodeset V(sram[669]->outb) vsp
Xsram[670] sram->in sram[670]->out sram[670]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[670]->out) 0
.nodeset V(sram[670]->outb) vsp
Xsram[671] sram->in sram[671]->out sram[671]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[671]->out) 0
.nodeset V(sram[671]->outb) vsp
Xsram[672] sram->in sram[672]->out sram[672]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[672]->out) 0
.nodeset V(sram[672]->outb) vsp
Xsram[673] sram->in sram[673]->out sram[673]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[673]->out) 0
.nodeset V(sram[673]->outb) vsp
Xsram[674] sram->in sram[674]->out sram[674]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[674]->out) 0
.nodeset V(sram[674]->outb) vsp
Xsram[675] sram->in sram[675]->out sram[675]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[675]->out) 0
.nodeset V(sram[675]->outb) vsp
Xsram[676] sram->in sram[676]->out sram[676]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[676]->out) 0
.nodeset V(sram[676]->outb) vsp
Xsram[677] sram->in sram[677]->out sram[677]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[677]->out) 0
.nodeset V(sram[677]->outb) vsp
Xsram[678] sram->in sram[678]->out sram[678]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[678]->out) 0
.nodeset V(sram[678]->outb) vsp
Xsram[679] sram->in sram[679]->out sram[679]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[679]->out) 0
.nodeset V(sram[679]->outb) vsp
Xsram[680] sram->in sram[680]->out sram[680]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[680]->out) 0
.nodeset V(sram[680]->outb) vsp
Xsram[681] sram->in sram[681]->out sram[681]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[681]->out) 0
.nodeset V(sram[681]->outb) vsp
Xmux_2level_size50[2] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[0]->in[2] sram[682]->outb sram[682]->out sram[683]->out sram[683]->outb sram[684]->out sram[684]->outb sram[685]->out sram[685]->outb sram[686]->out sram[686]->outb sram[687]->out sram[687]->outb sram[688]->out sram[688]->outb sram[689]->out sram[689]->outb sram[690]->outb sram[690]->out sram[691]->out sram[691]->outb sram[692]->out sram[692]->outb sram[693]->out sram[693]->outb sram[694]->out sram[694]->outb sram[695]->out sram[695]->outb sram[696]->out sram[696]->outb sram[697]->out sram[697]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[2], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[682] sram->in sram[682]->out sram[682]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[682]->out) 0
.nodeset V(sram[682]->outb) vsp
Xsram[683] sram->in sram[683]->out sram[683]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[683]->out) 0
.nodeset V(sram[683]->outb) vsp
Xsram[684] sram->in sram[684]->out sram[684]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[684]->out) 0
.nodeset V(sram[684]->outb) vsp
Xsram[685] sram->in sram[685]->out sram[685]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[685]->out) 0
.nodeset V(sram[685]->outb) vsp
Xsram[686] sram->in sram[686]->out sram[686]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[686]->out) 0
.nodeset V(sram[686]->outb) vsp
Xsram[687] sram->in sram[687]->out sram[687]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[687]->out) 0
.nodeset V(sram[687]->outb) vsp
Xsram[688] sram->in sram[688]->out sram[688]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[688]->out) 0
.nodeset V(sram[688]->outb) vsp
Xsram[689] sram->in sram[689]->out sram[689]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[689]->out) 0
.nodeset V(sram[689]->outb) vsp
Xsram[690] sram->in sram[690]->out sram[690]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[690]->out) 0
.nodeset V(sram[690]->outb) vsp
Xsram[691] sram->in sram[691]->out sram[691]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[691]->out) 0
.nodeset V(sram[691]->outb) vsp
Xsram[692] sram->in sram[692]->out sram[692]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[692]->out) 0
.nodeset V(sram[692]->outb) vsp
Xsram[693] sram->in sram[693]->out sram[693]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[693]->out) 0
.nodeset V(sram[693]->outb) vsp
Xsram[694] sram->in sram[694]->out sram[694]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[694]->out) 0
.nodeset V(sram[694]->outb) vsp
Xsram[695] sram->in sram[695]->out sram[695]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[695]->out) 0
.nodeset V(sram[695]->outb) vsp
Xsram[696] sram->in sram[696]->out sram[696]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[696]->out) 0
.nodeset V(sram[696]->outb) vsp
Xsram[697] sram->in sram[697]->out sram[697]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[697]->out) 0
.nodeset V(sram[697]->outb) vsp
Xmux_2level_size50[3] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[0]->in[3] sram[698]->outb sram[698]->out sram[699]->out sram[699]->outb sram[700]->out sram[700]->outb sram[701]->out sram[701]->outb sram[702]->out sram[702]->outb sram[703]->out sram[703]->outb sram[704]->out sram[704]->outb sram[705]->out sram[705]->outb sram[706]->outb sram[706]->out sram[707]->out sram[707]->outb sram[708]->out sram[708]->outb sram[709]->out sram[709]->outb sram[710]->out sram[710]->outb sram[711]->out sram[711]->outb sram[712]->out sram[712]->outb sram[713]->out sram[713]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[3], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[698] sram->in sram[698]->out sram[698]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[698]->out) 0
.nodeset V(sram[698]->outb) vsp
Xsram[699] sram->in sram[699]->out sram[699]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[699]->out) 0
.nodeset V(sram[699]->outb) vsp
Xsram[700] sram->in sram[700]->out sram[700]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[700]->out) 0
.nodeset V(sram[700]->outb) vsp
Xsram[701] sram->in sram[701]->out sram[701]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[701]->out) 0
.nodeset V(sram[701]->outb) vsp
Xsram[702] sram->in sram[702]->out sram[702]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[702]->out) 0
.nodeset V(sram[702]->outb) vsp
Xsram[703] sram->in sram[703]->out sram[703]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[703]->out) 0
.nodeset V(sram[703]->outb) vsp
Xsram[704] sram->in sram[704]->out sram[704]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[704]->out) 0
.nodeset V(sram[704]->outb) vsp
Xsram[705] sram->in sram[705]->out sram[705]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[705]->out) 0
.nodeset V(sram[705]->outb) vsp
Xsram[706] sram->in sram[706]->out sram[706]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[706]->out) 0
.nodeset V(sram[706]->outb) vsp
Xsram[707] sram->in sram[707]->out sram[707]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[707]->out) 0
.nodeset V(sram[707]->outb) vsp
Xsram[708] sram->in sram[708]->out sram[708]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[708]->out) 0
.nodeset V(sram[708]->outb) vsp
Xsram[709] sram->in sram[709]->out sram[709]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[709]->out) 0
.nodeset V(sram[709]->outb) vsp
Xsram[710] sram->in sram[710]->out sram[710]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[710]->out) 0
.nodeset V(sram[710]->outb) vsp
Xsram[711] sram->in sram[711]->out sram[711]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[711]->out) 0
.nodeset V(sram[711]->outb) vsp
Xsram[712] sram->in sram[712]->out sram[712]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[712]->out) 0
.nodeset V(sram[712]->outb) vsp
Xsram[713] sram->in sram[713]->out sram[713]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[713]->out) 0
.nodeset V(sram[713]->outb) vsp
Xmux_2level_size50[4] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[0]->in[4] sram[714]->outb sram[714]->out sram[715]->out sram[715]->outb sram[716]->out sram[716]->outb sram[717]->out sram[717]->outb sram[718]->out sram[718]->outb sram[719]->out sram[719]->outb sram[720]->out sram[720]->outb sram[721]->out sram[721]->outb sram[722]->outb sram[722]->out sram[723]->out sram[723]->outb sram[724]->out sram[724]->outb sram[725]->out sram[725]->outb sram[726]->out sram[726]->outb sram[727]->out sram[727]->outb sram[728]->out sram[728]->outb sram[729]->out sram[729]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[4], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[714] sram->in sram[714]->out sram[714]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[714]->out) 0
.nodeset V(sram[714]->outb) vsp
Xsram[715] sram->in sram[715]->out sram[715]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[715]->out) 0
.nodeset V(sram[715]->outb) vsp
Xsram[716] sram->in sram[716]->out sram[716]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[716]->out) 0
.nodeset V(sram[716]->outb) vsp
Xsram[717] sram->in sram[717]->out sram[717]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[717]->out) 0
.nodeset V(sram[717]->outb) vsp
Xsram[718] sram->in sram[718]->out sram[718]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[718]->out) 0
.nodeset V(sram[718]->outb) vsp
Xsram[719] sram->in sram[719]->out sram[719]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[719]->out) 0
.nodeset V(sram[719]->outb) vsp
Xsram[720] sram->in sram[720]->out sram[720]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[720]->out) 0
.nodeset V(sram[720]->outb) vsp
Xsram[721] sram->in sram[721]->out sram[721]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[721]->out) 0
.nodeset V(sram[721]->outb) vsp
Xsram[722] sram->in sram[722]->out sram[722]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[722]->out) 0
.nodeset V(sram[722]->outb) vsp
Xsram[723] sram->in sram[723]->out sram[723]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[723]->out) 0
.nodeset V(sram[723]->outb) vsp
Xsram[724] sram->in sram[724]->out sram[724]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[724]->out) 0
.nodeset V(sram[724]->outb) vsp
Xsram[725] sram->in sram[725]->out sram[725]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[725]->out) 0
.nodeset V(sram[725]->outb) vsp
Xsram[726] sram->in sram[726]->out sram[726]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[726]->out) 0
.nodeset V(sram[726]->outb) vsp
Xsram[727] sram->in sram[727]->out sram[727]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[727]->out) 0
.nodeset V(sram[727]->outb) vsp
Xsram[728] sram->in sram[728]->out sram[728]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[728]->out) 0
.nodeset V(sram[728]->outb) vsp
Xsram[729] sram->in sram[729]->out sram[729]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[729]->out) 0
.nodeset V(sram[729]->outb) vsp
Xmux_2level_size50[5] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[0]->in[5] sram[730]->outb sram[730]->out sram[731]->out sram[731]->outb sram[732]->out sram[732]->outb sram[733]->out sram[733]->outb sram[734]->out sram[734]->outb sram[735]->out sram[735]->outb sram[736]->out sram[736]->outb sram[737]->out sram[737]->outb sram[738]->outb sram[738]->out sram[739]->out sram[739]->outb sram[740]->out sram[740]->outb sram[741]->out sram[741]->outb sram[742]->out sram[742]->outb sram[743]->out sram[743]->outb sram[744]->out sram[744]->outb sram[745]->out sram[745]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[5], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[730] sram->in sram[730]->out sram[730]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[730]->out) 0
.nodeset V(sram[730]->outb) vsp
Xsram[731] sram->in sram[731]->out sram[731]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[731]->out) 0
.nodeset V(sram[731]->outb) vsp
Xsram[732] sram->in sram[732]->out sram[732]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[732]->out) 0
.nodeset V(sram[732]->outb) vsp
Xsram[733] sram->in sram[733]->out sram[733]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[733]->out) 0
.nodeset V(sram[733]->outb) vsp
Xsram[734] sram->in sram[734]->out sram[734]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[734]->out) 0
.nodeset V(sram[734]->outb) vsp
Xsram[735] sram->in sram[735]->out sram[735]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[735]->out) 0
.nodeset V(sram[735]->outb) vsp
Xsram[736] sram->in sram[736]->out sram[736]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[736]->out) 0
.nodeset V(sram[736]->outb) vsp
Xsram[737] sram->in sram[737]->out sram[737]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[737]->out) 0
.nodeset V(sram[737]->outb) vsp
Xsram[738] sram->in sram[738]->out sram[738]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[738]->out) 0
.nodeset V(sram[738]->outb) vsp
Xsram[739] sram->in sram[739]->out sram[739]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[739]->out) 0
.nodeset V(sram[739]->outb) vsp
Xsram[740] sram->in sram[740]->out sram[740]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[740]->out) 0
.nodeset V(sram[740]->outb) vsp
Xsram[741] sram->in sram[741]->out sram[741]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[741]->out) 0
.nodeset V(sram[741]->outb) vsp
Xsram[742] sram->in sram[742]->out sram[742]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[742]->out) 0
.nodeset V(sram[742]->outb) vsp
Xsram[743] sram->in sram[743]->out sram[743]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[743]->out) 0
.nodeset V(sram[743]->outb) vsp
Xsram[744] sram->in sram[744]->out sram[744]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[744]->out) 0
.nodeset V(sram[744]->outb) vsp
Xsram[745] sram->in sram[745]->out sram[745]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[745]->out) 0
.nodeset V(sram[745]->outb) vsp
Xdirect_interc[170] mode[clb]->clk[0] fle[0]->clk[0] gvdd_local_interc sgnd direct_interc
Xmux_2level_size50[6] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[1]->in[0] sram[746]->outb sram[746]->out sram[747]->out sram[747]->outb sram[748]->out sram[748]->outb sram[749]->out sram[749]->outb sram[750]->out sram[750]->outb sram[751]->out sram[751]->outb sram[752]->out sram[752]->outb sram[753]->out sram[753]->outb sram[754]->outb sram[754]->out sram[755]->out sram[755]->outb sram[756]->out sram[756]->outb sram[757]->out sram[757]->outb sram[758]->out sram[758]->outb sram[759]->out sram[759]->outb sram[760]->out sram[760]->outb sram[761]->out sram[761]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[6], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[746] sram->in sram[746]->out sram[746]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[746]->out) 0
.nodeset V(sram[746]->outb) vsp
Xsram[747] sram->in sram[747]->out sram[747]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[747]->out) 0
.nodeset V(sram[747]->outb) vsp
Xsram[748] sram->in sram[748]->out sram[748]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[748]->out) 0
.nodeset V(sram[748]->outb) vsp
Xsram[749] sram->in sram[749]->out sram[749]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[749]->out) 0
.nodeset V(sram[749]->outb) vsp
Xsram[750] sram->in sram[750]->out sram[750]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[750]->out) 0
.nodeset V(sram[750]->outb) vsp
Xsram[751] sram->in sram[751]->out sram[751]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[751]->out) 0
.nodeset V(sram[751]->outb) vsp
Xsram[752] sram->in sram[752]->out sram[752]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[752]->out) 0
.nodeset V(sram[752]->outb) vsp
Xsram[753] sram->in sram[753]->out sram[753]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[753]->out) 0
.nodeset V(sram[753]->outb) vsp
Xsram[754] sram->in sram[754]->out sram[754]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[754]->out) 0
.nodeset V(sram[754]->outb) vsp
Xsram[755] sram->in sram[755]->out sram[755]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[755]->out) 0
.nodeset V(sram[755]->outb) vsp
Xsram[756] sram->in sram[756]->out sram[756]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[756]->out) 0
.nodeset V(sram[756]->outb) vsp
Xsram[757] sram->in sram[757]->out sram[757]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[757]->out) 0
.nodeset V(sram[757]->outb) vsp
Xsram[758] sram->in sram[758]->out sram[758]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[758]->out) 0
.nodeset V(sram[758]->outb) vsp
Xsram[759] sram->in sram[759]->out sram[759]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[759]->out) 0
.nodeset V(sram[759]->outb) vsp
Xsram[760] sram->in sram[760]->out sram[760]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[760]->out) 0
.nodeset V(sram[760]->outb) vsp
Xsram[761] sram->in sram[761]->out sram[761]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[761]->out) 0
.nodeset V(sram[761]->outb) vsp
Xmux_2level_size50[7] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[1]->in[1] sram[762]->outb sram[762]->out sram[763]->out sram[763]->outb sram[764]->out sram[764]->outb sram[765]->out sram[765]->outb sram[766]->out sram[766]->outb sram[767]->out sram[767]->outb sram[768]->out sram[768]->outb sram[769]->out sram[769]->outb sram[770]->outb sram[770]->out sram[771]->out sram[771]->outb sram[772]->out sram[772]->outb sram[773]->out sram[773]->outb sram[774]->out sram[774]->outb sram[775]->out sram[775]->outb sram[776]->out sram[776]->outb sram[777]->out sram[777]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[7], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[762] sram->in sram[762]->out sram[762]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[762]->out) 0
.nodeset V(sram[762]->outb) vsp
Xsram[763] sram->in sram[763]->out sram[763]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[763]->out) 0
.nodeset V(sram[763]->outb) vsp
Xsram[764] sram->in sram[764]->out sram[764]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[764]->out) 0
.nodeset V(sram[764]->outb) vsp
Xsram[765] sram->in sram[765]->out sram[765]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[765]->out) 0
.nodeset V(sram[765]->outb) vsp
Xsram[766] sram->in sram[766]->out sram[766]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[766]->out) 0
.nodeset V(sram[766]->outb) vsp
Xsram[767] sram->in sram[767]->out sram[767]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[767]->out) 0
.nodeset V(sram[767]->outb) vsp
Xsram[768] sram->in sram[768]->out sram[768]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[768]->out) 0
.nodeset V(sram[768]->outb) vsp
Xsram[769] sram->in sram[769]->out sram[769]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[769]->out) 0
.nodeset V(sram[769]->outb) vsp
Xsram[770] sram->in sram[770]->out sram[770]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[770]->out) 0
.nodeset V(sram[770]->outb) vsp
Xsram[771] sram->in sram[771]->out sram[771]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[771]->out) 0
.nodeset V(sram[771]->outb) vsp
Xsram[772] sram->in sram[772]->out sram[772]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[772]->out) 0
.nodeset V(sram[772]->outb) vsp
Xsram[773] sram->in sram[773]->out sram[773]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[773]->out) 0
.nodeset V(sram[773]->outb) vsp
Xsram[774] sram->in sram[774]->out sram[774]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[774]->out) 0
.nodeset V(sram[774]->outb) vsp
Xsram[775] sram->in sram[775]->out sram[775]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[775]->out) 0
.nodeset V(sram[775]->outb) vsp
Xsram[776] sram->in sram[776]->out sram[776]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[776]->out) 0
.nodeset V(sram[776]->outb) vsp
Xsram[777] sram->in sram[777]->out sram[777]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[777]->out) 0
.nodeset V(sram[777]->outb) vsp
Xmux_2level_size50[8] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[1]->in[2] sram[778]->outb sram[778]->out sram[779]->out sram[779]->outb sram[780]->out sram[780]->outb sram[781]->out sram[781]->outb sram[782]->out sram[782]->outb sram[783]->out sram[783]->outb sram[784]->out sram[784]->outb sram[785]->out sram[785]->outb sram[786]->outb sram[786]->out sram[787]->out sram[787]->outb sram[788]->out sram[788]->outb sram[789]->out sram[789]->outb sram[790]->out sram[790]->outb sram[791]->out sram[791]->outb sram[792]->out sram[792]->outb sram[793]->out sram[793]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[8], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[778] sram->in sram[778]->out sram[778]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[778]->out) 0
.nodeset V(sram[778]->outb) vsp
Xsram[779] sram->in sram[779]->out sram[779]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[779]->out) 0
.nodeset V(sram[779]->outb) vsp
Xsram[780] sram->in sram[780]->out sram[780]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[780]->out) 0
.nodeset V(sram[780]->outb) vsp
Xsram[781] sram->in sram[781]->out sram[781]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[781]->out) 0
.nodeset V(sram[781]->outb) vsp
Xsram[782] sram->in sram[782]->out sram[782]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[782]->out) 0
.nodeset V(sram[782]->outb) vsp
Xsram[783] sram->in sram[783]->out sram[783]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[783]->out) 0
.nodeset V(sram[783]->outb) vsp
Xsram[784] sram->in sram[784]->out sram[784]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[784]->out) 0
.nodeset V(sram[784]->outb) vsp
Xsram[785] sram->in sram[785]->out sram[785]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[785]->out) 0
.nodeset V(sram[785]->outb) vsp
Xsram[786] sram->in sram[786]->out sram[786]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[786]->out) 0
.nodeset V(sram[786]->outb) vsp
Xsram[787] sram->in sram[787]->out sram[787]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[787]->out) 0
.nodeset V(sram[787]->outb) vsp
Xsram[788] sram->in sram[788]->out sram[788]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[788]->out) 0
.nodeset V(sram[788]->outb) vsp
Xsram[789] sram->in sram[789]->out sram[789]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[789]->out) 0
.nodeset V(sram[789]->outb) vsp
Xsram[790] sram->in sram[790]->out sram[790]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[790]->out) 0
.nodeset V(sram[790]->outb) vsp
Xsram[791] sram->in sram[791]->out sram[791]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[791]->out) 0
.nodeset V(sram[791]->outb) vsp
Xsram[792] sram->in sram[792]->out sram[792]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[792]->out) 0
.nodeset V(sram[792]->outb) vsp
Xsram[793] sram->in sram[793]->out sram[793]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[793]->out) 0
.nodeset V(sram[793]->outb) vsp
Xmux_2level_size50[9] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[1]->in[3] sram[794]->outb sram[794]->out sram[795]->out sram[795]->outb sram[796]->out sram[796]->outb sram[797]->out sram[797]->outb sram[798]->out sram[798]->outb sram[799]->out sram[799]->outb sram[800]->out sram[800]->outb sram[801]->out sram[801]->outb sram[802]->outb sram[802]->out sram[803]->out sram[803]->outb sram[804]->out sram[804]->outb sram[805]->out sram[805]->outb sram[806]->out sram[806]->outb sram[807]->out sram[807]->outb sram[808]->out sram[808]->outb sram[809]->out sram[809]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[9], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[794] sram->in sram[794]->out sram[794]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[794]->out) 0
.nodeset V(sram[794]->outb) vsp
Xsram[795] sram->in sram[795]->out sram[795]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[795]->out) 0
.nodeset V(sram[795]->outb) vsp
Xsram[796] sram->in sram[796]->out sram[796]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[796]->out) 0
.nodeset V(sram[796]->outb) vsp
Xsram[797] sram->in sram[797]->out sram[797]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[797]->out) 0
.nodeset V(sram[797]->outb) vsp
Xsram[798] sram->in sram[798]->out sram[798]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[798]->out) 0
.nodeset V(sram[798]->outb) vsp
Xsram[799] sram->in sram[799]->out sram[799]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[799]->out) 0
.nodeset V(sram[799]->outb) vsp
Xsram[800] sram->in sram[800]->out sram[800]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[800]->out) 0
.nodeset V(sram[800]->outb) vsp
Xsram[801] sram->in sram[801]->out sram[801]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[801]->out) 0
.nodeset V(sram[801]->outb) vsp
Xsram[802] sram->in sram[802]->out sram[802]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[802]->out) 0
.nodeset V(sram[802]->outb) vsp
Xsram[803] sram->in sram[803]->out sram[803]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[803]->out) 0
.nodeset V(sram[803]->outb) vsp
Xsram[804] sram->in sram[804]->out sram[804]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[804]->out) 0
.nodeset V(sram[804]->outb) vsp
Xsram[805] sram->in sram[805]->out sram[805]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[805]->out) 0
.nodeset V(sram[805]->outb) vsp
Xsram[806] sram->in sram[806]->out sram[806]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[806]->out) 0
.nodeset V(sram[806]->outb) vsp
Xsram[807] sram->in sram[807]->out sram[807]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[807]->out) 0
.nodeset V(sram[807]->outb) vsp
Xsram[808] sram->in sram[808]->out sram[808]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[808]->out) 0
.nodeset V(sram[808]->outb) vsp
Xsram[809] sram->in sram[809]->out sram[809]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[809]->out) 0
.nodeset V(sram[809]->outb) vsp
Xmux_2level_size50[10] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[1]->in[4] sram[810]->outb sram[810]->out sram[811]->out sram[811]->outb sram[812]->out sram[812]->outb sram[813]->out sram[813]->outb sram[814]->out sram[814]->outb sram[815]->out sram[815]->outb sram[816]->out sram[816]->outb sram[817]->out sram[817]->outb sram[818]->outb sram[818]->out sram[819]->out sram[819]->outb sram[820]->out sram[820]->outb sram[821]->out sram[821]->outb sram[822]->out sram[822]->outb sram[823]->out sram[823]->outb sram[824]->out sram[824]->outb sram[825]->out sram[825]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[10], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[810] sram->in sram[810]->out sram[810]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[810]->out) 0
.nodeset V(sram[810]->outb) vsp
Xsram[811] sram->in sram[811]->out sram[811]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[811]->out) 0
.nodeset V(sram[811]->outb) vsp
Xsram[812] sram->in sram[812]->out sram[812]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[812]->out) 0
.nodeset V(sram[812]->outb) vsp
Xsram[813] sram->in sram[813]->out sram[813]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[813]->out) 0
.nodeset V(sram[813]->outb) vsp
Xsram[814] sram->in sram[814]->out sram[814]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[814]->out) 0
.nodeset V(sram[814]->outb) vsp
Xsram[815] sram->in sram[815]->out sram[815]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[815]->out) 0
.nodeset V(sram[815]->outb) vsp
Xsram[816] sram->in sram[816]->out sram[816]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[816]->out) 0
.nodeset V(sram[816]->outb) vsp
Xsram[817] sram->in sram[817]->out sram[817]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[817]->out) 0
.nodeset V(sram[817]->outb) vsp
Xsram[818] sram->in sram[818]->out sram[818]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[818]->out) 0
.nodeset V(sram[818]->outb) vsp
Xsram[819] sram->in sram[819]->out sram[819]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[819]->out) 0
.nodeset V(sram[819]->outb) vsp
Xsram[820] sram->in sram[820]->out sram[820]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[820]->out) 0
.nodeset V(sram[820]->outb) vsp
Xsram[821] sram->in sram[821]->out sram[821]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[821]->out) 0
.nodeset V(sram[821]->outb) vsp
Xsram[822] sram->in sram[822]->out sram[822]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[822]->out) 0
.nodeset V(sram[822]->outb) vsp
Xsram[823] sram->in sram[823]->out sram[823]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[823]->out) 0
.nodeset V(sram[823]->outb) vsp
Xsram[824] sram->in sram[824]->out sram[824]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[824]->out) 0
.nodeset V(sram[824]->outb) vsp
Xsram[825] sram->in sram[825]->out sram[825]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[825]->out) 0
.nodeset V(sram[825]->outb) vsp
Xmux_2level_size50[11] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[1]->in[5] sram[826]->outb sram[826]->out sram[827]->out sram[827]->outb sram[828]->out sram[828]->outb sram[829]->out sram[829]->outb sram[830]->out sram[830]->outb sram[831]->out sram[831]->outb sram[832]->out sram[832]->outb sram[833]->out sram[833]->outb sram[834]->outb sram[834]->out sram[835]->out sram[835]->outb sram[836]->out sram[836]->outb sram[837]->out sram[837]->outb sram[838]->out sram[838]->outb sram[839]->out sram[839]->outb sram[840]->out sram[840]->outb sram[841]->out sram[841]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[11], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[826] sram->in sram[826]->out sram[826]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[826]->out) 0
.nodeset V(sram[826]->outb) vsp
Xsram[827] sram->in sram[827]->out sram[827]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[827]->out) 0
.nodeset V(sram[827]->outb) vsp
Xsram[828] sram->in sram[828]->out sram[828]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[828]->out) 0
.nodeset V(sram[828]->outb) vsp
Xsram[829] sram->in sram[829]->out sram[829]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[829]->out) 0
.nodeset V(sram[829]->outb) vsp
Xsram[830] sram->in sram[830]->out sram[830]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[830]->out) 0
.nodeset V(sram[830]->outb) vsp
Xsram[831] sram->in sram[831]->out sram[831]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[831]->out) 0
.nodeset V(sram[831]->outb) vsp
Xsram[832] sram->in sram[832]->out sram[832]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[832]->out) 0
.nodeset V(sram[832]->outb) vsp
Xsram[833] sram->in sram[833]->out sram[833]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[833]->out) 0
.nodeset V(sram[833]->outb) vsp
Xsram[834] sram->in sram[834]->out sram[834]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[834]->out) 0
.nodeset V(sram[834]->outb) vsp
Xsram[835] sram->in sram[835]->out sram[835]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[835]->out) 0
.nodeset V(sram[835]->outb) vsp
Xsram[836] sram->in sram[836]->out sram[836]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[836]->out) 0
.nodeset V(sram[836]->outb) vsp
Xsram[837] sram->in sram[837]->out sram[837]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[837]->out) 0
.nodeset V(sram[837]->outb) vsp
Xsram[838] sram->in sram[838]->out sram[838]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[838]->out) 0
.nodeset V(sram[838]->outb) vsp
Xsram[839] sram->in sram[839]->out sram[839]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[839]->out) 0
.nodeset V(sram[839]->outb) vsp
Xsram[840] sram->in sram[840]->out sram[840]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[840]->out) 0
.nodeset V(sram[840]->outb) vsp
Xsram[841] sram->in sram[841]->out sram[841]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[841]->out) 0
.nodeset V(sram[841]->outb) vsp
Xdirect_interc[171] mode[clb]->clk[0] fle[1]->clk[0] gvdd_local_interc sgnd direct_interc
Xmux_2level_size50[12] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[2]->in[0] sram[842]->outb sram[842]->out sram[843]->out sram[843]->outb sram[844]->out sram[844]->outb sram[845]->out sram[845]->outb sram[846]->out sram[846]->outb sram[847]->out sram[847]->outb sram[848]->out sram[848]->outb sram[849]->out sram[849]->outb sram[850]->outb sram[850]->out sram[851]->out sram[851]->outb sram[852]->out sram[852]->outb sram[853]->out sram[853]->outb sram[854]->out sram[854]->outb sram[855]->out sram[855]->outb sram[856]->out sram[856]->outb sram[857]->out sram[857]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[12], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[842] sram->in sram[842]->out sram[842]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[842]->out) 0
.nodeset V(sram[842]->outb) vsp
Xsram[843] sram->in sram[843]->out sram[843]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[843]->out) 0
.nodeset V(sram[843]->outb) vsp
Xsram[844] sram->in sram[844]->out sram[844]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[844]->out) 0
.nodeset V(sram[844]->outb) vsp
Xsram[845] sram->in sram[845]->out sram[845]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[845]->out) 0
.nodeset V(sram[845]->outb) vsp
Xsram[846] sram->in sram[846]->out sram[846]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[846]->out) 0
.nodeset V(sram[846]->outb) vsp
Xsram[847] sram->in sram[847]->out sram[847]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[847]->out) 0
.nodeset V(sram[847]->outb) vsp
Xsram[848] sram->in sram[848]->out sram[848]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[848]->out) 0
.nodeset V(sram[848]->outb) vsp
Xsram[849] sram->in sram[849]->out sram[849]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[849]->out) 0
.nodeset V(sram[849]->outb) vsp
Xsram[850] sram->in sram[850]->out sram[850]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[850]->out) 0
.nodeset V(sram[850]->outb) vsp
Xsram[851] sram->in sram[851]->out sram[851]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[851]->out) 0
.nodeset V(sram[851]->outb) vsp
Xsram[852] sram->in sram[852]->out sram[852]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[852]->out) 0
.nodeset V(sram[852]->outb) vsp
Xsram[853] sram->in sram[853]->out sram[853]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[853]->out) 0
.nodeset V(sram[853]->outb) vsp
Xsram[854] sram->in sram[854]->out sram[854]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[854]->out) 0
.nodeset V(sram[854]->outb) vsp
Xsram[855] sram->in sram[855]->out sram[855]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[855]->out) 0
.nodeset V(sram[855]->outb) vsp
Xsram[856] sram->in sram[856]->out sram[856]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[856]->out) 0
.nodeset V(sram[856]->outb) vsp
Xsram[857] sram->in sram[857]->out sram[857]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[857]->out) 0
.nodeset V(sram[857]->outb) vsp
Xmux_2level_size50[13] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[2]->in[1] sram[858]->outb sram[858]->out sram[859]->out sram[859]->outb sram[860]->out sram[860]->outb sram[861]->out sram[861]->outb sram[862]->out sram[862]->outb sram[863]->out sram[863]->outb sram[864]->out sram[864]->outb sram[865]->out sram[865]->outb sram[866]->outb sram[866]->out sram[867]->out sram[867]->outb sram[868]->out sram[868]->outb sram[869]->out sram[869]->outb sram[870]->out sram[870]->outb sram[871]->out sram[871]->outb sram[872]->out sram[872]->outb sram[873]->out sram[873]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[13], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[858] sram->in sram[858]->out sram[858]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[858]->out) 0
.nodeset V(sram[858]->outb) vsp
Xsram[859] sram->in sram[859]->out sram[859]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[859]->out) 0
.nodeset V(sram[859]->outb) vsp
Xsram[860] sram->in sram[860]->out sram[860]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[860]->out) 0
.nodeset V(sram[860]->outb) vsp
Xsram[861] sram->in sram[861]->out sram[861]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[861]->out) 0
.nodeset V(sram[861]->outb) vsp
Xsram[862] sram->in sram[862]->out sram[862]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[862]->out) 0
.nodeset V(sram[862]->outb) vsp
Xsram[863] sram->in sram[863]->out sram[863]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[863]->out) 0
.nodeset V(sram[863]->outb) vsp
Xsram[864] sram->in sram[864]->out sram[864]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[864]->out) 0
.nodeset V(sram[864]->outb) vsp
Xsram[865] sram->in sram[865]->out sram[865]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[865]->out) 0
.nodeset V(sram[865]->outb) vsp
Xsram[866] sram->in sram[866]->out sram[866]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[866]->out) 0
.nodeset V(sram[866]->outb) vsp
Xsram[867] sram->in sram[867]->out sram[867]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[867]->out) 0
.nodeset V(sram[867]->outb) vsp
Xsram[868] sram->in sram[868]->out sram[868]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[868]->out) 0
.nodeset V(sram[868]->outb) vsp
Xsram[869] sram->in sram[869]->out sram[869]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[869]->out) 0
.nodeset V(sram[869]->outb) vsp
Xsram[870] sram->in sram[870]->out sram[870]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[870]->out) 0
.nodeset V(sram[870]->outb) vsp
Xsram[871] sram->in sram[871]->out sram[871]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[871]->out) 0
.nodeset V(sram[871]->outb) vsp
Xsram[872] sram->in sram[872]->out sram[872]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[872]->out) 0
.nodeset V(sram[872]->outb) vsp
Xsram[873] sram->in sram[873]->out sram[873]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[873]->out) 0
.nodeset V(sram[873]->outb) vsp
Xmux_2level_size50[14] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[2]->in[2] sram[874]->outb sram[874]->out sram[875]->out sram[875]->outb sram[876]->out sram[876]->outb sram[877]->out sram[877]->outb sram[878]->out sram[878]->outb sram[879]->out sram[879]->outb sram[880]->out sram[880]->outb sram[881]->out sram[881]->outb sram[882]->outb sram[882]->out sram[883]->out sram[883]->outb sram[884]->out sram[884]->outb sram[885]->out sram[885]->outb sram[886]->out sram[886]->outb sram[887]->out sram[887]->outb sram[888]->out sram[888]->outb sram[889]->out sram[889]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[14], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[874] sram->in sram[874]->out sram[874]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[874]->out) 0
.nodeset V(sram[874]->outb) vsp
Xsram[875] sram->in sram[875]->out sram[875]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[875]->out) 0
.nodeset V(sram[875]->outb) vsp
Xsram[876] sram->in sram[876]->out sram[876]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[876]->out) 0
.nodeset V(sram[876]->outb) vsp
Xsram[877] sram->in sram[877]->out sram[877]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[877]->out) 0
.nodeset V(sram[877]->outb) vsp
Xsram[878] sram->in sram[878]->out sram[878]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[878]->out) 0
.nodeset V(sram[878]->outb) vsp
Xsram[879] sram->in sram[879]->out sram[879]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[879]->out) 0
.nodeset V(sram[879]->outb) vsp
Xsram[880] sram->in sram[880]->out sram[880]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[880]->out) 0
.nodeset V(sram[880]->outb) vsp
Xsram[881] sram->in sram[881]->out sram[881]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[881]->out) 0
.nodeset V(sram[881]->outb) vsp
Xsram[882] sram->in sram[882]->out sram[882]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[882]->out) 0
.nodeset V(sram[882]->outb) vsp
Xsram[883] sram->in sram[883]->out sram[883]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[883]->out) 0
.nodeset V(sram[883]->outb) vsp
Xsram[884] sram->in sram[884]->out sram[884]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[884]->out) 0
.nodeset V(sram[884]->outb) vsp
Xsram[885] sram->in sram[885]->out sram[885]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[885]->out) 0
.nodeset V(sram[885]->outb) vsp
Xsram[886] sram->in sram[886]->out sram[886]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[886]->out) 0
.nodeset V(sram[886]->outb) vsp
Xsram[887] sram->in sram[887]->out sram[887]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[887]->out) 0
.nodeset V(sram[887]->outb) vsp
Xsram[888] sram->in sram[888]->out sram[888]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[888]->out) 0
.nodeset V(sram[888]->outb) vsp
Xsram[889] sram->in sram[889]->out sram[889]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[889]->out) 0
.nodeset V(sram[889]->outb) vsp
Xmux_2level_size50[15] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[2]->in[3] sram[890]->outb sram[890]->out sram[891]->out sram[891]->outb sram[892]->out sram[892]->outb sram[893]->out sram[893]->outb sram[894]->out sram[894]->outb sram[895]->out sram[895]->outb sram[896]->out sram[896]->outb sram[897]->out sram[897]->outb sram[898]->outb sram[898]->out sram[899]->out sram[899]->outb sram[900]->out sram[900]->outb sram[901]->out sram[901]->outb sram[902]->out sram[902]->outb sram[903]->out sram[903]->outb sram[904]->out sram[904]->outb sram[905]->out sram[905]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[15], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[890] sram->in sram[890]->out sram[890]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[890]->out) 0
.nodeset V(sram[890]->outb) vsp
Xsram[891] sram->in sram[891]->out sram[891]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[891]->out) 0
.nodeset V(sram[891]->outb) vsp
Xsram[892] sram->in sram[892]->out sram[892]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[892]->out) 0
.nodeset V(sram[892]->outb) vsp
Xsram[893] sram->in sram[893]->out sram[893]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[893]->out) 0
.nodeset V(sram[893]->outb) vsp
Xsram[894] sram->in sram[894]->out sram[894]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[894]->out) 0
.nodeset V(sram[894]->outb) vsp
Xsram[895] sram->in sram[895]->out sram[895]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[895]->out) 0
.nodeset V(sram[895]->outb) vsp
Xsram[896] sram->in sram[896]->out sram[896]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[896]->out) 0
.nodeset V(sram[896]->outb) vsp
Xsram[897] sram->in sram[897]->out sram[897]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[897]->out) 0
.nodeset V(sram[897]->outb) vsp
Xsram[898] sram->in sram[898]->out sram[898]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[898]->out) 0
.nodeset V(sram[898]->outb) vsp
Xsram[899] sram->in sram[899]->out sram[899]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[899]->out) 0
.nodeset V(sram[899]->outb) vsp
Xsram[900] sram->in sram[900]->out sram[900]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[900]->out) 0
.nodeset V(sram[900]->outb) vsp
Xsram[901] sram->in sram[901]->out sram[901]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[901]->out) 0
.nodeset V(sram[901]->outb) vsp
Xsram[902] sram->in sram[902]->out sram[902]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[902]->out) 0
.nodeset V(sram[902]->outb) vsp
Xsram[903] sram->in sram[903]->out sram[903]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[903]->out) 0
.nodeset V(sram[903]->outb) vsp
Xsram[904] sram->in sram[904]->out sram[904]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[904]->out) 0
.nodeset V(sram[904]->outb) vsp
Xsram[905] sram->in sram[905]->out sram[905]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[905]->out) 0
.nodeset V(sram[905]->outb) vsp
Xmux_2level_size50[16] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[2]->in[4] sram[906]->outb sram[906]->out sram[907]->out sram[907]->outb sram[908]->out sram[908]->outb sram[909]->out sram[909]->outb sram[910]->out sram[910]->outb sram[911]->out sram[911]->outb sram[912]->out sram[912]->outb sram[913]->out sram[913]->outb sram[914]->outb sram[914]->out sram[915]->out sram[915]->outb sram[916]->out sram[916]->outb sram[917]->out sram[917]->outb sram[918]->out sram[918]->outb sram[919]->out sram[919]->outb sram[920]->out sram[920]->outb sram[921]->out sram[921]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[16], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[906] sram->in sram[906]->out sram[906]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[906]->out) 0
.nodeset V(sram[906]->outb) vsp
Xsram[907] sram->in sram[907]->out sram[907]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[907]->out) 0
.nodeset V(sram[907]->outb) vsp
Xsram[908] sram->in sram[908]->out sram[908]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[908]->out) 0
.nodeset V(sram[908]->outb) vsp
Xsram[909] sram->in sram[909]->out sram[909]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[909]->out) 0
.nodeset V(sram[909]->outb) vsp
Xsram[910] sram->in sram[910]->out sram[910]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[910]->out) 0
.nodeset V(sram[910]->outb) vsp
Xsram[911] sram->in sram[911]->out sram[911]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[911]->out) 0
.nodeset V(sram[911]->outb) vsp
Xsram[912] sram->in sram[912]->out sram[912]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[912]->out) 0
.nodeset V(sram[912]->outb) vsp
Xsram[913] sram->in sram[913]->out sram[913]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[913]->out) 0
.nodeset V(sram[913]->outb) vsp
Xsram[914] sram->in sram[914]->out sram[914]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[914]->out) 0
.nodeset V(sram[914]->outb) vsp
Xsram[915] sram->in sram[915]->out sram[915]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[915]->out) 0
.nodeset V(sram[915]->outb) vsp
Xsram[916] sram->in sram[916]->out sram[916]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[916]->out) 0
.nodeset V(sram[916]->outb) vsp
Xsram[917] sram->in sram[917]->out sram[917]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[917]->out) 0
.nodeset V(sram[917]->outb) vsp
Xsram[918] sram->in sram[918]->out sram[918]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[918]->out) 0
.nodeset V(sram[918]->outb) vsp
Xsram[919] sram->in sram[919]->out sram[919]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[919]->out) 0
.nodeset V(sram[919]->outb) vsp
Xsram[920] sram->in sram[920]->out sram[920]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[920]->out) 0
.nodeset V(sram[920]->outb) vsp
Xsram[921] sram->in sram[921]->out sram[921]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[921]->out) 0
.nodeset V(sram[921]->outb) vsp
Xmux_2level_size50[17] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[2]->in[5] sram[922]->outb sram[922]->out sram[923]->out sram[923]->outb sram[924]->out sram[924]->outb sram[925]->out sram[925]->outb sram[926]->out sram[926]->outb sram[927]->out sram[927]->outb sram[928]->out sram[928]->outb sram[929]->out sram[929]->outb sram[930]->outb sram[930]->out sram[931]->out sram[931]->outb sram[932]->out sram[932]->outb sram[933]->out sram[933]->outb sram[934]->out sram[934]->outb sram[935]->out sram[935]->outb sram[936]->out sram[936]->outb sram[937]->out sram[937]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[17], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[922] sram->in sram[922]->out sram[922]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[922]->out) 0
.nodeset V(sram[922]->outb) vsp
Xsram[923] sram->in sram[923]->out sram[923]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[923]->out) 0
.nodeset V(sram[923]->outb) vsp
Xsram[924] sram->in sram[924]->out sram[924]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[924]->out) 0
.nodeset V(sram[924]->outb) vsp
Xsram[925] sram->in sram[925]->out sram[925]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[925]->out) 0
.nodeset V(sram[925]->outb) vsp
Xsram[926] sram->in sram[926]->out sram[926]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[926]->out) 0
.nodeset V(sram[926]->outb) vsp
Xsram[927] sram->in sram[927]->out sram[927]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[927]->out) 0
.nodeset V(sram[927]->outb) vsp
Xsram[928] sram->in sram[928]->out sram[928]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[928]->out) 0
.nodeset V(sram[928]->outb) vsp
Xsram[929] sram->in sram[929]->out sram[929]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[929]->out) 0
.nodeset V(sram[929]->outb) vsp
Xsram[930] sram->in sram[930]->out sram[930]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[930]->out) 0
.nodeset V(sram[930]->outb) vsp
Xsram[931] sram->in sram[931]->out sram[931]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[931]->out) 0
.nodeset V(sram[931]->outb) vsp
Xsram[932] sram->in sram[932]->out sram[932]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[932]->out) 0
.nodeset V(sram[932]->outb) vsp
Xsram[933] sram->in sram[933]->out sram[933]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[933]->out) 0
.nodeset V(sram[933]->outb) vsp
Xsram[934] sram->in sram[934]->out sram[934]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[934]->out) 0
.nodeset V(sram[934]->outb) vsp
Xsram[935] sram->in sram[935]->out sram[935]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[935]->out) 0
.nodeset V(sram[935]->outb) vsp
Xsram[936] sram->in sram[936]->out sram[936]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[936]->out) 0
.nodeset V(sram[936]->outb) vsp
Xsram[937] sram->in sram[937]->out sram[937]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[937]->out) 0
.nodeset V(sram[937]->outb) vsp
Xdirect_interc[172] mode[clb]->clk[0] fle[2]->clk[0] gvdd_local_interc sgnd direct_interc
Xmux_2level_size50[18] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[3]->in[0] sram[938]->outb sram[938]->out sram[939]->out sram[939]->outb sram[940]->out sram[940]->outb sram[941]->out sram[941]->outb sram[942]->out sram[942]->outb sram[943]->out sram[943]->outb sram[944]->out sram[944]->outb sram[945]->out sram[945]->outb sram[946]->outb sram[946]->out sram[947]->out sram[947]->outb sram[948]->out sram[948]->outb sram[949]->out sram[949]->outb sram[950]->out sram[950]->outb sram[951]->out sram[951]->outb sram[952]->out sram[952]->outb sram[953]->out sram[953]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[18], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[938] sram->in sram[938]->out sram[938]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[938]->out) 0
.nodeset V(sram[938]->outb) vsp
Xsram[939] sram->in sram[939]->out sram[939]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[939]->out) 0
.nodeset V(sram[939]->outb) vsp
Xsram[940] sram->in sram[940]->out sram[940]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[940]->out) 0
.nodeset V(sram[940]->outb) vsp
Xsram[941] sram->in sram[941]->out sram[941]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[941]->out) 0
.nodeset V(sram[941]->outb) vsp
Xsram[942] sram->in sram[942]->out sram[942]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[942]->out) 0
.nodeset V(sram[942]->outb) vsp
Xsram[943] sram->in sram[943]->out sram[943]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[943]->out) 0
.nodeset V(sram[943]->outb) vsp
Xsram[944] sram->in sram[944]->out sram[944]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[944]->out) 0
.nodeset V(sram[944]->outb) vsp
Xsram[945] sram->in sram[945]->out sram[945]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[945]->out) 0
.nodeset V(sram[945]->outb) vsp
Xsram[946] sram->in sram[946]->out sram[946]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[946]->out) 0
.nodeset V(sram[946]->outb) vsp
Xsram[947] sram->in sram[947]->out sram[947]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[947]->out) 0
.nodeset V(sram[947]->outb) vsp
Xsram[948] sram->in sram[948]->out sram[948]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[948]->out) 0
.nodeset V(sram[948]->outb) vsp
Xsram[949] sram->in sram[949]->out sram[949]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[949]->out) 0
.nodeset V(sram[949]->outb) vsp
Xsram[950] sram->in sram[950]->out sram[950]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[950]->out) 0
.nodeset V(sram[950]->outb) vsp
Xsram[951] sram->in sram[951]->out sram[951]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[951]->out) 0
.nodeset V(sram[951]->outb) vsp
Xsram[952] sram->in sram[952]->out sram[952]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[952]->out) 0
.nodeset V(sram[952]->outb) vsp
Xsram[953] sram->in sram[953]->out sram[953]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[953]->out) 0
.nodeset V(sram[953]->outb) vsp
Xmux_2level_size50[19] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[3]->in[1] sram[954]->outb sram[954]->out sram[955]->out sram[955]->outb sram[956]->out sram[956]->outb sram[957]->out sram[957]->outb sram[958]->out sram[958]->outb sram[959]->out sram[959]->outb sram[960]->out sram[960]->outb sram[961]->out sram[961]->outb sram[962]->outb sram[962]->out sram[963]->out sram[963]->outb sram[964]->out sram[964]->outb sram[965]->out sram[965]->outb sram[966]->out sram[966]->outb sram[967]->out sram[967]->outb sram[968]->out sram[968]->outb sram[969]->out sram[969]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[19], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[954] sram->in sram[954]->out sram[954]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[954]->out) 0
.nodeset V(sram[954]->outb) vsp
Xsram[955] sram->in sram[955]->out sram[955]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[955]->out) 0
.nodeset V(sram[955]->outb) vsp
Xsram[956] sram->in sram[956]->out sram[956]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[956]->out) 0
.nodeset V(sram[956]->outb) vsp
Xsram[957] sram->in sram[957]->out sram[957]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[957]->out) 0
.nodeset V(sram[957]->outb) vsp
Xsram[958] sram->in sram[958]->out sram[958]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[958]->out) 0
.nodeset V(sram[958]->outb) vsp
Xsram[959] sram->in sram[959]->out sram[959]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[959]->out) 0
.nodeset V(sram[959]->outb) vsp
Xsram[960] sram->in sram[960]->out sram[960]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[960]->out) 0
.nodeset V(sram[960]->outb) vsp
Xsram[961] sram->in sram[961]->out sram[961]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[961]->out) 0
.nodeset V(sram[961]->outb) vsp
Xsram[962] sram->in sram[962]->out sram[962]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[962]->out) 0
.nodeset V(sram[962]->outb) vsp
Xsram[963] sram->in sram[963]->out sram[963]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[963]->out) 0
.nodeset V(sram[963]->outb) vsp
Xsram[964] sram->in sram[964]->out sram[964]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[964]->out) 0
.nodeset V(sram[964]->outb) vsp
Xsram[965] sram->in sram[965]->out sram[965]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[965]->out) 0
.nodeset V(sram[965]->outb) vsp
Xsram[966] sram->in sram[966]->out sram[966]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[966]->out) 0
.nodeset V(sram[966]->outb) vsp
Xsram[967] sram->in sram[967]->out sram[967]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[967]->out) 0
.nodeset V(sram[967]->outb) vsp
Xsram[968] sram->in sram[968]->out sram[968]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[968]->out) 0
.nodeset V(sram[968]->outb) vsp
Xsram[969] sram->in sram[969]->out sram[969]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[969]->out) 0
.nodeset V(sram[969]->outb) vsp
Xmux_2level_size50[20] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[3]->in[2] sram[970]->outb sram[970]->out sram[971]->out sram[971]->outb sram[972]->out sram[972]->outb sram[973]->out sram[973]->outb sram[974]->out sram[974]->outb sram[975]->out sram[975]->outb sram[976]->out sram[976]->outb sram[977]->out sram[977]->outb sram[978]->outb sram[978]->out sram[979]->out sram[979]->outb sram[980]->out sram[980]->outb sram[981]->out sram[981]->outb sram[982]->out sram[982]->outb sram[983]->out sram[983]->outb sram[984]->out sram[984]->outb sram[985]->out sram[985]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[20], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[970] sram->in sram[970]->out sram[970]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[970]->out) 0
.nodeset V(sram[970]->outb) vsp
Xsram[971] sram->in sram[971]->out sram[971]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[971]->out) 0
.nodeset V(sram[971]->outb) vsp
Xsram[972] sram->in sram[972]->out sram[972]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[972]->out) 0
.nodeset V(sram[972]->outb) vsp
Xsram[973] sram->in sram[973]->out sram[973]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[973]->out) 0
.nodeset V(sram[973]->outb) vsp
Xsram[974] sram->in sram[974]->out sram[974]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[974]->out) 0
.nodeset V(sram[974]->outb) vsp
Xsram[975] sram->in sram[975]->out sram[975]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[975]->out) 0
.nodeset V(sram[975]->outb) vsp
Xsram[976] sram->in sram[976]->out sram[976]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[976]->out) 0
.nodeset V(sram[976]->outb) vsp
Xsram[977] sram->in sram[977]->out sram[977]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[977]->out) 0
.nodeset V(sram[977]->outb) vsp
Xsram[978] sram->in sram[978]->out sram[978]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[978]->out) 0
.nodeset V(sram[978]->outb) vsp
Xsram[979] sram->in sram[979]->out sram[979]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[979]->out) 0
.nodeset V(sram[979]->outb) vsp
Xsram[980] sram->in sram[980]->out sram[980]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[980]->out) 0
.nodeset V(sram[980]->outb) vsp
Xsram[981] sram->in sram[981]->out sram[981]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[981]->out) 0
.nodeset V(sram[981]->outb) vsp
Xsram[982] sram->in sram[982]->out sram[982]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[982]->out) 0
.nodeset V(sram[982]->outb) vsp
Xsram[983] sram->in sram[983]->out sram[983]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[983]->out) 0
.nodeset V(sram[983]->outb) vsp
Xsram[984] sram->in sram[984]->out sram[984]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[984]->out) 0
.nodeset V(sram[984]->outb) vsp
Xsram[985] sram->in sram[985]->out sram[985]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[985]->out) 0
.nodeset V(sram[985]->outb) vsp
Xmux_2level_size50[21] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[3]->in[3] sram[986]->outb sram[986]->out sram[987]->out sram[987]->outb sram[988]->out sram[988]->outb sram[989]->out sram[989]->outb sram[990]->out sram[990]->outb sram[991]->out sram[991]->outb sram[992]->out sram[992]->outb sram[993]->out sram[993]->outb sram[994]->outb sram[994]->out sram[995]->out sram[995]->outb sram[996]->out sram[996]->outb sram[997]->out sram[997]->outb sram[998]->out sram[998]->outb sram[999]->out sram[999]->outb sram[1000]->out sram[1000]->outb sram[1001]->out sram[1001]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[21], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[986] sram->in sram[986]->out sram[986]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[986]->out) 0
.nodeset V(sram[986]->outb) vsp
Xsram[987] sram->in sram[987]->out sram[987]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[987]->out) 0
.nodeset V(sram[987]->outb) vsp
Xsram[988] sram->in sram[988]->out sram[988]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[988]->out) 0
.nodeset V(sram[988]->outb) vsp
Xsram[989] sram->in sram[989]->out sram[989]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[989]->out) 0
.nodeset V(sram[989]->outb) vsp
Xsram[990] sram->in sram[990]->out sram[990]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[990]->out) 0
.nodeset V(sram[990]->outb) vsp
Xsram[991] sram->in sram[991]->out sram[991]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[991]->out) 0
.nodeset V(sram[991]->outb) vsp
Xsram[992] sram->in sram[992]->out sram[992]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[992]->out) 0
.nodeset V(sram[992]->outb) vsp
Xsram[993] sram->in sram[993]->out sram[993]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[993]->out) 0
.nodeset V(sram[993]->outb) vsp
Xsram[994] sram->in sram[994]->out sram[994]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[994]->out) 0
.nodeset V(sram[994]->outb) vsp
Xsram[995] sram->in sram[995]->out sram[995]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[995]->out) 0
.nodeset V(sram[995]->outb) vsp
Xsram[996] sram->in sram[996]->out sram[996]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[996]->out) 0
.nodeset V(sram[996]->outb) vsp
Xsram[997] sram->in sram[997]->out sram[997]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[997]->out) 0
.nodeset V(sram[997]->outb) vsp
Xsram[998] sram->in sram[998]->out sram[998]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[998]->out) 0
.nodeset V(sram[998]->outb) vsp
Xsram[999] sram->in sram[999]->out sram[999]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[999]->out) 0
.nodeset V(sram[999]->outb) vsp
Xsram[1000] sram->in sram[1000]->out sram[1000]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1000]->out) 0
.nodeset V(sram[1000]->outb) vsp
Xsram[1001] sram->in sram[1001]->out sram[1001]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1001]->out) 0
.nodeset V(sram[1001]->outb) vsp
Xmux_2level_size50[22] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[3]->in[4] sram[1002]->outb sram[1002]->out sram[1003]->out sram[1003]->outb sram[1004]->out sram[1004]->outb sram[1005]->out sram[1005]->outb sram[1006]->out sram[1006]->outb sram[1007]->out sram[1007]->outb sram[1008]->out sram[1008]->outb sram[1009]->out sram[1009]->outb sram[1010]->outb sram[1010]->out sram[1011]->out sram[1011]->outb sram[1012]->out sram[1012]->outb sram[1013]->out sram[1013]->outb sram[1014]->out sram[1014]->outb sram[1015]->out sram[1015]->outb sram[1016]->out sram[1016]->outb sram[1017]->out sram[1017]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[22], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1002] sram->in sram[1002]->out sram[1002]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1002]->out) 0
.nodeset V(sram[1002]->outb) vsp
Xsram[1003] sram->in sram[1003]->out sram[1003]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1003]->out) 0
.nodeset V(sram[1003]->outb) vsp
Xsram[1004] sram->in sram[1004]->out sram[1004]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1004]->out) 0
.nodeset V(sram[1004]->outb) vsp
Xsram[1005] sram->in sram[1005]->out sram[1005]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1005]->out) 0
.nodeset V(sram[1005]->outb) vsp
Xsram[1006] sram->in sram[1006]->out sram[1006]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1006]->out) 0
.nodeset V(sram[1006]->outb) vsp
Xsram[1007] sram->in sram[1007]->out sram[1007]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1007]->out) 0
.nodeset V(sram[1007]->outb) vsp
Xsram[1008] sram->in sram[1008]->out sram[1008]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1008]->out) 0
.nodeset V(sram[1008]->outb) vsp
Xsram[1009] sram->in sram[1009]->out sram[1009]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1009]->out) 0
.nodeset V(sram[1009]->outb) vsp
Xsram[1010] sram->in sram[1010]->out sram[1010]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1010]->out) 0
.nodeset V(sram[1010]->outb) vsp
Xsram[1011] sram->in sram[1011]->out sram[1011]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1011]->out) 0
.nodeset V(sram[1011]->outb) vsp
Xsram[1012] sram->in sram[1012]->out sram[1012]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1012]->out) 0
.nodeset V(sram[1012]->outb) vsp
Xsram[1013] sram->in sram[1013]->out sram[1013]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1013]->out) 0
.nodeset V(sram[1013]->outb) vsp
Xsram[1014] sram->in sram[1014]->out sram[1014]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1014]->out) 0
.nodeset V(sram[1014]->outb) vsp
Xsram[1015] sram->in sram[1015]->out sram[1015]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1015]->out) 0
.nodeset V(sram[1015]->outb) vsp
Xsram[1016] sram->in sram[1016]->out sram[1016]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1016]->out) 0
.nodeset V(sram[1016]->outb) vsp
Xsram[1017] sram->in sram[1017]->out sram[1017]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1017]->out) 0
.nodeset V(sram[1017]->outb) vsp
Xmux_2level_size50[23] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[3]->in[5] sram[1018]->outb sram[1018]->out sram[1019]->out sram[1019]->outb sram[1020]->out sram[1020]->outb sram[1021]->out sram[1021]->outb sram[1022]->out sram[1022]->outb sram[1023]->out sram[1023]->outb sram[1024]->out sram[1024]->outb sram[1025]->out sram[1025]->outb sram[1026]->outb sram[1026]->out sram[1027]->out sram[1027]->outb sram[1028]->out sram[1028]->outb sram[1029]->out sram[1029]->outb sram[1030]->out sram[1030]->outb sram[1031]->out sram[1031]->outb sram[1032]->out sram[1032]->outb sram[1033]->out sram[1033]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[23], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1018] sram->in sram[1018]->out sram[1018]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1018]->out) 0
.nodeset V(sram[1018]->outb) vsp
Xsram[1019] sram->in sram[1019]->out sram[1019]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1019]->out) 0
.nodeset V(sram[1019]->outb) vsp
Xsram[1020] sram->in sram[1020]->out sram[1020]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1020]->out) 0
.nodeset V(sram[1020]->outb) vsp
Xsram[1021] sram->in sram[1021]->out sram[1021]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1021]->out) 0
.nodeset V(sram[1021]->outb) vsp
Xsram[1022] sram->in sram[1022]->out sram[1022]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1022]->out) 0
.nodeset V(sram[1022]->outb) vsp
Xsram[1023] sram->in sram[1023]->out sram[1023]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1023]->out) 0
.nodeset V(sram[1023]->outb) vsp
Xsram[1024] sram->in sram[1024]->out sram[1024]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1024]->out) 0
.nodeset V(sram[1024]->outb) vsp
Xsram[1025] sram->in sram[1025]->out sram[1025]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1025]->out) 0
.nodeset V(sram[1025]->outb) vsp
Xsram[1026] sram->in sram[1026]->out sram[1026]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1026]->out) 0
.nodeset V(sram[1026]->outb) vsp
Xsram[1027] sram->in sram[1027]->out sram[1027]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1027]->out) 0
.nodeset V(sram[1027]->outb) vsp
Xsram[1028] sram->in sram[1028]->out sram[1028]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1028]->out) 0
.nodeset V(sram[1028]->outb) vsp
Xsram[1029] sram->in sram[1029]->out sram[1029]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1029]->out) 0
.nodeset V(sram[1029]->outb) vsp
Xsram[1030] sram->in sram[1030]->out sram[1030]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1030]->out) 0
.nodeset V(sram[1030]->outb) vsp
Xsram[1031] sram->in sram[1031]->out sram[1031]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1031]->out) 0
.nodeset V(sram[1031]->outb) vsp
Xsram[1032] sram->in sram[1032]->out sram[1032]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1032]->out) 0
.nodeset V(sram[1032]->outb) vsp
Xsram[1033] sram->in sram[1033]->out sram[1033]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1033]->out) 0
.nodeset V(sram[1033]->outb) vsp
Xdirect_interc[173] mode[clb]->clk[0] fle[3]->clk[0] gvdd_local_interc sgnd direct_interc
Xmux_2level_size50[24] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[4]->in[0] sram[1034]->outb sram[1034]->out sram[1035]->out sram[1035]->outb sram[1036]->out sram[1036]->outb sram[1037]->out sram[1037]->outb sram[1038]->out sram[1038]->outb sram[1039]->out sram[1039]->outb sram[1040]->out sram[1040]->outb sram[1041]->out sram[1041]->outb sram[1042]->outb sram[1042]->out sram[1043]->out sram[1043]->outb sram[1044]->out sram[1044]->outb sram[1045]->out sram[1045]->outb sram[1046]->out sram[1046]->outb sram[1047]->out sram[1047]->outb sram[1048]->out sram[1048]->outb sram[1049]->out sram[1049]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[24], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1034] sram->in sram[1034]->out sram[1034]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1034]->out) 0
.nodeset V(sram[1034]->outb) vsp
Xsram[1035] sram->in sram[1035]->out sram[1035]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1035]->out) 0
.nodeset V(sram[1035]->outb) vsp
Xsram[1036] sram->in sram[1036]->out sram[1036]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1036]->out) 0
.nodeset V(sram[1036]->outb) vsp
Xsram[1037] sram->in sram[1037]->out sram[1037]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1037]->out) 0
.nodeset V(sram[1037]->outb) vsp
Xsram[1038] sram->in sram[1038]->out sram[1038]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1038]->out) 0
.nodeset V(sram[1038]->outb) vsp
Xsram[1039] sram->in sram[1039]->out sram[1039]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1039]->out) 0
.nodeset V(sram[1039]->outb) vsp
Xsram[1040] sram->in sram[1040]->out sram[1040]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1040]->out) 0
.nodeset V(sram[1040]->outb) vsp
Xsram[1041] sram->in sram[1041]->out sram[1041]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1041]->out) 0
.nodeset V(sram[1041]->outb) vsp
Xsram[1042] sram->in sram[1042]->out sram[1042]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1042]->out) 0
.nodeset V(sram[1042]->outb) vsp
Xsram[1043] sram->in sram[1043]->out sram[1043]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1043]->out) 0
.nodeset V(sram[1043]->outb) vsp
Xsram[1044] sram->in sram[1044]->out sram[1044]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1044]->out) 0
.nodeset V(sram[1044]->outb) vsp
Xsram[1045] sram->in sram[1045]->out sram[1045]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1045]->out) 0
.nodeset V(sram[1045]->outb) vsp
Xsram[1046] sram->in sram[1046]->out sram[1046]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1046]->out) 0
.nodeset V(sram[1046]->outb) vsp
Xsram[1047] sram->in sram[1047]->out sram[1047]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1047]->out) 0
.nodeset V(sram[1047]->outb) vsp
Xsram[1048] sram->in sram[1048]->out sram[1048]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1048]->out) 0
.nodeset V(sram[1048]->outb) vsp
Xsram[1049] sram->in sram[1049]->out sram[1049]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1049]->out) 0
.nodeset V(sram[1049]->outb) vsp
Xmux_2level_size50[25] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[4]->in[1] sram[1050]->outb sram[1050]->out sram[1051]->out sram[1051]->outb sram[1052]->out sram[1052]->outb sram[1053]->out sram[1053]->outb sram[1054]->out sram[1054]->outb sram[1055]->out sram[1055]->outb sram[1056]->out sram[1056]->outb sram[1057]->out sram[1057]->outb sram[1058]->outb sram[1058]->out sram[1059]->out sram[1059]->outb sram[1060]->out sram[1060]->outb sram[1061]->out sram[1061]->outb sram[1062]->out sram[1062]->outb sram[1063]->out sram[1063]->outb sram[1064]->out sram[1064]->outb sram[1065]->out sram[1065]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[25], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1050] sram->in sram[1050]->out sram[1050]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1050]->out) 0
.nodeset V(sram[1050]->outb) vsp
Xsram[1051] sram->in sram[1051]->out sram[1051]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1051]->out) 0
.nodeset V(sram[1051]->outb) vsp
Xsram[1052] sram->in sram[1052]->out sram[1052]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1052]->out) 0
.nodeset V(sram[1052]->outb) vsp
Xsram[1053] sram->in sram[1053]->out sram[1053]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1053]->out) 0
.nodeset V(sram[1053]->outb) vsp
Xsram[1054] sram->in sram[1054]->out sram[1054]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1054]->out) 0
.nodeset V(sram[1054]->outb) vsp
Xsram[1055] sram->in sram[1055]->out sram[1055]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1055]->out) 0
.nodeset V(sram[1055]->outb) vsp
Xsram[1056] sram->in sram[1056]->out sram[1056]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1056]->out) 0
.nodeset V(sram[1056]->outb) vsp
Xsram[1057] sram->in sram[1057]->out sram[1057]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1057]->out) 0
.nodeset V(sram[1057]->outb) vsp
Xsram[1058] sram->in sram[1058]->out sram[1058]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1058]->out) 0
.nodeset V(sram[1058]->outb) vsp
Xsram[1059] sram->in sram[1059]->out sram[1059]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1059]->out) 0
.nodeset V(sram[1059]->outb) vsp
Xsram[1060] sram->in sram[1060]->out sram[1060]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1060]->out) 0
.nodeset V(sram[1060]->outb) vsp
Xsram[1061] sram->in sram[1061]->out sram[1061]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1061]->out) 0
.nodeset V(sram[1061]->outb) vsp
Xsram[1062] sram->in sram[1062]->out sram[1062]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1062]->out) 0
.nodeset V(sram[1062]->outb) vsp
Xsram[1063] sram->in sram[1063]->out sram[1063]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1063]->out) 0
.nodeset V(sram[1063]->outb) vsp
Xsram[1064] sram->in sram[1064]->out sram[1064]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1064]->out) 0
.nodeset V(sram[1064]->outb) vsp
Xsram[1065] sram->in sram[1065]->out sram[1065]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1065]->out) 0
.nodeset V(sram[1065]->outb) vsp
Xmux_2level_size50[26] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[4]->in[2] sram[1066]->outb sram[1066]->out sram[1067]->out sram[1067]->outb sram[1068]->out sram[1068]->outb sram[1069]->out sram[1069]->outb sram[1070]->out sram[1070]->outb sram[1071]->out sram[1071]->outb sram[1072]->out sram[1072]->outb sram[1073]->out sram[1073]->outb sram[1074]->outb sram[1074]->out sram[1075]->out sram[1075]->outb sram[1076]->out sram[1076]->outb sram[1077]->out sram[1077]->outb sram[1078]->out sram[1078]->outb sram[1079]->out sram[1079]->outb sram[1080]->out sram[1080]->outb sram[1081]->out sram[1081]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[26], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1066] sram->in sram[1066]->out sram[1066]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1066]->out) 0
.nodeset V(sram[1066]->outb) vsp
Xsram[1067] sram->in sram[1067]->out sram[1067]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1067]->out) 0
.nodeset V(sram[1067]->outb) vsp
Xsram[1068] sram->in sram[1068]->out sram[1068]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1068]->out) 0
.nodeset V(sram[1068]->outb) vsp
Xsram[1069] sram->in sram[1069]->out sram[1069]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1069]->out) 0
.nodeset V(sram[1069]->outb) vsp
Xsram[1070] sram->in sram[1070]->out sram[1070]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1070]->out) 0
.nodeset V(sram[1070]->outb) vsp
Xsram[1071] sram->in sram[1071]->out sram[1071]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1071]->out) 0
.nodeset V(sram[1071]->outb) vsp
Xsram[1072] sram->in sram[1072]->out sram[1072]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1072]->out) 0
.nodeset V(sram[1072]->outb) vsp
Xsram[1073] sram->in sram[1073]->out sram[1073]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1073]->out) 0
.nodeset V(sram[1073]->outb) vsp
Xsram[1074] sram->in sram[1074]->out sram[1074]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1074]->out) 0
.nodeset V(sram[1074]->outb) vsp
Xsram[1075] sram->in sram[1075]->out sram[1075]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1075]->out) 0
.nodeset V(sram[1075]->outb) vsp
Xsram[1076] sram->in sram[1076]->out sram[1076]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1076]->out) 0
.nodeset V(sram[1076]->outb) vsp
Xsram[1077] sram->in sram[1077]->out sram[1077]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1077]->out) 0
.nodeset V(sram[1077]->outb) vsp
Xsram[1078] sram->in sram[1078]->out sram[1078]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1078]->out) 0
.nodeset V(sram[1078]->outb) vsp
Xsram[1079] sram->in sram[1079]->out sram[1079]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1079]->out) 0
.nodeset V(sram[1079]->outb) vsp
Xsram[1080] sram->in sram[1080]->out sram[1080]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1080]->out) 0
.nodeset V(sram[1080]->outb) vsp
Xsram[1081] sram->in sram[1081]->out sram[1081]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1081]->out) 0
.nodeset V(sram[1081]->outb) vsp
Xmux_2level_size50[27] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[4]->in[3] sram[1082]->outb sram[1082]->out sram[1083]->out sram[1083]->outb sram[1084]->out sram[1084]->outb sram[1085]->out sram[1085]->outb sram[1086]->out sram[1086]->outb sram[1087]->out sram[1087]->outb sram[1088]->out sram[1088]->outb sram[1089]->out sram[1089]->outb sram[1090]->outb sram[1090]->out sram[1091]->out sram[1091]->outb sram[1092]->out sram[1092]->outb sram[1093]->out sram[1093]->outb sram[1094]->out sram[1094]->outb sram[1095]->out sram[1095]->outb sram[1096]->out sram[1096]->outb sram[1097]->out sram[1097]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[27], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1082] sram->in sram[1082]->out sram[1082]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1082]->out) 0
.nodeset V(sram[1082]->outb) vsp
Xsram[1083] sram->in sram[1083]->out sram[1083]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1083]->out) 0
.nodeset V(sram[1083]->outb) vsp
Xsram[1084] sram->in sram[1084]->out sram[1084]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1084]->out) 0
.nodeset V(sram[1084]->outb) vsp
Xsram[1085] sram->in sram[1085]->out sram[1085]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1085]->out) 0
.nodeset V(sram[1085]->outb) vsp
Xsram[1086] sram->in sram[1086]->out sram[1086]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1086]->out) 0
.nodeset V(sram[1086]->outb) vsp
Xsram[1087] sram->in sram[1087]->out sram[1087]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1087]->out) 0
.nodeset V(sram[1087]->outb) vsp
Xsram[1088] sram->in sram[1088]->out sram[1088]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1088]->out) 0
.nodeset V(sram[1088]->outb) vsp
Xsram[1089] sram->in sram[1089]->out sram[1089]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1089]->out) 0
.nodeset V(sram[1089]->outb) vsp
Xsram[1090] sram->in sram[1090]->out sram[1090]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1090]->out) 0
.nodeset V(sram[1090]->outb) vsp
Xsram[1091] sram->in sram[1091]->out sram[1091]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1091]->out) 0
.nodeset V(sram[1091]->outb) vsp
Xsram[1092] sram->in sram[1092]->out sram[1092]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1092]->out) 0
.nodeset V(sram[1092]->outb) vsp
Xsram[1093] sram->in sram[1093]->out sram[1093]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1093]->out) 0
.nodeset V(sram[1093]->outb) vsp
Xsram[1094] sram->in sram[1094]->out sram[1094]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1094]->out) 0
.nodeset V(sram[1094]->outb) vsp
Xsram[1095] sram->in sram[1095]->out sram[1095]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1095]->out) 0
.nodeset V(sram[1095]->outb) vsp
Xsram[1096] sram->in sram[1096]->out sram[1096]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1096]->out) 0
.nodeset V(sram[1096]->outb) vsp
Xsram[1097] sram->in sram[1097]->out sram[1097]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1097]->out) 0
.nodeset V(sram[1097]->outb) vsp
Xmux_2level_size50[28] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[4]->in[4] sram[1098]->outb sram[1098]->out sram[1099]->out sram[1099]->outb sram[1100]->out sram[1100]->outb sram[1101]->out sram[1101]->outb sram[1102]->out sram[1102]->outb sram[1103]->out sram[1103]->outb sram[1104]->out sram[1104]->outb sram[1105]->out sram[1105]->outb sram[1106]->outb sram[1106]->out sram[1107]->out sram[1107]->outb sram[1108]->out sram[1108]->outb sram[1109]->out sram[1109]->outb sram[1110]->out sram[1110]->outb sram[1111]->out sram[1111]->outb sram[1112]->out sram[1112]->outb sram[1113]->out sram[1113]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[28], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1098] sram->in sram[1098]->out sram[1098]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1098]->out) 0
.nodeset V(sram[1098]->outb) vsp
Xsram[1099] sram->in sram[1099]->out sram[1099]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1099]->out) 0
.nodeset V(sram[1099]->outb) vsp
Xsram[1100] sram->in sram[1100]->out sram[1100]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1100]->out) 0
.nodeset V(sram[1100]->outb) vsp
Xsram[1101] sram->in sram[1101]->out sram[1101]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1101]->out) 0
.nodeset V(sram[1101]->outb) vsp
Xsram[1102] sram->in sram[1102]->out sram[1102]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1102]->out) 0
.nodeset V(sram[1102]->outb) vsp
Xsram[1103] sram->in sram[1103]->out sram[1103]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1103]->out) 0
.nodeset V(sram[1103]->outb) vsp
Xsram[1104] sram->in sram[1104]->out sram[1104]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1104]->out) 0
.nodeset V(sram[1104]->outb) vsp
Xsram[1105] sram->in sram[1105]->out sram[1105]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1105]->out) 0
.nodeset V(sram[1105]->outb) vsp
Xsram[1106] sram->in sram[1106]->out sram[1106]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1106]->out) 0
.nodeset V(sram[1106]->outb) vsp
Xsram[1107] sram->in sram[1107]->out sram[1107]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1107]->out) 0
.nodeset V(sram[1107]->outb) vsp
Xsram[1108] sram->in sram[1108]->out sram[1108]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1108]->out) 0
.nodeset V(sram[1108]->outb) vsp
Xsram[1109] sram->in sram[1109]->out sram[1109]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1109]->out) 0
.nodeset V(sram[1109]->outb) vsp
Xsram[1110] sram->in sram[1110]->out sram[1110]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1110]->out) 0
.nodeset V(sram[1110]->outb) vsp
Xsram[1111] sram->in sram[1111]->out sram[1111]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1111]->out) 0
.nodeset V(sram[1111]->outb) vsp
Xsram[1112] sram->in sram[1112]->out sram[1112]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1112]->out) 0
.nodeset V(sram[1112]->outb) vsp
Xsram[1113] sram->in sram[1113]->out sram[1113]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1113]->out) 0
.nodeset V(sram[1113]->outb) vsp
Xmux_2level_size50[29] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[4]->in[5] sram[1114]->outb sram[1114]->out sram[1115]->out sram[1115]->outb sram[1116]->out sram[1116]->outb sram[1117]->out sram[1117]->outb sram[1118]->out sram[1118]->outb sram[1119]->out sram[1119]->outb sram[1120]->out sram[1120]->outb sram[1121]->out sram[1121]->outb sram[1122]->outb sram[1122]->out sram[1123]->out sram[1123]->outb sram[1124]->out sram[1124]->outb sram[1125]->out sram[1125]->outb sram[1126]->out sram[1126]->outb sram[1127]->out sram[1127]->outb sram[1128]->out sram[1128]->outb sram[1129]->out sram[1129]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[29], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1114] sram->in sram[1114]->out sram[1114]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1114]->out) 0
.nodeset V(sram[1114]->outb) vsp
Xsram[1115] sram->in sram[1115]->out sram[1115]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1115]->out) 0
.nodeset V(sram[1115]->outb) vsp
Xsram[1116] sram->in sram[1116]->out sram[1116]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1116]->out) 0
.nodeset V(sram[1116]->outb) vsp
Xsram[1117] sram->in sram[1117]->out sram[1117]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1117]->out) 0
.nodeset V(sram[1117]->outb) vsp
Xsram[1118] sram->in sram[1118]->out sram[1118]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1118]->out) 0
.nodeset V(sram[1118]->outb) vsp
Xsram[1119] sram->in sram[1119]->out sram[1119]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1119]->out) 0
.nodeset V(sram[1119]->outb) vsp
Xsram[1120] sram->in sram[1120]->out sram[1120]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1120]->out) 0
.nodeset V(sram[1120]->outb) vsp
Xsram[1121] sram->in sram[1121]->out sram[1121]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1121]->out) 0
.nodeset V(sram[1121]->outb) vsp
Xsram[1122] sram->in sram[1122]->out sram[1122]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1122]->out) 0
.nodeset V(sram[1122]->outb) vsp
Xsram[1123] sram->in sram[1123]->out sram[1123]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1123]->out) 0
.nodeset V(sram[1123]->outb) vsp
Xsram[1124] sram->in sram[1124]->out sram[1124]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1124]->out) 0
.nodeset V(sram[1124]->outb) vsp
Xsram[1125] sram->in sram[1125]->out sram[1125]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1125]->out) 0
.nodeset V(sram[1125]->outb) vsp
Xsram[1126] sram->in sram[1126]->out sram[1126]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1126]->out) 0
.nodeset V(sram[1126]->outb) vsp
Xsram[1127] sram->in sram[1127]->out sram[1127]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1127]->out) 0
.nodeset V(sram[1127]->outb) vsp
Xsram[1128] sram->in sram[1128]->out sram[1128]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1128]->out) 0
.nodeset V(sram[1128]->outb) vsp
Xsram[1129] sram->in sram[1129]->out sram[1129]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1129]->out) 0
.nodeset V(sram[1129]->outb) vsp
Xdirect_interc[174] mode[clb]->clk[0] fle[4]->clk[0] gvdd_local_interc sgnd direct_interc
Xmux_2level_size50[30] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[5]->in[0] sram[1130]->outb sram[1130]->out sram[1131]->out sram[1131]->outb sram[1132]->out sram[1132]->outb sram[1133]->out sram[1133]->outb sram[1134]->out sram[1134]->outb sram[1135]->out sram[1135]->outb sram[1136]->out sram[1136]->outb sram[1137]->out sram[1137]->outb sram[1138]->outb sram[1138]->out sram[1139]->out sram[1139]->outb sram[1140]->out sram[1140]->outb sram[1141]->out sram[1141]->outb sram[1142]->out sram[1142]->outb sram[1143]->out sram[1143]->outb sram[1144]->out sram[1144]->outb sram[1145]->out sram[1145]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[30], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1130] sram->in sram[1130]->out sram[1130]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1130]->out) 0
.nodeset V(sram[1130]->outb) vsp
Xsram[1131] sram->in sram[1131]->out sram[1131]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1131]->out) 0
.nodeset V(sram[1131]->outb) vsp
Xsram[1132] sram->in sram[1132]->out sram[1132]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1132]->out) 0
.nodeset V(sram[1132]->outb) vsp
Xsram[1133] sram->in sram[1133]->out sram[1133]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1133]->out) 0
.nodeset V(sram[1133]->outb) vsp
Xsram[1134] sram->in sram[1134]->out sram[1134]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1134]->out) 0
.nodeset V(sram[1134]->outb) vsp
Xsram[1135] sram->in sram[1135]->out sram[1135]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1135]->out) 0
.nodeset V(sram[1135]->outb) vsp
Xsram[1136] sram->in sram[1136]->out sram[1136]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1136]->out) 0
.nodeset V(sram[1136]->outb) vsp
Xsram[1137] sram->in sram[1137]->out sram[1137]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1137]->out) 0
.nodeset V(sram[1137]->outb) vsp
Xsram[1138] sram->in sram[1138]->out sram[1138]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1138]->out) 0
.nodeset V(sram[1138]->outb) vsp
Xsram[1139] sram->in sram[1139]->out sram[1139]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1139]->out) 0
.nodeset V(sram[1139]->outb) vsp
Xsram[1140] sram->in sram[1140]->out sram[1140]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1140]->out) 0
.nodeset V(sram[1140]->outb) vsp
Xsram[1141] sram->in sram[1141]->out sram[1141]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1141]->out) 0
.nodeset V(sram[1141]->outb) vsp
Xsram[1142] sram->in sram[1142]->out sram[1142]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1142]->out) 0
.nodeset V(sram[1142]->outb) vsp
Xsram[1143] sram->in sram[1143]->out sram[1143]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1143]->out) 0
.nodeset V(sram[1143]->outb) vsp
Xsram[1144] sram->in sram[1144]->out sram[1144]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1144]->out) 0
.nodeset V(sram[1144]->outb) vsp
Xsram[1145] sram->in sram[1145]->out sram[1145]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1145]->out) 0
.nodeset V(sram[1145]->outb) vsp
Xmux_2level_size50[31] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[5]->in[1] sram[1146]->outb sram[1146]->out sram[1147]->out sram[1147]->outb sram[1148]->out sram[1148]->outb sram[1149]->out sram[1149]->outb sram[1150]->out sram[1150]->outb sram[1151]->out sram[1151]->outb sram[1152]->out sram[1152]->outb sram[1153]->out sram[1153]->outb sram[1154]->outb sram[1154]->out sram[1155]->out sram[1155]->outb sram[1156]->out sram[1156]->outb sram[1157]->out sram[1157]->outb sram[1158]->out sram[1158]->outb sram[1159]->out sram[1159]->outb sram[1160]->out sram[1160]->outb sram[1161]->out sram[1161]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[31], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1146] sram->in sram[1146]->out sram[1146]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1146]->out) 0
.nodeset V(sram[1146]->outb) vsp
Xsram[1147] sram->in sram[1147]->out sram[1147]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1147]->out) 0
.nodeset V(sram[1147]->outb) vsp
Xsram[1148] sram->in sram[1148]->out sram[1148]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1148]->out) 0
.nodeset V(sram[1148]->outb) vsp
Xsram[1149] sram->in sram[1149]->out sram[1149]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1149]->out) 0
.nodeset V(sram[1149]->outb) vsp
Xsram[1150] sram->in sram[1150]->out sram[1150]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1150]->out) 0
.nodeset V(sram[1150]->outb) vsp
Xsram[1151] sram->in sram[1151]->out sram[1151]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1151]->out) 0
.nodeset V(sram[1151]->outb) vsp
Xsram[1152] sram->in sram[1152]->out sram[1152]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1152]->out) 0
.nodeset V(sram[1152]->outb) vsp
Xsram[1153] sram->in sram[1153]->out sram[1153]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1153]->out) 0
.nodeset V(sram[1153]->outb) vsp
Xsram[1154] sram->in sram[1154]->out sram[1154]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1154]->out) 0
.nodeset V(sram[1154]->outb) vsp
Xsram[1155] sram->in sram[1155]->out sram[1155]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1155]->out) 0
.nodeset V(sram[1155]->outb) vsp
Xsram[1156] sram->in sram[1156]->out sram[1156]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1156]->out) 0
.nodeset V(sram[1156]->outb) vsp
Xsram[1157] sram->in sram[1157]->out sram[1157]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1157]->out) 0
.nodeset V(sram[1157]->outb) vsp
Xsram[1158] sram->in sram[1158]->out sram[1158]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1158]->out) 0
.nodeset V(sram[1158]->outb) vsp
Xsram[1159] sram->in sram[1159]->out sram[1159]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1159]->out) 0
.nodeset V(sram[1159]->outb) vsp
Xsram[1160] sram->in sram[1160]->out sram[1160]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1160]->out) 0
.nodeset V(sram[1160]->outb) vsp
Xsram[1161] sram->in sram[1161]->out sram[1161]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1161]->out) 0
.nodeset V(sram[1161]->outb) vsp
Xmux_2level_size50[32] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[5]->in[2] sram[1162]->outb sram[1162]->out sram[1163]->out sram[1163]->outb sram[1164]->out sram[1164]->outb sram[1165]->out sram[1165]->outb sram[1166]->out sram[1166]->outb sram[1167]->out sram[1167]->outb sram[1168]->out sram[1168]->outb sram[1169]->out sram[1169]->outb sram[1170]->outb sram[1170]->out sram[1171]->out sram[1171]->outb sram[1172]->out sram[1172]->outb sram[1173]->out sram[1173]->outb sram[1174]->out sram[1174]->outb sram[1175]->out sram[1175]->outb sram[1176]->out sram[1176]->outb sram[1177]->out sram[1177]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[32], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1162] sram->in sram[1162]->out sram[1162]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1162]->out) 0
.nodeset V(sram[1162]->outb) vsp
Xsram[1163] sram->in sram[1163]->out sram[1163]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1163]->out) 0
.nodeset V(sram[1163]->outb) vsp
Xsram[1164] sram->in sram[1164]->out sram[1164]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1164]->out) 0
.nodeset V(sram[1164]->outb) vsp
Xsram[1165] sram->in sram[1165]->out sram[1165]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1165]->out) 0
.nodeset V(sram[1165]->outb) vsp
Xsram[1166] sram->in sram[1166]->out sram[1166]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1166]->out) 0
.nodeset V(sram[1166]->outb) vsp
Xsram[1167] sram->in sram[1167]->out sram[1167]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1167]->out) 0
.nodeset V(sram[1167]->outb) vsp
Xsram[1168] sram->in sram[1168]->out sram[1168]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1168]->out) 0
.nodeset V(sram[1168]->outb) vsp
Xsram[1169] sram->in sram[1169]->out sram[1169]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1169]->out) 0
.nodeset V(sram[1169]->outb) vsp
Xsram[1170] sram->in sram[1170]->out sram[1170]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1170]->out) 0
.nodeset V(sram[1170]->outb) vsp
Xsram[1171] sram->in sram[1171]->out sram[1171]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1171]->out) 0
.nodeset V(sram[1171]->outb) vsp
Xsram[1172] sram->in sram[1172]->out sram[1172]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1172]->out) 0
.nodeset V(sram[1172]->outb) vsp
Xsram[1173] sram->in sram[1173]->out sram[1173]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1173]->out) 0
.nodeset V(sram[1173]->outb) vsp
Xsram[1174] sram->in sram[1174]->out sram[1174]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1174]->out) 0
.nodeset V(sram[1174]->outb) vsp
Xsram[1175] sram->in sram[1175]->out sram[1175]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1175]->out) 0
.nodeset V(sram[1175]->outb) vsp
Xsram[1176] sram->in sram[1176]->out sram[1176]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1176]->out) 0
.nodeset V(sram[1176]->outb) vsp
Xsram[1177] sram->in sram[1177]->out sram[1177]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1177]->out) 0
.nodeset V(sram[1177]->outb) vsp
Xmux_2level_size50[33] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[5]->in[3] sram[1178]->outb sram[1178]->out sram[1179]->out sram[1179]->outb sram[1180]->out sram[1180]->outb sram[1181]->out sram[1181]->outb sram[1182]->out sram[1182]->outb sram[1183]->out sram[1183]->outb sram[1184]->out sram[1184]->outb sram[1185]->out sram[1185]->outb sram[1186]->outb sram[1186]->out sram[1187]->out sram[1187]->outb sram[1188]->out sram[1188]->outb sram[1189]->out sram[1189]->outb sram[1190]->out sram[1190]->outb sram[1191]->out sram[1191]->outb sram[1192]->out sram[1192]->outb sram[1193]->out sram[1193]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[33], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1178] sram->in sram[1178]->out sram[1178]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1178]->out) 0
.nodeset V(sram[1178]->outb) vsp
Xsram[1179] sram->in sram[1179]->out sram[1179]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1179]->out) 0
.nodeset V(sram[1179]->outb) vsp
Xsram[1180] sram->in sram[1180]->out sram[1180]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1180]->out) 0
.nodeset V(sram[1180]->outb) vsp
Xsram[1181] sram->in sram[1181]->out sram[1181]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1181]->out) 0
.nodeset V(sram[1181]->outb) vsp
Xsram[1182] sram->in sram[1182]->out sram[1182]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1182]->out) 0
.nodeset V(sram[1182]->outb) vsp
Xsram[1183] sram->in sram[1183]->out sram[1183]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1183]->out) 0
.nodeset V(sram[1183]->outb) vsp
Xsram[1184] sram->in sram[1184]->out sram[1184]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1184]->out) 0
.nodeset V(sram[1184]->outb) vsp
Xsram[1185] sram->in sram[1185]->out sram[1185]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1185]->out) 0
.nodeset V(sram[1185]->outb) vsp
Xsram[1186] sram->in sram[1186]->out sram[1186]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1186]->out) 0
.nodeset V(sram[1186]->outb) vsp
Xsram[1187] sram->in sram[1187]->out sram[1187]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1187]->out) 0
.nodeset V(sram[1187]->outb) vsp
Xsram[1188] sram->in sram[1188]->out sram[1188]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1188]->out) 0
.nodeset V(sram[1188]->outb) vsp
Xsram[1189] sram->in sram[1189]->out sram[1189]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1189]->out) 0
.nodeset V(sram[1189]->outb) vsp
Xsram[1190] sram->in sram[1190]->out sram[1190]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1190]->out) 0
.nodeset V(sram[1190]->outb) vsp
Xsram[1191] sram->in sram[1191]->out sram[1191]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1191]->out) 0
.nodeset V(sram[1191]->outb) vsp
Xsram[1192] sram->in sram[1192]->out sram[1192]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1192]->out) 0
.nodeset V(sram[1192]->outb) vsp
Xsram[1193] sram->in sram[1193]->out sram[1193]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1193]->out) 0
.nodeset V(sram[1193]->outb) vsp
Xmux_2level_size50[34] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[5]->in[4] sram[1194]->outb sram[1194]->out sram[1195]->out sram[1195]->outb sram[1196]->out sram[1196]->outb sram[1197]->out sram[1197]->outb sram[1198]->out sram[1198]->outb sram[1199]->out sram[1199]->outb sram[1200]->out sram[1200]->outb sram[1201]->out sram[1201]->outb sram[1202]->outb sram[1202]->out sram[1203]->out sram[1203]->outb sram[1204]->out sram[1204]->outb sram[1205]->out sram[1205]->outb sram[1206]->out sram[1206]->outb sram[1207]->out sram[1207]->outb sram[1208]->out sram[1208]->outb sram[1209]->out sram[1209]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[34], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1194] sram->in sram[1194]->out sram[1194]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1194]->out) 0
.nodeset V(sram[1194]->outb) vsp
Xsram[1195] sram->in sram[1195]->out sram[1195]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1195]->out) 0
.nodeset V(sram[1195]->outb) vsp
Xsram[1196] sram->in sram[1196]->out sram[1196]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1196]->out) 0
.nodeset V(sram[1196]->outb) vsp
Xsram[1197] sram->in sram[1197]->out sram[1197]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1197]->out) 0
.nodeset V(sram[1197]->outb) vsp
Xsram[1198] sram->in sram[1198]->out sram[1198]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1198]->out) 0
.nodeset V(sram[1198]->outb) vsp
Xsram[1199] sram->in sram[1199]->out sram[1199]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1199]->out) 0
.nodeset V(sram[1199]->outb) vsp
Xsram[1200] sram->in sram[1200]->out sram[1200]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1200]->out) 0
.nodeset V(sram[1200]->outb) vsp
Xsram[1201] sram->in sram[1201]->out sram[1201]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1201]->out) 0
.nodeset V(sram[1201]->outb) vsp
Xsram[1202] sram->in sram[1202]->out sram[1202]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1202]->out) 0
.nodeset V(sram[1202]->outb) vsp
Xsram[1203] sram->in sram[1203]->out sram[1203]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1203]->out) 0
.nodeset V(sram[1203]->outb) vsp
Xsram[1204] sram->in sram[1204]->out sram[1204]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1204]->out) 0
.nodeset V(sram[1204]->outb) vsp
Xsram[1205] sram->in sram[1205]->out sram[1205]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1205]->out) 0
.nodeset V(sram[1205]->outb) vsp
Xsram[1206] sram->in sram[1206]->out sram[1206]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1206]->out) 0
.nodeset V(sram[1206]->outb) vsp
Xsram[1207] sram->in sram[1207]->out sram[1207]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1207]->out) 0
.nodeset V(sram[1207]->outb) vsp
Xsram[1208] sram->in sram[1208]->out sram[1208]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1208]->out) 0
.nodeset V(sram[1208]->outb) vsp
Xsram[1209] sram->in sram[1209]->out sram[1209]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1209]->out) 0
.nodeset V(sram[1209]->outb) vsp
Xmux_2level_size50[35] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[5]->in[5] sram[1210]->outb sram[1210]->out sram[1211]->out sram[1211]->outb sram[1212]->out sram[1212]->outb sram[1213]->out sram[1213]->outb sram[1214]->out sram[1214]->outb sram[1215]->out sram[1215]->outb sram[1216]->out sram[1216]->outb sram[1217]->out sram[1217]->outb sram[1218]->outb sram[1218]->out sram[1219]->out sram[1219]->outb sram[1220]->out sram[1220]->outb sram[1221]->out sram[1221]->outb sram[1222]->out sram[1222]->outb sram[1223]->out sram[1223]->outb sram[1224]->out sram[1224]->outb sram[1225]->out sram[1225]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[35], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1210] sram->in sram[1210]->out sram[1210]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1210]->out) 0
.nodeset V(sram[1210]->outb) vsp
Xsram[1211] sram->in sram[1211]->out sram[1211]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1211]->out) 0
.nodeset V(sram[1211]->outb) vsp
Xsram[1212] sram->in sram[1212]->out sram[1212]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1212]->out) 0
.nodeset V(sram[1212]->outb) vsp
Xsram[1213] sram->in sram[1213]->out sram[1213]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1213]->out) 0
.nodeset V(sram[1213]->outb) vsp
Xsram[1214] sram->in sram[1214]->out sram[1214]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1214]->out) 0
.nodeset V(sram[1214]->outb) vsp
Xsram[1215] sram->in sram[1215]->out sram[1215]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1215]->out) 0
.nodeset V(sram[1215]->outb) vsp
Xsram[1216] sram->in sram[1216]->out sram[1216]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1216]->out) 0
.nodeset V(sram[1216]->outb) vsp
Xsram[1217] sram->in sram[1217]->out sram[1217]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1217]->out) 0
.nodeset V(sram[1217]->outb) vsp
Xsram[1218] sram->in sram[1218]->out sram[1218]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1218]->out) 0
.nodeset V(sram[1218]->outb) vsp
Xsram[1219] sram->in sram[1219]->out sram[1219]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1219]->out) 0
.nodeset V(sram[1219]->outb) vsp
Xsram[1220] sram->in sram[1220]->out sram[1220]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1220]->out) 0
.nodeset V(sram[1220]->outb) vsp
Xsram[1221] sram->in sram[1221]->out sram[1221]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1221]->out) 0
.nodeset V(sram[1221]->outb) vsp
Xsram[1222] sram->in sram[1222]->out sram[1222]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1222]->out) 0
.nodeset V(sram[1222]->outb) vsp
Xsram[1223] sram->in sram[1223]->out sram[1223]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1223]->out) 0
.nodeset V(sram[1223]->outb) vsp
Xsram[1224] sram->in sram[1224]->out sram[1224]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1224]->out) 0
.nodeset V(sram[1224]->outb) vsp
Xsram[1225] sram->in sram[1225]->out sram[1225]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1225]->out) 0
.nodeset V(sram[1225]->outb) vsp
Xdirect_interc[175] mode[clb]->clk[0] fle[5]->clk[0] gvdd_local_interc sgnd direct_interc
Xmux_2level_size50[36] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[6]->in[0] sram[1226]->outb sram[1226]->out sram[1227]->out sram[1227]->outb sram[1228]->out sram[1228]->outb sram[1229]->out sram[1229]->outb sram[1230]->out sram[1230]->outb sram[1231]->out sram[1231]->outb sram[1232]->out sram[1232]->outb sram[1233]->out sram[1233]->outb sram[1234]->outb sram[1234]->out sram[1235]->out sram[1235]->outb sram[1236]->out sram[1236]->outb sram[1237]->out sram[1237]->outb sram[1238]->out sram[1238]->outb sram[1239]->out sram[1239]->outb sram[1240]->out sram[1240]->outb sram[1241]->out sram[1241]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[36], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1226] sram->in sram[1226]->out sram[1226]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1226]->out) 0
.nodeset V(sram[1226]->outb) vsp
Xsram[1227] sram->in sram[1227]->out sram[1227]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1227]->out) 0
.nodeset V(sram[1227]->outb) vsp
Xsram[1228] sram->in sram[1228]->out sram[1228]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1228]->out) 0
.nodeset V(sram[1228]->outb) vsp
Xsram[1229] sram->in sram[1229]->out sram[1229]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1229]->out) 0
.nodeset V(sram[1229]->outb) vsp
Xsram[1230] sram->in sram[1230]->out sram[1230]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1230]->out) 0
.nodeset V(sram[1230]->outb) vsp
Xsram[1231] sram->in sram[1231]->out sram[1231]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1231]->out) 0
.nodeset V(sram[1231]->outb) vsp
Xsram[1232] sram->in sram[1232]->out sram[1232]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1232]->out) 0
.nodeset V(sram[1232]->outb) vsp
Xsram[1233] sram->in sram[1233]->out sram[1233]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1233]->out) 0
.nodeset V(sram[1233]->outb) vsp
Xsram[1234] sram->in sram[1234]->out sram[1234]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1234]->out) 0
.nodeset V(sram[1234]->outb) vsp
Xsram[1235] sram->in sram[1235]->out sram[1235]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1235]->out) 0
.nodeset V(sram[1235]->outb) vsp
Xsram[1236] sram->in sram[1236]->out sram[1236]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1236]->out) 0
.nodeset V(sram[1236]->outb) vsp
Xsram[1237] sram->in sram[1237]->out sram[1237]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1237]->out) 0
.nodeset V(sram[1237]->outb) vsp
Xsram[1238] sram->in sram[1238]->out sram[1238]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1238]->out) 0
.nodeset V(sram[1238]->outb) vsp
Xsram[1239] sram->in sram[1239]->out sram[1239]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1239]->out) 0
.nodeset V(sram[1239]->outb) vsp
Xsram[1240] sram->in sram[1240]->out sram[1240]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1240]->out) 0
.nodeset V(sram[1240]->outb) vsp
Xsram[1241] sram->in sram[1241]->out sram[1241]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1241]->out) 0
.nodeset V(sram[1241]->outb) vsp
Xmux_2level_size50[37] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[6]->in[1] sram[1242]->outb sram[1242]->out sram[1243]->out sram[1243]->outb sram[1244]->out sram[1244]->outb sram[1245]->out sram[1245]->outb sram[1246]->out sram[1246]->outb sram[1247]->out sram[1247]->outb sram[1248]->out sram[1248]->outb sram[1249]->out sram[1249]->outb sram[1250]->outb sram[1250]->out sram[1251]->out sram[1251]->outb sram[1252]->out sram[1252]->outb sram[1253]->out sram[1253]->outb sram[1254]->out sram[1254]->outb sram[1255]->out sram[1255]->outb sram[1256]->out sram[1256]->outb sram[1257]->out sram[1257]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[37], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1242] sram->in sram[1242]->out sram[1242]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1242]->out) 0
.nodeset V(sram[1242]->outb) vsp
Xsram[1243] sram->in sram[1243]->out sram[1243]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1243]->out) 0
.nodeset V(sram[1243]->outb) vsp
Xsram[1244] sram->in sram[1244]->out sram[1244]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1244]->out) 0
.nodeset V(sram[1244]->outb) vsp
Xsram[1245] sram->in sram[1245]->out sram[1245]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1245]->out) 0
.nodeset V(sram[1245]->outb) vsp
Xsram[1246] sram->in sram[1246]->out sram[1246]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1246]->out) 0
.nodeset V(sram[1246]->outb) vsp
Xsram[1247] sram->in sram[1247]->out sram[1247]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1247]->out) 0
.nodeset V(sram[1247]->outb) vsp
Xsram[1248] sram->in sram[1248]->out sram[1248]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1248]->out) 0
.nodeset V(sram[1248]->outb) vsp
Xsram[1249] sram->in sram[1249]->out sram[1249]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1249]->out) 0
.nodeset V(sram[1249]->outb) vsp
Xsram[1250] sram->in sram[1250]->out sram[1250]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1250]->out) 0
.nodeset V(sram[1250]->outb) vsp
Xsram[1251] sram->in sram[1251]->out sram[1251]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1251]->out) 0
.nodeset V(sram[1251]->outb) vsp
Xsram[1252] sram->in sram[1252]->out sram[1252]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1252]->out) 0
.nodeset V(sram[1252]->outb) vsp
Xsram[1253] sram->in sram[1253]->out sram[1253]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1253]->out) 0
.nodeset V(sram[1253]->outb) vsp
Xsram[1254] sram->in sram[1254]->out sram[1254]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1254]->out) 0
.nodeset V(sram[1254]->outb) vsp
Xsram[1255] sram->in sram[1255]->out sram[1255]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1255]->out) 0
.nodeset V(sram[1255]->outb) vsp
Xsram[1256] sram->in sram[1256]->out sram[1256]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1256]->out) 0
.nodeset V(sram[1256]->outb) vsp
Xsram[1257] sram->in sram[1257]->out sram[1257]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1257]->out) 0
.nodeset V(sram[1257]->outb) vsp
Xmux_2level_size50[38] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[6]->in[2] sram[1258]->outb sram[1258]->out sram[1259]->out sram[1259]->outb sram[1260]->out sram[1260]->outb sram[1261]->out sram[1261]->outb sram[1262]->out sram[1262]->outb sram[1263]->out sram[1263]->outb sram[1264]->out sram[1264]->outb sram[1265]->out sram[1265]->outb sram[1266]->outb sram[1266]->out sram[1267]->out sram[1267]->outb sram[1268]->out sram[1268]->outb sram[1269]->out sram[1269]->outb sram[1270]->out sram[1270]->outb sram[1271]->out sram[1271]->outb sram[1272]->out sram[1272]->outb sram[1273]->out sram[1273]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[38], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1258] sram->in sram[1258]->out sram[1258]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1258]->out) 0
.nodeset V(sram[1258]->outb) vsp
Xsram[1259] sram->in sram[1259]->out sram[1259]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1259]->out) 0
.nodeset V(sram[1259]->outb) vsp
Xsram[1260] sram->in sram[1260]->out sram[1260]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1260]->out) 0
.nodeset V(sram[1260]->outb) vsp
Xsram[1261] sram->in sram[1261]->out sram[1261]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1261]->out) 0
.nodeset V(sram[1261]->outb) vsp
Xsram[1262] sram->in sram[1262]->out sram[1262]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1262]->out) 0
.nodeset V(sram[1262]->outb) vsp
Xsram[1263] sram->in sram[1263]->out sram[1263]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1263]->out) 0
.nodeset V(sram[1263]->outb) vsp
Xsram[1264] sram->in sram[1264]->out sram[1264]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1264]->out) 0
.nodeset V(sram[1264]->outb) vsp
Xsram[1265] sram->in sram[1265]->out sram[1265]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1265]->out) 0
.nodeset V(sram[1265]->outb) vsp
Xsram[1266] sram->in sram[1266]->out sram[1266]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1266]->out) 0
.nodeset V(sram[1266]->outb) vsp
Xsram[1267] sram->in sram[1267]->out sram[1267]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1267]->out) 0
.nodeset V(sram[1267]->outb) vsp
Xsram[1268] sram->in sram[1268]->out sram[1268]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1268]->out) 0
.nodeset V(sram[1268]->outb) vsp
Xsram[1269] sram->in sram[1269]->out sram[1269]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1269]->out) 0
.nodeset V(sram[1269]->outb) vsp
Xsram[1270] sram->in sram[1270]->out sram[1270]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1270]->out) 0
.nodeset V(sram[1270]->outb) vsp
Xsram[1271] sram->in sram[1271]->out sram[1271]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1271]->out) 0
.nodeset V(sram[1271]->outb) vsp
Xsram[1272] sram->in sram[1272]->out sram[1272]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1272]->out) 0
.nodeset V(sram[1272]->outb) vsp
Xsram[1273] sram->in sram[1273]->out sram[1273]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1273]->out) 0
.nodeset V(sram[1273]->outb) vsp
Xmux_2level_size50[39] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[6]->in[3] sram[1274]->outb sram[1274]->out sram[1275]->out sram[1275]->outb sram[1276]->out sram[1276]->outb sram[1277]->out sram[1277]->outb sram[1278]->out sram[1278]->outb sram[1279]->out sram[1279]->outb sram[1280]->out sram[1280]->outb sram[1281]->out sram[1281]->outb sram[1282]->outb sram[1282]->out sram[1283]->out sram[1283]->outb sram[1284]->out sram[1284]->outb sram[1285]->out sram[1285]->outb sram[1286]->out sram[1286]->outb sram[1287]->out sram[1287]->outb sram[1288]->out sram[1288]->outb sram[1289]->out sram[1289]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[39], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1274] sram->in sram[1274]->out sram[1274]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1274]->out) 0
.nodeset V(sram[1274]->outb) vsp
Xsram[1275] sram->in sram[1275]->out sram[1275]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1275]->out) 0
.nodeset V(sram[1275]->outb) vsp
Xsram[1276] sram->in sram[1276]->out sram[1276]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1276]->out) 0
.nodeset V(sram[1276]->outb) vsp
Xsram[1277] sram->in sram[1277]->out sram[1277]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1277]->out) 0
.nodeset V(sram[1277]->outb) vsp
Xsram[1278] sram->in sram[1278]->out sram[1278]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1278]->out) 0
.nodeset V(sram[1278]->outb) vsp
Xsram[1279] sram->in sram[1279]->out sram[1279]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1279]->out) 0
.nodeset V(sram[1279]->outb) vsp
Xsram[1280] sram->in sram[1280]->out sram[1280]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1280]->out) 0
.nodeset V(sram[1280]->outb) vsp
Xsram[1281] sram->in sram[1281]->out sram[1281]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1281]->out) 0
.nodeset V(sram[1281]->outb) vsp
Xsram[1282] sram->in sram[1282]->out sram[1282]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1282]->out) 0
.nodeset V(sram[1282]->outb) vsp
Xsram[1283] sram->in sram[1283]->out sram[1283]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1283]->out) 0
.nodeset V(sram[1283]->outb) vsp
Xsram[1284] sram->in sram[1284]->out sram[1284]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1284]->out) 0
.nodeset V(sram[1284]->outb) vsp
Xsram[1285] sram->in sram[1285]->out sram[1285]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1285]->out) 0
.nodeset V(sram[1285]->outb) vsp
Xsram[1286] sram->in sram[1286]->out sram[1286]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1286]->out) 0
.nodeset V(sram[1286]->outb) vsp
Xsram[1287] sram->in sram[1287]->out sram[1287]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1287]->out) 0
.nodeset V(sram[1287]->outb) vsp
Xsram[1288] sram->in sram[1288]->out sram[1288]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1288]->out) 0
.nodeset V(sram[1288]->outb) vsp
Xsram[1289] sram->in sram[1289]->out sram[1289]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1289]->out) 0
.nodeset V(sram[1289]->outb) vsp
Xmux_2level_size50[40] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[6]->in[4] sram[1290]->outb sram[1290]->out sram[1291]->out sram[1291]->outb sram[1292]->out sram[1292]->outb sram[1293]->out sram[1293]->outb sram[1294]->out sram[1294]->outb sram[1295]->out sram[1295]->outb sram[1296]->out sram[1296]->outb sram[1297]->out sram[1297]->outb sram[1298]->outb sram[1298]->out sram[1299]->out sram[1299]->outb sram[1300]->out sram[1300]->outb sram[1301]->out sram[1301]->outb sram[1302]->out sram[1302]->outb sram[1303]->out sram[1303]->outb sram[1304]->out sram[1304]->outb sram[1305]->out sram[1305]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[40], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1290] sram->in sram[1290]->out sram[1290]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1290]->out) 0
.nodeset V(sram[1290]->outb) vsp
Xsram[1291] sram->in sram[1291]->out sram[1291]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1291]->out) 0
.nodeset V(sram[1291]->outb) vsp
Xsram[1292] sram->in sram[1292]->out sram[1292]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1292]->out) 0
.nodeset V(sram[1292]->outb) vsp
Xsram[1293] sram->in sram[1293]->out sram[1293]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1293]->out) 0
.nodeset V(sram[1293]->outb) vsp
Xsram[1294] sram->in sram[1294]->out sram[1294]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1294]->out) 0
.nodeset V(sram[1294]->outb) vsp
Xsram[1295] sram->in sram[1295]->out sram[1295]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1295]->out) 0
.nodeset V(sram[1295]->outb) vsp
Xsram[1296] sram->in sram[1296]->out sram[1296]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1296]->out) 0
.nodeset V(sram[1296]->outb) vsp
Xsram[1297] sram->in sram[1297]->out sram[1297]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1297]->out) 0
.nodeset V(sram[1297]->outb) vsp
Xsram[1298] sram->in sram[1298]->out sram[1298]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1298]->out) 0
.nodeset V(sram[1298]->outb) vsp
Xsram[1299] sram->in sram[1299]->out sram[1299]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1299]->out) 0
.nodeset V(sram[1299]->outb) vsp
Xsram[1300] sram->in sram[1300]->out sram[1300]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1300]->out) 0
.nodeset V(sram[1300]->outb) vsp
Xsram[1301] sram->in sram[1301]->out sram[1301]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1301]->out) 0
.nodeset V(sram[1301]->outb) vsp
Xsram[1302] sram->in sram[1302]->out sram[1302]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1302]->out) 0
.nodeset V(sram[1302]->outb) vsp
Xsram[1303] sram->in sram[1303]->out sram[1303]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1303]->out) 0
.nodeset V(sram[1303]->outb) vsp
Xsram[1304] sram->in sram[1304]->out sram[1304]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1304]->out) 0
.nodeset V(sram[1304]->outb) vsp
Xsram[1305] sram->in sram[1305]->out sram[1305]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1305]->out) 0
.nodeset V(sram[1305]->outb) vsp
Xmux_2level_size50[41] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[6]->in[5] sram[1306]->outb sram[1306]->out sram[1307]->out sram[1307]->outb sram[1308]->out sram[1308]->outb sram[1309]->out sram[1309]->outb sram[1310]->out sram[1310]->outb sram[1311]->out sram[1311]->outb sram[1312]->out sram[1312]->outb sram[1313]->out sram[1313]->outb sram[1314]->outb sram[1314]->out sram[1315]->out sram[1315]->outb sram[1316]->out sram[1316]->outb sram[1317]->out sram[1317]->outb sram[1318]->out sram[1318]->outb sram[1319]->out sram[1319]->outb sram[1320]->out sram[1320]->outb sram[1321]->out sram[1321]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[41], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1306] sram->in sram[1306]->out sram[1306]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1306]->out) 0
.nodeset V(sram[1306]->outb) vsp
Xsram[1307] sram->in sram[1307]->out sram[1307]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1307]->out) 0
.nodeset V(sram[1307]->outb) vsp
Xsram[1308] sram->in sram[1308]->out sram[1308]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1308]->out) 0
.nodeset V(sram[1308]->outb) vsp
Xsram[1309] sram->in sram[1309]->out sram[1309]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1309]->out) 0
.nodeset V(sram[1309]->outb) vsp
Xsram[1310] sram->in sram[1310]->out sram[1310]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1310]->out) 0
.nodeset V(sram[1310]->outb) vsp
Xsram[1311] sram->in sram[1311]->out sram[1311]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1311]->out) 0
.nodeset V(sram[1311]->outb) vsp
Xsram[1312] sram->in sram[1312]->out sram[1312]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1312]->out) 0
.nodeset V(sram[1312]->outb) vsp
Xsram[1313] sram->in sram[1313]->out sram[1313]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1313]->out) 0
.nodeset V(sram[1313]->outb) vsp
Xsram[1314] sram->in sram[1314]->out sram[1314]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1314]->out) 0
.nodeset V(sram[1314]->outb) vsp
Xsram[1315] sram->in sram[1315]->out sram[1315]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1315]->out) 0
.nodeset V(sram[1315]->outb) vsp
Xsram[1316] sram->in sram[1316]->out sram[1316]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1316]->out) 0
.nodeset V(sram[1316]->outb) vsp
Xsram[1317] sram->in sram[1317]->out sram[1317]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1317]->out) 0
.nodeset V(sram[1317]->outb) vsp
Xsram[1318] sram->in sram[1318]->out sram[1318]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1318]->out) 0
.nodeset V(sram[1318]->outb) vsp
Xsram[1319] sram->in sram[1319]->out sram[1319]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1319]->out) 0
.nodeset V(sram[1319]->outb) vsp
Xsram[1320] sram->in sram[1320]->out sram[1320]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1320]->out) 0
.nodeset V(sram[1320]->outb) vsp
Xsram[1321] sram->in sram[1321]->out sram[1321]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1321]->out) 0
.nodeset V(sram[1321]->outb) vsp
Xdirect_interc[176] mode[clb]->clk[0] fle[6]->clk[0] gvdd_local_interc sgnd direct_interc
Xmux_2level_size50[42] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[7]->in[0] sram[1322]->outb sram[1322]->out sram[1323]->out sram[1323]->outb sram[1324]->out sram[1324]->outb sram[1325]->out sram[1325]->outb sram[1326]->out sram[1326]->outb sram[1327]->out sram[1327]->outb sram[1328]->out sram[1328]->outb sram[1329]->out sram[1329]->outb sram[1330]->outb sram[1330]->out sram[1331]->out sram[1331]->outb sram[1332]->out sram[1332]->outb sram[1333]->out sram[1333]->outb sram[1334]->out sram[1334]->outb sram[1335]->out sram[1335]->outb sram[1336]->out sram[1336]->outb sram[1337]->out sram[1337]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[42], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1322] sram->in sram[1322]->out sram[1322]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1322]->out) 0
.nodeset V(sram[1322]->outb) vsp
Xsram[1323] sram->in sram[1323]->out sram[1323]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1323]->out) 0
.nodeset V(sram[1323]->outb) vsp
Xsram[1324] sram->in sram[1324]->out sram[1324]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1324]->out) 0
.nodeset V(sram[1324]->outb) vsp
Xsram[1325] sram->in sram[1325]->out sram[1325]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1325]->out) 0
.nodeset V(sram[1325]->outb) vsp
Xsram[1326] sram->in sram[1326]->out sram[1326]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1326]->out) 0
.nodeset V(sram[1326]->outb) vsp
Xsram[1327] sram->in sram[1327]->out sram[1327]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1327]->out) 0
.nodeset V(sram[1327]->outb) vsp
Xsram[1328] sram->in sram[1328]->out sram[1328]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1328]->out) 0
.nodeset V(sram[1328]->outb) vsp
Xsram[1329] sram->in sram[1329]->out sram[1329]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1329]->out) 0
.nodeset V(sram[1329]->outb) vsp
Xsram[1330] sram->in sram[1330]->out sram[1330]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1330]->out) 0
.nodeset V(sram[1330]->outb) vsp
Xsram[1331] sram->in sram[1331]->out sram[1331]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1331]->out) 0
.nodeset V(sram[1331]->outb) vsp
Xsram[1332] sram->in sram[1332]->out sram[1332]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1332]->out) 0
.nodeset V(sram[1332]->outb) vsp
Xsram[1333] sram->in sram[1333]->out sram[1333]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1333]->out) 0
.nodeset V(sram[1333]->outb) vsp
Xsram[1334] sram->in sram[1334]->out sram[1334]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1334]->out) 0
.nodeset V(sram[1334]->outb) vsp
Xsram[1335] sram->in sram[1335]->out sram[1335]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1335]->out) 0
.nodeset V(sram[1335]->outb) vsp
Xsram[1336] sram->in sram[1336]->out sram[1336]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1336]->out) 0
.nodeset V(sram[1336]->outb) vsp
Xsram[1337] sram->in sram[1337]->out sram[1337]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1337]->out) 0
.nodeset V(sram[1337]->outb) vsp
Xmux_2level_size50[43] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[7]->in[1] sram[1338]->outb sram[1338]->out sram[1339]->out sram[1339]->outb sram[1340]->out sram[1340]->outb sram[1341]->out sram[1341]->outb sram[1342]->out sram[1342]->outb sram[1343]->out sram[1343]->outb sram[1344]->out sram[1344]->outb sram[1345]->out sram[1345]->outb sram[1346]->outb sram[1346]->out sram[1347]->out sram[1347]->outb sram[1348]->out sram[1348]->outb sram[1349]->out sram[1349]->outb sram[1350]->out sram[1350]->outb sram[1351]->out sram[1351]->outb sram[1352]->out sram[1352]->outb sram[1353]->out sram[1353]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[43], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1338] sram->in sram[1338]->out sram[1338]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1338]->out) 0
.nodeset V(sram[1338]->outb) vsp
Xsram[1339] sram->in sram[1339]->out sram[1339]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1339]->out) 0
.nodeset V(sram[1339]->outb) vsp
Xsram[1340] sram->in sram[1340]->out sram[1340]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1340]->out) 0
.nodeset V(sram[1340]->outb) vsp
Xsram[1341] sram->in sram[1341]->out sram[1341]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1341]->out) 0
.nodeset V(sram[1341]->outb) vsp
Xsram[1342] sram->in sram[1342]->out sram[1342]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1342]->out) 0
.nodeset V(sram[1342]->outb) vsp
Xsram[1343] sram->in sram[1343]->out sram[1343]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1343]->out) 0
.nodeset V(sram[1343]->outb) vsp
Xsram[1344] sram->in sram[1344]->out sram[1344]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1344]->out) 0
.nodeset V(sram[1344]->outb) vsp
Xsram[1345] sram->in sram[1345]->out sram[1345]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1345]->out) 0
.nodeset V(sram[1345]->outb) vsp
Xsram[1346] sram->in sram[1346]->out sram[1346]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1346]->out) 0
.nodeset V(sram[1346]->outb) vsp
Xsram[1347] sram->in sram[1347]->out sram[1347]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1347]->out) 0
.nodeset V(sram[1347]->outb) vsp
Xsram[1348] sram->in sram[1348]->out sram[1348]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1348]->out) 0
.nodeset V(sram[1348]->outb) vsp
Xsram[1349] sram->in sram[1349]->out sram[1349]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1349]->out) 0
.nodeset V(sram[1349]->outb) vsp
Xsram[1350] sram->in sram[1350]->out sram[1350]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1350]->out) 0
.nodeset V(sram[1350]->outb) vsp
Xsram[1351] sram->in sram[1351]->out sram[1351]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1351]->out) 0
.nodeset V(sram[1351]->outb) vsp
Xsram[1352] sram->in sram[1352]->out sram[1352]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1352]->out) 0
.nodeset V(sram[1352]->outb) vsp
Xsram[1353] sram->in sram[1353]->out sram[1353]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1353]->out) 0
.nodeset V(sram[1353]->outb) vsp
Xmux_2level_size50[44] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[7]->in[2] sram[1354]->outb sram[1354]->out sram[1355]->out sram[1355]->outb sram[1356]->out sram[1356]->outb sram[1357]->out sram[1357]->outb sram[1358]->out sram[1358]->outb sram[1359]->out sram[1359]->outb sram[1360]->out sram[1360]->outb sram[1361]->out sram[1361]->outb sram[1362]->outb sram[1362]->out sram[1363]->out sram[1363]->outb sram[1364]->out sram[1364]->outb sram[1365]->out sram[1365]->outb sram[1366]->out sram[1366]->outb sram[1367]->out sram[1367]->outb sram[1368]->out sram[1368]->outb sram[1369]->out sram[1369]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[44], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1354] sram->in sram[1354]->out sram[1354]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1354]->out) 0
.nodeset V(sram[1354]->outb) vsp
Xsram[1355] sram->in sram[1355]->out sram[1355]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1355]->out) 0
.nodeset V(sram[1355]->outb) vsp
Xsram[1356] sram->in sram[1356]->out sram[1356]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1356]->out) 0
.nodeset V(sram[1356]->outb) vsp
Xsram[1357] sram->in sram[1357]->out sram[1357]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1357]->out) 0
.nodeset V(sram[1357]->outb) vsp
Xsram[1358] sram->in sram[1358]->out sram[1358]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1358]->out) 0
.nodeset V(sram[1358]->outb) vsp
Xsram[1359] sram->in sram[1359]->out sram[1359]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1359]->out) 0
.nodeset V(sram[1359]->outb) vsp
Xsram[1360] sram->in sram[1360]->out sram[1360]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1360]->out) 0
.nodeset V(sram[1360]->outb) vsp
Xsram[1361] sram->in sram[1361]->out sram[1361]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1361]->out) 0
.nodeset V(sram[1361]->outb) vsp
Xsram[1362] sram->in sram[1362]->out sram[1362]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1362]->out) 0
.nodeset V(sram[1362]->outb) vsp
Xsram[1363] sram->in sram[1363]->out sram[1363]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1363]->out) 0
.nodeset V(sram[1363]->outb) vsp
Xsram[1364] sram->in sram[1364]->out sram[1364]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1364]->out) 0
.nodeset V(sram[1364]->outb) vsp
Xsram[1365] sram->in sram[1365]->out sram[1365]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1365]->out) 0
.nodeset V(sram[1365]->outb) vsp
Xsram[1366] sram->in sram[1366]->out sram[1366]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1366]->out) 0
.nodeset V(sram[1366]->outb) vsp
Xsram[1367] sram->in sram[1367]->out sram[1367]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1367]->out) 0
.nodeset V(sram[1367]->outb) vsp
Xsram[1368] sram->in sram[1368]->out sram[1368]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1368]->out) 0
.nodeset V(sram[1368]->outb) vsp
Xsram[1369] sram->in sram[1369]->out sram[1369]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1369]->out) 0
.nodeset V(sram[1369]->outb) vsp
Xmux_2level_size50[45] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[7]->in[3] sram[1370]->outb sram[1370]->out sram[1371]->out sram[1371]->outb sram[1372]->out sram[1372]->outb sram[1373]->out sram[1373]->outb sram[1374]->out sram[1374]->outb sram[1375]->out sram[1375]->outb sram[1376]->out sram[1376]->outb sram[1377]->out sram[1377]->outb sram[1378]->outb sram[1378]->out sram[1379]->out sram[1379]->outb sram[1380]->out sram[1380]->outb sram[1381]->out sram[1381]->outb sram[1382]->out sram[1382]->outb sram[1383]->out sram[1383]->outb sram[1384]->out sram[1384]->outb sram[1385]->out sram[1385]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[45], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1370] sram->in sram[1370]->out sram[1370]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1370]->out) 0
.nodeset V(sram[1370]->outb) vsp
Xsram[1371] sram->in sram[1371]->out sram[1371]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1371]->out) 0
.nodeset V(sram[1371]->outb) vsp
Xsram[1372] sram->in sram[1372]->out sram[1372]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1372]->out) 0
.nodeset V(sram[1372]->outb) vsp
Xsram[1373] sram->in sram[1373]->out sram[1373]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1373]->out) 0
.nodeset V(sram[1373]->outb) vsp
Xsram[1374] sram->in sram[1374]->out sram[1374]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1374]->out) 0
.nodeset V(sram[1374]->outb) vsp
Xsram[1375] sram->in sram[1375]->out sram[1375]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1375]->out) 0
.nodeset V(sram[1375]->outb) vsp
Xsram[1376] sram->in sram[1376]->out sram[1376]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1376]->out) 0
.nodeset V(sram[1376]->outb) vsp
Xsram[1377] sram->in sram[1377]->out sram[1377]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1377]->out) 0
.nodeset V(sram[1377]->outb) vsp
Xsram[1378] sram->in sram[1378]->out sram[1378]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1378]->out) 0
.nodeset V(sram[1378]->outb) vsp
Xsram[1379] sram->in sram[1379]->out sram[1379]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1379]->out) 0
.nodeset V(sram[1379]->outb) vsp
Xsram[1380] sram->in sram[1380]->out sram[1380]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1380]->out) 0
.nodeset V(sram[1380]->outb) vsp
Xsram[1381] sram->in sram[1381]->out sram[1381]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1381]->out) 0
.nodeset V(sram[1381]->outb) vsp
Xsram[1382] sram->in sram[1382]->out sram[1382]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1382]->out) 0
.nodeset V(sram[1382]->outb) vsp
Xsram[1383] sram->in sram[1383]->out sram[1383]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1383]->out) 0
.nodeset V(sram[1383]->outb) vsp
Xsram[1384] sram->in sram[1384]->out sram[1384]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1384]->out) 0
.nodeset V(sram[1384]->outb) vsp
Xsram[1385] sram->in sram[1385]->out sram[1385]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1385]->out) 0
.nodeset V(sram[1385]->outb) vsp
Xmux_2level_size50[46] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[7]->in[4] sram[1386]->outb sram[1386]->out sram[1387]->out sram[1387]->outb sram[1388]->out sram[1388]->outb sram[1389]->out sram[1389]->outb sram[1390]->out sram[1390]->outb sram[1391]->out sram[1391]->outb sram[1392]->out sram[1392]->outb sram[1393]->out sram[1393]->outb sram[1394]->outb sram[1394]->out sram[1395]->out sram[1395]->outb sram[1396]->out sram[1396]->outb sram[1397]->out sram[1397]->outb sram[1398]->out sram[1398]->outb sram[1399]->out sram[1399]->outb sram[1400]->out sram[1400]->outb sram[1401]->out sram[1401]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[46], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1386] sram->in sram[1386]->out sram[1386]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1386]->out) 0
.nodeset V(sram[1386]->outb) vsp
Xsram[1387] sram->in sram[1387]->out sram[1387]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1387]->out) 0
.nodeset V(sram[1387]->outb) vsp
Xsram[1388] sram->in sram[1388]->out sram[1388]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1388]->out) 0
.nodeset V(sram[1388]->outb) vsp
Xsram[1389] sram->in sram[1389]->out sram[1389]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1389]->out) 0
.nodeset V(sram[1389]->outb) vsp
Xsram[1390] sram->in sram[1390]->out sram[1390]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1390]->out) 0
.nodeset V(sram[1390]->outb) vsp
Xsram[1391] sram->in sram[1391]->out sram[1391]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1391]->out) 0
.nodeset V(sram[1391]->outb) vsp
Xsram[1392] sram->in sram[1392]->out sram[1392]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1392]->out) 0
.nodeset V(sram[1392]->outb) vsp
Xsram[1393] sram->in sram[1393]->out sram[1393]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1393]->out) 0
.nodeset V(sram[1393]->outb) vsp
Xsram[1394] sram->in sram[1394]->out sram[1394]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1394]->out) 0
.nodeset V(sram[1394]->outb) vsp
Xsram[1395] sram->in sram[1395]->out sram[1395]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1395]->out) 0
.nodeset V(sram[1395]->outb) vsp
Xsram[1396] sram->in sram[1396]->out sram[1396]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1396]->out) 0
.nodeset V(sram[1396]->outb) vsp
Xsram[1397] sram->in sram[1397]->out sram[1397]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1397]->out) 0
.nodeset V(sram[1397]->outb) vsp
Xsram[1398] sram->in sram[1398]->out sram[1398]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1398]->out) 0
.nodeset V(sram[1398]->outb) vsp
Xsram[1399] sram->in sram[1399]->out sram[1399]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1399]->out) 0
.nodeset V(sram[1399]->outb) vsp
Xsram[1400] sram->in sram[1400]->out sram[1400]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1400]->out) 0
.nodeset V(sram[1400]->outb) vsp
Xsram[1401] sram->in sram[1401]->out sram[1401]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1401]->out) 0
.nodeset V(sram[1401]->outb) vsp
Xmux_2level_size50[47] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[7]->in[5] sram[1402]->outb sram[1402]->out sram[1403]->out sram[1403]->outb sram[1404]->out sram[1404]->outb sram[1405]->out sram[1405]->outb sram[1406]->out sram[1406]->outb sram[1407]->out sram[1407]->outb sram[1408]->out sram[1408]->outb sram[1409]->out sram[1409]->outb sram[1410]->outb sram[1410]->out sram[1411]->out sram[1411]->outb sram[1412]->out sram[1412]->outb sram[1413]->out sram[1413]->outb sram[1414]->out sram[1414]->outb sram[1415]->out sram[1415]->outb sram[1416]->out sram[1416]->outb sram[1417]->out sram[1417]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[47], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1402] sram->in sram[1402]->out sram[1402]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1402]->out) 0
.nodeset V(sram[1402]->outb) vsp
Xsram[1403] sram->in sram[1403]->out sram[1403]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1403]->out) 0
.nodeset V(sram[1403]->outb) vsp
Xsram[1404] sram->in sram[1404]->out sram[1404]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1404]->out) 0
.nodeset V(sram[1404]->outb) vsp
Xsram[1405] sram->in sram[1405]->out sram[1405]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1405]->out) 0
.nodeset V(sram[1405]->outb) vsp
Xsram[1406] sram->in sram[1406]->out sram[1406]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1406]->out) 0
.nodeset V(sram[1406]->outb) vsp
Xsram[1407] sram->in sram[1407]->out sram[1407]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1407]->out) 0
.nodeset V(sram[1407]->outb) vsp
Xsram[1408] sram->in sram[1408]->out sram[1408]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1408]->out) 0
.nodeset V(sram[1408]->outb) vsp
Xsram[1409] sram->in sram[1409]->out sram[1409]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1409]->out) 0
.nodeset V(sram[1409]->outb) vsp
Xsram[1410] sram->in sram[1410]->out sram[1410]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1410]->out) 0
.nodeset V(sram[1410]->outb) vsp
Xsram[1411] sram->in sram[1411]->out sram[1411]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1411]->out) 0
.nodeset V(sram[1411]->outb) vsp
Xsram[1412] sram->in sram[1412]->out sram[1412]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1412]->out) 0
.nodeset V(sram[1412]->outb) vsp
Xsram[1413] sram->in sram[1413]->out sram[1413]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1413]->out) 0
.nodeset V(sram[1413]->outb) vsp
Xsram[1414] sram->in sram[1414]->out sram[1414]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1414]->out) 0
.nodeset V(sram[1414]->outb) vsp
Xsram[1415] sram->in sram[1415]->out sram[1415]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1415]->out) 0
.nodeset V(sram[1415]->outb) vsp
Xsram[1416] sram->in sram[1416]->out sram[1416]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1416]->out) 0
.nodeset V(sram[1416]->outb) vsp
Xsram[1417] sram->in sram[1417]->out sram[1417]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1417]->out) 0
.nodeset V(sram[1417]->outb) vsp
Xdirect_interc[177] mode[clb]->clk[0] fle[7]->clk[0] gvdd_local_interc sgnd direct_interc
Xmux_2level_size50[48] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[8]->in[0] sram[1418]->outb sram[1418]->out sram[1419]->out sram[1419]->outb sram[1420]->out sram[1420]->outb sram[1421]->out sram[1421]->outb sram[1422]->out sram[1422]->outb sram[1423]->out sram[1423]->outb sram[1424]->out sram[1424]->outb sram[1425]->out sram[1425]->outb sram[1426]->outb sram[1426]->out sram[1427]->out sram[1427]->outb sram[1428]->out sram[1428]->outb sram[1429]->out sram[1429]->outb sram[1430]->out sram[1430]->outb sram[1431]->out sram[1431]->outb sram[1432]->out sram[1432]->outb sram[1433]->out sram[1433]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[48], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1418] sram->in sram[1418]->out sram[1418]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1418]->out) 0
.nodeset V(sram[1418]->outb) vsp
Xsram[1419] sram->in sram[1419]->out sram[1419]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1419]->out) 0
.nodeset V(sram[1419]->outb) vsp
Xsram[1420] sram->in sram[1420]->out sram[1420]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1420]->out) 0
.nodeset V(sram[1420]->outb) vsp
Xsram[1421] sram->in sram[1421]->out sram[1421]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1421]->out) 0
.nodeset V(sram[1421]->outb) vsp
Xsram[1422] sram->in sram[1422]->out sram[1422]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1422]->out) 0
.nodeset V(sram[1422]->outb) vsp
Xsram[1423] sram->in sram[1423]->out sram[1423]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1423]->out) 0
.nodeset V(sram[1423]->outb) vsp
Xsram[1424] sram->in sram[1424]->out sram[1424]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1424]->out) 0
.nodeset V(sram[1424]->outb) vsp
Xsram[1425] sram->in sram[1425]->out sram[1425]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1425]->out) 0
.nodeset V(sram[1425]->outb) vsp
Xsram[1426] sram->in sram[1426]->out sram[1426]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1426]->out) 0
.nodeset V(sram[1426]->outb) vsp
Xsram[1427] sram->in sram[1427]->out sram[1427]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1427]->out) 0
.nodeset V(sram[1427]->outb) vsp
Xsram[1428] sram->in sram[1428]->out sram[1428]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1428]->out) 0
.nodeset V(sram[1428]->outb) vsp
Xsram[1429] sram->in sram[1429]->out sram[1429]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1429]->out) 0
.nodeset V(sram[1429]->outb) vsp
Xsram[1430] sram->in sram[1430]->out sram[1430]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1430]->out) 0
.nodeset V(sram[1430]->outb) vsp
Xsram[1431] sram->in sram[1431]->out sram[1431]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1431]->out) 0
.nodeset V(sram[1431]->outb) vsp
Xsram[1432] sram->in sram[1432]->out sram[1432]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1432]->out) 0
.nodeset V(sram[1432]->outb) vsp
Xsram[1433] sram->in sram[1433]->out sram[1433]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1433]->out) 0
.nodeset V(sram[1433]->outb) vsp
Xmux_2level_size50[49] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[8]->in[1] sram[1434]->outb sram[1434]->out sram[1435]->out sram[1435]->outb sram[1436]->out sram[1436]->outb sram[1437]->out sram[1437]->outb sram[1438]->out sram[1438]->outb sram[1439]->out sram[1439]->outb sram[1440]->out sram[1440]->outb sram[1441]->out sram[1441]->outb sram[1442]->outb sram[1442]->out sram[1443]->out sram[1443]->outb sram[1444]->out sram[1444]->outb sram[1445]->out sram[1445]->outb sram[1446]->out sram[1446]->outb sram[1447]->out sram[1447]->outb sram[1448]->out sram[1448]->outb sram[1449]->out sram[1449]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[49], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1434] sram->in sram[1434]->out sram[1434]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1434]->out) 0
.nodeset V(sram[1434]->outb) vsp
Xsram[1435] sram->in sram[1435]->out sram[1435]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1435]->out) 0
.nodeset V(sram[1435]->outb) vsp
Xsram[1436] sram->in sram[1436]->out sram[1436]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1436]->out) 0
.nodeset V(sram[1436]->outb) vsp
Xsram[1437] sram->in sram[1437]->out sram[1437]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1437]->out) 0
.nodeset V(sram[1437]->outb) vsp
Xsram[1438] sram->in sram[1438]->out sram[1438]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1438]->out) 0
.nodeset V(sram[1438]->outb) vsp
Xsram[1439] sram->in sram[1439]->out sram[1439]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1439]->out) 0
.nodeset V(sram[1439]->outb) vsp
Xsram[1440] sram->in sram[1440]->out sram[1440]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1440]->out) 0
.nodeset V(sram[1440]->outb) vsp
Xsram[1441] sram->in sram[1441]->out sram[1441]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1441]->out) 0
.nodeset V(sram[1441]->outb) vsp
Xsram[1442] sram->in sram[1442]->out sram[1442]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1442]->out) 0
.nodeset V(sram[1442]->outb) vsp
Xsram[1443] sram->in sram[1443]->out sram[1443]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1443]->out) 0
.nodeset V(sram[1443]->outb) vsp
Xsram[1444] sram->in sram[1444]->out sram[1444]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1444]->out) 0
.nodeset V(sram[1444]->outb) vsp
Xsram[1445] sram->in sram[1445]->out sram[1445]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1445]->out) 0
.nodeset V(sram[1445]->outb) vsp
Xsram[1446] sram->in sram[1446]->out sram[1446]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1446]->out) 0
.nodeset V(sram[1446]->outb) vsp
Xsram[1447] sram->in sram[1447]->out sram[1447]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1447]->out) 0
.nodeset V(sram[1447]->outb) vsp
Xsram[1448] sram->in sram[1448]->out sram[1448]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1448]->out) 0
.nodeset V(sram[1448]->outb) vsp
Xsram[1449] sram->in sram[1449]->out sram[1449]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1449]->out) 0
.nodeset V(sram[1449]->outb) vsp
Xmux_2level_size50[50] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[8]->in[2] sram[1450]->outb sram[1450]->out sram[1451]->out sram[1451]->outb sram[1452]->out sram[1452]->outb sram[1453]->out sram[1453]->outb sram[1454]->out sram[1454]->outb sram[1455]->out sram[1455]->outb sram[1456]->out sram[1456]->outb sram[1457]->out sram[1457]->outb sram[1458]->outb sram[1458]->out sram[1459]->out sram[1459]->outb sram[1460]->out sram[1460]->outb sram[1461]->out sram[1461]->outb sram[1462]->out sram[1462]->outb sram[1463]->out sram[1463]->outb sram[1464]->out sram[1464]->outb sram[1465]->out sram[1465]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[50], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1450] sram->in sram[1450]->out sram[1450]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1450]->out) 0
.nodeset V(sram[1450]->outb) vsp
Xsram[1451] sram->in sram[1451]->out sram[1451]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1451]->out) 0
.nodeset V(sram[1451]->outb) vsp
Xsram[1452] sram->in sram[1452]->out sram[1452]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1452]->out) 0
.nodeset V(sram[1452]->outb) vsp
Xsram[1453] sram->in sram[1453]->out sram[1453]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1453]->out) 0
.nodeset V(sram[1453]->outb) vsp
Xsram[1454] sram->in sram[1454]->out sram[1454]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1454]->out) 0
.nodeset V(sram[1454]->outb) vsp
Xsram[1455] sram->in sram[1455]->out sram[1455]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1455]->out) 0
.nodeset V(sram[1455]->outb) vsp
Xsram[1456] sram->in sram[1456]->out sram[1456]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1456]->out) 0
.nodeset V(sram[1456]->outb) vsp
Xsram[1457] sram->in sram[1457]->out sram[1457]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1457]->out) 0
.nodeset V(sram[1457]->outb) vsp
Xsram[1458] sram->in sram[1458]->out sram[1458]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1458]->out) 0
.nodeset V(sram[1458]->outb) vsp
Xsram[1459] sram->in sram[1459]->out sram[1459]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1459]->out) 0
.nodeset V(sram[1459]->outb) vsp
Xsram[1460] sram->in sram[1460]->out sram[1460]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1460]->out) 0
.nodeset V(sram[1460]->outb) vsp
Xsram[1461] sram->in sram[1461]->out sram[1461]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1461]->out) 0
.nodeset V(sram[1461]->outb) vsp
Xsram[1462] sram->in sram[1462]->out sram[1462]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1462]->out) 0
.nodeset V(sram[1462]->outb) vsp
Xsram[1463] sram->in sram[1463]->out sram[1463]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1463]->out) 0
.nodeset V(sram[1463]->outb) vsp
Xsram[1464] sram->in sram[1464]->out sram[1464]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1464]->out) 0
.nodeset V(sram[1464]->outb) vsp
Xsram[1465] sram->in sram[1465]->out sram[1465]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1465]->out) 0
.nodeset V(sram[1465]->outb) vsp
Xmux_2level_size50[51] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[8]->in[3] sram[1466]->outb sram[1466]->out sram[1467]->out sram[1467]->outb sram[1468]->out sram[1468]->outb sram[1469]->out sram[1469]->outb sram[1470]->out sram[1470]->outb sram[1471]->out sram[1471]->outb sram[1472]->out sram[1472]->outb sram[1473]->out sram[1473]->outb sram[1474]->outb sram[1474]->out sram[1475]->out sram[1475]->outb sram[1476]->out sram[1476]->outb sram[1477]->out sram[1477]->outb sram[1478]->out sram[1478]->outb sram[1479]->out sram[1479]->outb sram[1480]->out sram[1480]->outb sram[1481]->out sram[1481]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[51], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1466] sram->in sram[1466]->out sram[1466]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1466]->out) 0
.nodeset V(sram[1466]->outb) vsp
Xsram[1467] sram->in sram[1467]->out sram[1467]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1467]->out) 0
.nodeset V(sram[1467]->outb) vsp
Xsram[1468] sram->in sram[1468]->out sram[1468]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1468]->out) 0
.nodeset V(sram[1468]->outb) vsp
Xsram[1469] sram->in sram[1469]->out sram[1469]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1469]->out) 0
.nodeset V(sram[1469]->outb) vsp
Xsram[1470] sram->in sram[1470]->out sram[1470]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1470]->out) 0
.nodeset V(sram[1470]->outb) vsp
Xsram[1471] sram->in sram[1471]->out sram[1471]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1471]->out) 0
.nodeset V(sram[1471]->outb) vsp
Xsram[1472] sram->in sram[1472]->out sram[1472]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1472]->out) 0
.nodeset V(sram[1472]->outb) vsp
Xsram[1473] sram->in sram[1473]->out sram[1473]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1473]->out) 0
.nodeset V(sram[1473]->outb) vsp
Xsram[1474] sram->in sram[1474]->out sram[1474]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1474]->out) 0
.nodeset V(sram[1474]->outb) vsp
Xsram[1475] sram->in sram[1475]->out sram[1475]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1475]->out) 0
.nodeset V(sram[1475]->outb) vsp
Xsram[1476] sram->in sram[1476]->out sram[1476]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1476]->out) 0
.nodeset V(sram[1476]->outb) vsp
Xsram[1477] sram->in sram[1477]->out sram[1477]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1477]->out) 0
.nodeset V(sram[1477]->outb) vsp
Xsram[1478] sram->in sram[1478]->out sram[1478]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1478]->out) 0
.nodeset V(sram[1478]->outb) vsp
Xsram[1479] sram->in sram[1479]->out sram[1479]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1479]->out) 0
.nodeset V(sram[1479]->outb) vsp
Xsram[1480] sram->in sram[1480]->out sram[1480]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1480]->out) 0
.nodeset V(sram[1480]->outb) vsp
Xsram[1481] sram->in sram[1481]->out sram[1481]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1481]->out) 0
.nodeset V(sram[1481]->outb) vsp
Xmux_2level_size50[52] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[8]->in[4] sram[1482]->outb sram[1482]->out sram[1483]->out sram[1483]->outb sram[1484]->out sram[1484]->outb sram[1485]->out sram[1485]->outb sram[1486]->out sram[1486]->outb sram[1487]->out sram[1487]->outb sram[1488]->out sram[1488]->outb sram[1489]->out sram[1489]->outb sram[1490]->outb sram[1490]->out sram[1491]->out sram[1491]->outb sram[1492]->out sram[1492]->outb sram[1493]->out sram[1493]->outb sram[1494]->out sram[1494]->outb sram[1495]->out sram[1495]->outb sram[1496]->out sram[1496]->outb sram[1497]->out sram[1497]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[52], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1482] sram->in sram[1482]->out sram[1482]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1482]->out) 0
.nodeset V(sram[1482]->outb) vsp
Xsram[1483] sram->in sram[1483]->out sram[1483]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1483]->out) 0
.nodeset V(sram[1483]->outb) vsp
Xsram[1484] sram->in sram[1484]->out sram[1484]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1484]->out) 0
.nodeset V(sram[1484]->outb) vsp
Xsram[1485] sram->in sram[1485]->out sram[1485]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1485]->out) 0
.nodeset V(sram[1485]->outb) vsp
Xsram[1486] sram->in sram[1486]->out sram[1486]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1486]->out) 0
.nodeset V(sram[1486]->outb) vsp
Xsram[1487] sram->in sram[1487]->out sram[1487]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1487]->out) 0
.nodeset V(sram[1487]->outb) vsp
Xsram[1488] sram->in sram[1488]->out sram[1488]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1488]->out) 0
.nodeset V(sram[1488]->outb) vsp
Xsram[1489] sram->in sram[1489]->out sram[1489]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1489]->out) 0
.nodeset V(sram[1489]->outb) vsp
Xsram[1490] sram->in sram[1490]->out sram[1490]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1490]->out) 0
.nodeset V(sram[1490]->outb) vsp
Xsram[1491] sram->in sram[1491]->out sram[1491]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1491]->out) 0
.nodeset V(sram[1491]->outb) vsp
Xsram[1492] sram->in sram[1492]->out sram[1492]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1492]->out) 0
.nodeset V(sram[1492]->outb) vsp
Xsram[1493] sram->in sram[1493]->out sram[1493]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1493]->out) 0
.nodeset V(sram[1493]->outb) vsp
Xsram[1494] sram->in sram[1494]->out sram[1494]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1494]->out) 0
.nodeset V(sram[1494]->outb) vsp
Xsram[1495] sram->in sram[1495]->out sram[1495]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1495]->out) 0
.nodeset V(sram[1495]->outb) vsp
Xsram[1496] sram->in sram[1496]->out sram[1496]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1496]->out) 0
.nodeset V(sram[1496]->outb) vsp
Xsram[1497] sram->in sram[1497]->out sram[1497]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1497]->out) 0
.nodeset V(sram[1497]->outb) vsp
Xmux_2level_size50[53] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[8]->in[5] sram[1498]->outb sram[1498]->out sram[1499]->out sram[1499]->outb sram[1500]->out sram[1500]->outb sram[1501]->out sram[1501]->outb sram[1502]->out sram[1502]->outb sram[1503]->out sram[1503]->outb sram[1504]->out sram[1504]->outb sram[1505]->out sram[1505]->outb sram[1506]->outb sram[1506]->out sram[1507]->out sram[1507]->outb sram[1508]->out sram[1508]->outb sram[1509]->out sram[1509]->outb sram[1510]->out sram[1510]->outb sram[1511]->out sram[1511]->outb sram[1512]->out sram[1512]->outb sram[1513]->out sram[1513]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[53], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1498] sram->in sram[1498]->out sram[1498]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1498]->out) 0
.nodeset V(sram[1498]->outb) vsp
Xsram[1499] sram->in sram[1499]->out sram[1499]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1499]->out) 0
.nodeset V(sram[1499]->outb) vsp
Xsram[1500] sram->in sram[1500]->out sram[1500]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1500]->out) 0
.nodeset V(sram[1500]->outb) vsp
Xsram[1501] sram->in sram[1501]->out sram[1501]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1501]->out) 0
.nodeset V(sram[1501]->outb) vsp
Xsram[1502] sram->in sram[1502]->out sram[1502]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1502]->out) 0
.nodeset V(sram[1502]->outb) vsp
Xsram[1503] sram->in sram[1503]->out sram[1503]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1503]->out) 0
.nodeset V(sram[1503]->outb) vsp
Xsram[1504] sram->in sram[1504]->out sram[1504]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1504]->out) 0
.nodeset V(sram[1504]->outb) vsp
Xsram[1505] sram->in sram[1505]->out sram[1505]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1505]->out) 0
.nodeset V(sram[1505]->outb) vsp
Xsram[1506] sram->in sram[1506]->out sram[1506]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1506]->out) 0
.nodeset V(sram[1506]->outb) vsp
Xsram[1507] sram->in sram[1507]->out sram[1507]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1507]->out) 0
.nodeset V(sram[1507]->outb) vsp
Xsram[1508] sram->in sram[1508]->out sram[1508]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1508]->out) 0
.nodeset V(sram[1508]->outb) vsp
Xsram[1509] sram->in sram[1509]->out sram[1509]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1509]->out) 0
.nodeset V(sram[1509]->outb) vsp
Xsram[1510] sram->in sram[1510]->out sram[1510]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1510]->out) 0
.nodeset V(sram[1510]->outb) vsp
Xsram[1511] sram->in sram[1511]->out sram[1511]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1511]->out) 0
.nodeset V(sram[1511]->outb) vsp
Xsram[1512] sram->in sram[1512]->out sram[1512]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1512]->out) 0
.nodeset V(sram[1512]->outb) vsp
Xsram[1513] sram->in sram[1513]->out sram[1513]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1513]->out) 0
.nodeset V(sram[1513]->outb) vsp
Xdirect_interc[178] mode[clb]->clk[0] fle[8]->clk[0] gvdd_local_interc sgnd direct_interc
Xmux_2level_size50[54] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[9]->in[0] sram[1514]->out sram[1514]->outb sram[1515]->out sram[1515]->outb sram[1516]->outb sram[1516]->out sram[1517]->out sram[1517]->outb sram[1518]->out sram[1518]->outb sram[1519]->out sram[1519]->outb sram[1520]->out sram[1520]->outb sram[1521]->out sram[1521]->outb sram[1522]->out sram[1522]->outb sram[1523]->out sram[1523]->outb sram[1524]->out sram[1524]->outb sram[1525]->out sram[1525]->outb sram[1526]->out sram[1526]->outb sram[1527]->out sram[1527]->outb sram[1528]->outb sram[1528]->out sram[1529]->out sram[1529]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[54], level=2, select_path_id=22. *****
*****0010000000000010*****
Xsram[1514] sram->in sram[1514]->out sram[1514]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1514]->out) 0
.nodeset V(sram[1514]->outb) vsp
Xsram[1515] sram->in sram[1515]->out sram[1515]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1515]->out) 0
.nodeset V(sram[1515]->outb) vsp
Xsram[1516] sram->in sram[1516]->out sram[1516]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1516]->out) 0
.nodeset V(sram[1516]->outb) vsp
Xsram[1517] sram->in sram[1517]->out sram[1517]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1517]->out) 0
.nodeset V(sram[1517]->outb) vsp
Xsram[1518] sram->in sram[1518]->out sram[1518]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1518]->out) 0
.nodeset V(sram[1518]->outb) vsp
Xsram[1519] sram->in sram[1519]->out sram[1519]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1519]->out) 0
.nodeset V(sram[1519]->outb) vsp
Xsram[1520] sram->in sram[1520]->out sram[1520]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1520]->out) 0
.nodeset V(sram[1520]->outb) vsp
Xsram[1521] sram->in sram[1521]->out sram[1521]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1521]->out) 0
.nodeset V(sram[1521]->outb) vsp
Xsram[1522] sram->in sram[1522]->out sram[1522]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1522]->out) 0
.nodeset V(sram[1522]->outb) vsp
Xsram[1523] sram->in sram[1523]->out sram[1523]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1523]->out) 0
.nodeset V(sram[1523]->outb) vsp
Xsram[1524] sram->in sram[1524]->out sram[1524]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1524]->out) 0
.nodeset V(sram[1524]->outb) vsp
Xsram[1525] sram->in sram[1525]->out sram[1525]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1525]->out) 0
.nodeset V(sram[1525]->outb) vsp
Xsram[1526] sram->in sram[1526]->out sram[1526]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1526]->out) 0
.nodeset V(sram[1526]->outb) vsp
Xsram[1527] sram->in sram[1527]->out sram[1527]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1527]->out) 0
.nodeset V(sram[1527]->outb) vsp
Xsram[1528] sram->in sram[1528]->out sram[1528]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1528]->out) 0
.nodeset V(sram[1528]->outb) vsp
Xsram[1529] sram->in sram[1529]->out sram[1529]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1529]->out) 0
.nodeset V(sram[1529]->outb) vsp
Xmux_2level_size50[55] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[9]->in[1] sram[1530]->outb sram[1530]->out sram[1531]->out sram[1531]->outb sram[1532]->out sram[1532]->outb sram[1533]->out sram[1533]->outb sram[1534]->out sram[1534]->outb sram[1535]->out sram[1535]->outb sram[1536]->out sram[1536]->outb sram[1537]->out sram[1537]->outb sram[1538]->outb sram[1538]->out sram[1539]->out sram[1539]->outb sram[1540]->out sram[1540]->outb sram[1541]->out sram[1541]->outb sram[1542]->out sram[1542]->outb sram[1543]->out sram[1543]->outb sram[1544]->out sram[1544]->outb sram[1545]->out sram[1545]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[55], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1530] sram->in sram[1530]->out sram[1530]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1530]->out) 0
.nodeset V(sram[1530]->outb) vsp
Xsram[1531] sram->in sram[1531]->out sram[1531]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1531]->out) 0
.nodeset V(sram[1531]->outb) vsp
Xsram[1532] sram->in sram[1532]->out sram[1532]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1532]->out) 0
.nodeset V(sram[1532]->outb) vsp
Xsram[1533] sram->in sram[1533]->out sram[1533]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1533]->out) 0
.nodeset V(sram[1533]->outb) vsp
Xsram[1534] sram->in sram[1534]->out sram[1534]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1534]->out) 0
.nodeset V(sram[1534]->outb) vsp
Xsram[1535] sram->in sram[1535]->out sram[1535]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1535]->out) 0
.nodeset V(sram[1535]->outb) vsp
Xsram[1536] sram->in sram[1536]->out sram[1536]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1536]->out) 0
.nodeset V(sram[1536]->outb) vsp
Xsram[1537] sram->in sram[1537]->out sram[1537]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1537]->out) 0
.nodeset V(sram[1537]->outb) vsp
Xsram[1538] sram->in sram[1538]->out sram[1538]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1538]->out) 0
.nodeset V(sram[1538]->outb) vsp
Xsram[1539] sram->in sram[1539]->out sram[1539]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1539]->out) 0
.nodeset V(sram[1539]->outb) vsp
Xsram[1540] sram->in sram[1540]->out sram[1540]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1540]->out) 0
.nodeset V(sram[1540]->outb) vsp
Xsram[1541] sram->in sram[1541]->out sram[1541]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1541]->out) 0
.nodeset V(sram[1541]->outb) vsp
Xsram[1542] sram->in sram[1542]->out sram[1542]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1542]->out) 0
.nodeset V(sram[1542]->outb) vsp
Xsram[1543] sram->in sram[1543]->out sram[1543]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1543]->out) 0
.nodeset V(sram[1543]->outb) vsp
Xsram[1544] sram->in sram[1544]->out sram[1544]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1544]->out) 0
.nodeset V(sram[1544]->outb) vsp
Xsram[1545] sram->in sram[1545]->out sram[1545]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1545]->out) 0
.nodeset V(sram[1545]->outb) vsp
Xmux_2level_size50[56] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[9]->in[2] sram[1546]->outb sram[1546]->out sram[1547]->out sram[1547]->outb sram[1548]->out sram[1548]->outb sram[1549]->out sram[1549]->outb sram[1550]->out sram[1550]->outb sram[1551]->out sram[1551]->outb sram[1552]->out sram[1552]->outb sram[1553]->out sram[1553]->outb sram[1554]->outb sram[1554]->out sram[1555]->out sram[1555]->outb sram[1556]->out sram[1556]->outb sram[1557]->out sram[1557]->outb sram[1558]->out sram[1558]->outb sram[1559]->out sram[1559]->outb sram[1560]->out sram[1560]->outb sram[1561]->out sram[1561]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[56], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1546] sram->in sram[1546]->out sram[1546]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1546]->out) 0
.nodeset V(sram[1546]->outb) vsp
Xsram[1547] sram->in sram[1547]->out sram[1547]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1547]->out) 0
.nodeset V(sram[1547]->outb) vsp
Xsram[1548] sram->in sram[1548]->out sram[1548]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1548]->out) 0
.nodeset V(sram[1548]->outb) vsp
Xsram[1549] sram->in sram[1549]->out sram[1549]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1549]->out) 0
.nodeset V(sram[1549]->outb) vsp
Xsram[1550] sram->in sram[1550]->out sram[1550]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1550]->out) 0
.nodeset V(sram[1550]->outb) vsp
Xsram[1551] sram->in sram[1551]->out sram[1551]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1551]->out) 0
.nodeset V(sram[1551]->outb) vsp
Xsram[1552] sram->in sram[1552]->out sram[1552]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1552]->out) 0
.nodeset V(sram[1552]->outb) vsp
Xsram[1553] sram->in sram[1553]->out sram[1553]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1553]->out) 0
.nodeset V(sram[1553]->outb) vsp
Xsram[1554] sram->in sram[1554]->out sram[1554]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1554]->out) 0
.nodeset V(sram[1554]->outb) vsp
Xsram[1555] sram->in sram[1555]->out sram[1555]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1555]->out) 0
.nodeset V(sram[1555]->outb) vsp
Xsram[1556] sram->in sram[1556]->out sram[1556]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1556]->out) 0
.nodeset V(sram[1556]->outb) vsp
Xsram[1557] sram->in sram[1557]->out sram[1557]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1557]->out) 0
.nodeset V(sram[1557]->outb) vsp
Xsram[1558] sram->in sram[1558]->out sram[1558]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1558]->out) 0
.nodeset V(sram[1558]->outb) vsp
Xsram[1559] sram->in sram[1559]->out sram[1559]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1559]->out) 0
.nodeset V(sram[1559]->outb) vsp
Xsram[1560] sram->in sram[1560]->out sram[1560]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1560]->out) 0
.nodeset V(sram[1560]->outb) vsp
Xsram[1561] sram->in sram[1561]->out sram[1561]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1561]->out) 0
.nodeset V(sram[1561]->outb) vsp
Xmux_2level_size50[57] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[9]->in[3] sram[1562]->outb sram[1562]->out sram[1563]->out sram[1563]->outb sram[1564]->out sram[1564]->outb sram[1565]->out sram[1565]->outb sram[1566]->out sram[1566]->outb sram[1567]->out sram[1567]->outb sram[1568]->out sram[1568]->outb sram[1569]->out sram[1569]->outb sram[1570]->outb sram[1570]->out sram[1571]->out sram[1571]->outb sram[1572]->out sram[1572]->outb sram[1573]->out sram[1573]->outb sram[1574]->out sram[1574]->outb sram[1575]->out sram[1575]->outb sram[1576]->out sram[1576]->outb sram[1577]->out sram[1577]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[57], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1562] sram->in sram[1562]->out sram[1562]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1562]->out) 0
.nodeset V(sram[1562]->outb) vsp
Xsram[1563] sram->in sram[1563]->out sram[1563]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1563]->out) 0
.nodeset V(sram[1563]->outb) vsp
Xsram[1564] sram->in sram[1564]->out sram[1564]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1564]->out) 0
.nodeset V(sram[1564]->outb) vsp
Xsram[1565] sram->in sram[1565]->out sram[1565]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1565]->out) 0
.nodeset V(sram[1565]->outb) vsp
Xsram[1566] sram->in sram[1566]->out sram[1566]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1566]->out) 0
.nodeset V(sram[1566]->outb) vsp
Xsram[1567] sram->in sram[1567]->out sram[1567]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1567]->out) 0
.nodeset V(sram[1567]->outb) vsp
Xsram[1568] sram->in sram[1568]->out sram[1568]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1568]->out) 0
.nodeset V(sram[1568]->outb) vsp
Xsram[1569] sram->in sram[1569]->out sram[1569]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1569]->out) 0
.nodeset V(sram[1569]->outb) vsp
Xsram[1570] sram->in sram[1570]->out sram[1570]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1570]->out) 0
.nodeset V(sram[1570]->outb) vsp
Xsram[1571] sram->in sram[1571]->out sram[1571]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1571]->out) 0
.nodeset V(sram[1571]->outb) vsp
Xsram[1572] sram->in sram[1572]->out sram[1572]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1572]->out) 0
.nodeset V(sram[1572]->outb) vsp
Xsram[1573] sram->in sram[1573]->out sram[1573]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1573]->out) 0
.nodeset V(sram[1573]->outb) vsp
Xsram[1574] sram->in sram[1574]->out sram[1574]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1574]->out) 0
.nodeset V(sram[1574]->outb) vsp
Xsram[1575] sram->in sram[1575]->out sram[1575]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1575]->out) 0
.nodeset V(sram[1575]->outb) vsp
Xsram[1576] sram->in sram[1576]->out sram[1576]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1576]->out) 0
.nodeset V(sram[1576]->outb) vsp
Xsram[1577] sram->in sram[1577]->out sram[1577]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1577]->out) 0
.nodeset V(sram[1577]->outb) vsp
Xmux_2level_size50[58] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[9]->in[4] sram[1578]->outb sram[1578]->out sram[1579]->out sram[1579]->outb sram[1580]->out sram[1580]->outb sram[1581]->out sram[1581]->outb sram[1582]->out sram[1582]->outb sram[1583]->out sram[1583]->outb sram[1584]->out sram[1584]->outb sram[1585]->out sram[1585]->outb sram[1586]->outb sram[1586]->out sram[1587]->out sram[1587]->outb sram[1588]->out sram[1588]->outb sram[1589]->out sram[1589]->outb sram[1590]->out sram[1590]->outb sram[1591]->out sram[1591]->outb sram[1592]->out sram[1592]->outb sram[1593]->out sram[1593]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[58], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1578] sram->in sram[1578]->out sram[1578]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1578]->out) 0
.nodeset V(sram[1578]->outb) vsp
Xsram[1579] sram->in sram[1579]->out sram[1579]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1579]->out) 0
.nodeset V(sram[1579]->outb) vsp
Xsram[1580] sram->in sram[1580]->out sram[1580]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1580]->out) 0
.nodeset V(sram[1580]->outb) vsp
Xsram[1581] sram->in sram[1581]->out sram[1581]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1581]->out) 0
.nodeset V(sram[1581]->outb) vsp
Xsram[1582] sram->in sram[1582]->out sram[1582]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1582]->out) 0
.nodeset V(sram[1582]->outb) vsp
Xsram[1583] sram->in sram[1583]->out sram[1583]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1583]->out) 0
.nodeset V(sram[1583]->outb) vsp
Xsram[1584] sram->in sram[1584]->out sram[1584]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1584]->out) 0
.nodeset V(sram[1584]->outb) vsp
Xsram[1585] sram->in sram[1585]->out sram[1585]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1585]->out) 0
.nodeset V(sram[1585]->outb) vsp
Xsram[1586] sram->in sram[1586]->out sram[1586]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1586]->out) 0
.nodeset V(sram[1586]->outb) vsp
Xsram[1587] sram->in sram[1587]->out sram[1587]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1587]->out) 0
.nodeset V(sram[1587]->outb) vsp
Xsram[1588] sram->in sram[1588]->out sram[1588]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1588]->out) 0
.nodeset V(sram[1588]->outb) vsp
Xsram[1589] sram->in sram[1589]->out sram[1589]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1589]->out) 0
.nodeset V(sram[1589]->outb) vsp
Xsram[1590] sram->in sram[1590]->out sram[1590]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1590]->out) 0
.nodeset V(sram[1590]->outb) vsp
Xsram[1591] sram->in sram[1591]->out sram[1591]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1591]->out) 0
.nodeset V(sram[1591]->outb) vsp
Xsram[1592] sram->in sram[1592]->out sram[1592]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1592]->out) 0
.nodeset V(sram[1592]->outb) vsp
Xsram[1593] sram->in sram[1593]->out sram[1593]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1593]->out) 0
.nodeset V(sram[1593]->outb) vsp
Xmux_2level_size50[59] mode[clb]->I[0] mode[clb]->I[1] mode[clb]->I[2] mode[clb]->I[3] mode[clb]->I[4] mode[clb]->I[5] mode[clb]->I[6] mode[clb]->I[7] mode[clb]->I[8] mode[clb]->I[9] mode[clb]->I[10] mode[clb]->I[11] mode[clb]->I[12] mode[clb]->I[13] mode[clb]->I[14] mode[clb]->I[15] mode[clb]->I[16] mode[clb]->I[17] mode[clb]->I[18] mode[clb]->I[19] mode[clb]->I[20] mode[clb]->I[21] mode[clb]->I[22] mode[clb]->I[23] mode[clb]->I[24] mode[clb]->I[25] mode[clb]->I[26] mode[clb]->I[27] mode[clb]->I[28] mode[clb]->I[29] mode[clb]->I[30] mode[clb]->I[31] mode[clb]->I[32] mode[clb]->I[33] mode[clb]->I[34] mode[clb]->I[35] mode[clb]->I[36] mode[clb]->I[37] mode[clb]->I[38] mode[clb]->I[39] fle[0]->out[0] fle[1]->out[0] fle[2]->out[0] fle[3]->out[0] fle[4]->out[0] fle[5]->out[0] fle[6]->out[0] fle[7]->out[0] fle[8]->out[0] fle[9]->out[0] fle[9]->in[5] sram[1594]->outb sram[1594]->out sram[1595]->out sram[1595]->outb sram[1596]->out sram[1596]->outb sram[1597]->out sram[1597]->outb sram[1598]->out sram[1598]->outb sram[1599]->out sram[1599]->outb sram[1600]->out sram[1600]->outb sram[1601]->out sram[1601]->outb sram[1602]->outb sram[1602]->out sram[1603]->out sram[1603]->outb sram[1604]->out sram[1604]->outb sram[1605]->out sram[1605]->outb sram[1606]->out sram[1606]->outb sram[1607]->out sram[1607]->outb sram[1608]->out sram[1608]->outb sram[1609]->out sram[1609]->outb gvdd_local_interc sgnd mux_2level_size50
***** SRAM bits for MUX[59], level=2, select_path_id=0. *****
*****1000000010000000*****
Xsram[1594] sram->in sram[1594]->out sram[1594]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1594]->out) 0
.nodeset V(sram[1594]->outb) vsp
Xsram[1595] sram->in sram[1595]->out sram[1595]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1595]->out) 0
.nodeset V(sram[1595]->outb) vsp
Xsram[1596] sram->in sram[1596]->out sram[1596]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1596]->out) 0
.nodeset V(sram[1596]->outb) vsp
Xsram[1597] sram->in sram[1597]->out sram[1597]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1597]->out) 0
.nodeset V(sram[1597]->outb) vsp
Xsram[1598] sram->in sram[1598]->out sram[1598]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1598]->out) 0
.nodeset V(sram[1598]->outb) vsp
Xsram[1599] sram->in sram[1599]->out sram[1599]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1599]->out) 0
.nodeset V(sram[1599]->outb) vsp
Xsram[1600] sram->in sram[1600]->out sram[1600]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1600]->out) 0
.nodeset V(sram[1600]->outb) vsp
Xsram[1601] sram->in sram[1601]->out sram[1601]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1601]->out) 0
.nodeset V(sram[1601]->outb) vsp
Xsram[1602] sram->in sram[1602]->out sram[1602]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1602]->out) 0
.nodeset V(sram[1602]->outb) vsp
Xsram[1603] sram->in sram[1603]->out sram[1603]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1603]->out) 0
.nodeset V(sram[1603]->outb) vsp
Xsram[1604] sram->in sram[1604]->out sram[1604]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1604]->out) 0
.nodeset V(sram[1604]->outb) vsp
Xsram[1605] sram->in sram[1605]->out sram[1605]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1605]->out) 0
.nodeset V(sram[1605]->outb) vsp
Xsram[1606] sram->in sram[1606]->out sram[1606]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1606]->out) 0
.nodeset V(sram[1606]->outb) vsp
Xsram[1607] sram->in sram[1607]->out sram[1607]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1607]->out) 0
.nodeset V(sram[1607]->outb) vsp
Xsram[1608] sram->in sram[1608]->out sram[1608]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1608]->out) 0
.nodeset V(sram[1608]->outb) vsp
Xsram[1609] sram->in sram[1609]->out sram[1609]->outb gvdd_sram_local_routing sgnd  sram6T
.nodeset V(sram[1609]->out) 0
.nodeset V(sram[1609]->outb) vsp
Xdirect_interc[179] mode[clb]->clk[0] fle[9]->clk[0] gvdd_local_interc sgnd direct_interc
.eom
***** END *****

***** Grid[1][1], Capactity: 1 *****
***** Top Protocol *****
.subckt grid[1][1] 
+ top_height[0]_pin[0] 
+ top_height[0]_pin[4] 
+ top_height[0]_pin[8] 
+ top_height[0]_pin[12] 
+ top_height[0]_pin[16] 
+ top_height[0]_pin[20] 
+ top_height[0]_pin[24] 
+ top_height[0]_pin[28] 
+ top_height[0]_pin[32] 
+ top_height[0]_pin[36] 
+ top_height[0]_pin[40] 
+ top_height[0]_pin[44] 
+ top_height[0]_pin[48] 
+ right_height[0]_pin[1] 
+ right_height[0]_pin[5] 
+ right_height[0]_pin[9] 
+ right_height[0]_pin[13] 
+ right_height[0]_pin[17] 
+ right_height[0]_pin[21] 
+ right_height[0]_pin[25] 
+ right_height[0]_pin[29] 
+ right_height[0]_pin[33] 
+ right_height[0]_pin[37] 
+ right_height[0]_pin[41] 
+ right_height[0]_pin[45] 
+ right_height[0]_pin[49] 
+ bottom_height[0]_pin[2] 
+ bottom_height[0]_pin[6] 
+ bottom_height[0]_pin[10] 
+ bottom_height[0]_pin[14] 
+ bottom_height[0]_pin[18] 
+ bottom_height[0]_pin[22] 
+ bottom_height[0]_pin[26] 
+ bottom_height[0]_pin[30] 
+ bottom_height[0]_pin[34] 
+ bottom_height[0]_pin[38] 
+ bottom_height[0]_pin[42] 
+ bottom_height[0]_pin[46] 
+ bottom_height[0]_pin[50] 
+ left_height[0]_pin[3] 
+ left_height[0]_pin[7] 
+ left_height[0]_pin[11] 
+ left_height[0]_pin[15] 
+ left_height[0]_pin[19] 
+ left_height[0]_pin[23] 
+ left_height[0]_pin[27] 
+ left_height[0]_pin[31] 
+ left_height[0]_pin[35] 
+ left_height[0]_pin[39] 
+ left_height[0]_pin[43] 
+ left_height[0]_pin[47] 
+ svdd sgnd
Xgrid[1][1][0] 
+ top_height[0]_pin[0] 
+ right_height[0]_pin[1] 
+ bottom_height[0]_pin[2] 
+ left_height[0]_pin[3] 
+ top_height[0]_pin[4] 
+ right_height[0]_pin[5] 
+ bottom_height[0]_pin[6] 
+ left_height[0]_pin[7] 
+ top_height[0]_pin[8] 
+ right_height[0]_pin[9] 
+ bottom_height[0]_pin[10] 
+ left_height[0]_pin[11] 
+ top_height[0]_pin[12] 
+ right_height[0]_pin[13] 
+ bottom_height[0]_pin[14] 
+ left_height[0]_pin[15] 
+ top_height[0]_pin[16] 
+ right_height[0]_pin[17] 
+ bottom_height[0]_pin[18] 
+ left_height[0]_pin[19] 
+ top_height[0]_pin[20] 
+ right_height[0]_pin[21] 
+ bottom_height[0]_pin[22] 
+ left_height[0]_pin[23] 
+ top_height[0]_pin[24] 
+ right_height[0]_pin[25] 
+ bottom_height[0]_pin[26] 
+ left_height[0]_pin[27] 
+ top_height[0]_pin[28] 
+ right_height[0]_pin[29] 
+ bottom_height[0]_pin[30] 
+ left_height[0]_pin[31] 
+ top_height[0]_pin[32] 
+ right_height[0]_pin[33] 
+ bottom_height[0]_pin[34] 
+ left_height[0]_pin[35] 
+ top_height[0]_pin[36] 
+ right_height[0]_pin[37] 
+ bottom_height[0]_pin[38] 
+ left_height[0]_pin[39] 
+ top_height[0]_pin[40] 
+ right_height[0]_pin[41] 
+ bottom_height[0]_pin[42] 
+ left_height[0]_pin[43] 
+ top_height[0]_pin[44] 
+ right_height[0]_pin[45] 
+ bottom_height[0]_pin[46] 
+ left_height[0]_pin[47] 
+ top_height[0]_pin[48] 
+ right_height[0]_pin[49] 
+ bottom_height[0]_pin[50] 
+ svdd sgnd grid[1][1]_clb[0]_mode[clb]
.eom
