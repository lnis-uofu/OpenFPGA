// Benchmark "TOP" written by ABC on Mon Feb  4 17:31:57 2019

module ex5p ( 
    i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_,
    o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_,
    o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_,
    o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_,
    o_31_, o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_, o_40_,
    o_41_, o_42_, o_43_, o_44_, o_45_, o_46_, o_47_, o_48_, o_49_, o_50_,
    o_51_, o_52_, o_53_, o_54_, o_55_, o_56_, o_57_, o_58_, o_59_, o_60_,
    o_61_, o_62_  );
  input  i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_;
  output o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_,
    o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_,
    o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_,
    o_31_, o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_, o_40_,
    o_41_, o_42_, o_43_, o_44_, o_45_, o_46_, o_47_, o_48_, o_49_, o_50_,
    o_51_, o_52_, o_53_, o_54_, o_55_, o_56_, o_57_, o_58_, o_59_, o_60_,
    o_61_, o_62_;
  wire n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
    n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
    n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
    n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
    n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
    n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
    n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
    n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
    n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
    n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
    n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
    n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
    n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
    n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
    n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
    n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
    n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
    n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
    n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
    n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
    n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
    n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
    n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
    n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
    n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
    n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
    n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
    n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
    n589, n590, n591, n592, n593, n594, n595, n596, n597;
  assign o_0_ = ~n365;
  assign o_1_ = ~n361;
  assign o_2_ = ~n403;
  assign o_3_ = ~n370;
  assign o_4_ = ~n450;
  assign o_5_ = ~n357;
  assign o_6_ = ~n136;
  assign o_7_ = ~n180;
  assign o_8_ = ~n452;
  assign o_9_ = ~n491;
  assign o_10_ = ~n139;
  assign o_11_ = ~n179;
  assign o_12_ = ~n385;
  assign o_13_ = ~n471;
  assign o_14_ = ~n507;
  assign o_15_ = ~n138;
  assign o_16_ = ~n407;
  assign o_17_ = ~n354;
  assign o_18_ = ~n421;
  assign o_19_ = ~n420;
  assign o_20_ = ~n142;
  assign o_21_ = ~n145;
  assign o_22_ = ~n148;
  assign o_23_ = ~n352;
  assign o_24_ = ~n504;
  assign o_25_ = ~n200;
  assign o_26_ = ~n151;
  assign o_27_ = ~n260;
  assign o_28_ = ~n556;
  assign o_29_ = ~n506;
  assign o_30_ = ~n150;
  assign o_31_ = ~n347;
  assign o_32_ = ~n344;
  assign o_33_ = ~n340;
  assign o_34_ = ~n336;
  assign o_35_ = ~n332;
  assign o_36_ = ~n328;
  assign o_37_ = ~n321;
  assign o_38_ = ~n314;
  assign o_39_ = ~n308;
  assign o_40_ = ~n303;
  assign o_41_ = ~n296;
  assign o_42_ = ~n291;
  assign o_43_ = ~n284;
  assign o_44_ = ~n276;
  assign o_45_ = ~n274;
  assign o_46_ = ~n268;
  assign o_47_ = ~n264;
  assign o_48_ = ~n259;
  assign o_49_ = ~n257;
  assign o_50_ = ~n252;
  assign o_51_ = ~n245;
  assign o_52_ = ~n238;
  assign o_53_ = ~n232;
  assign o_54_ = ~n226;
  assign o_55_ = ~n220;
  assign o_56_ = ~n214;
  assign o_57_ = ~n205;
  assign o_58_ = ~n197;
  assign o_59_ = ~n189;
  assign o_60_ = ~n182;
  assign o_61_ = ~n173;
  assign o_62_ = ~n164;
  assign n134 = n155 | n439;
  assign n135 = n155 | n441;
  assign n136 = n134 & n135;
  assign n137 = n436 | n339;
  assign n138 = n445 | n339;
  assign n139 = n137 & n138;
  assign n140 = n462 | n152;
  assign n141 = n463 | n152;
  assign n142 = n140 & n141;
  assign n143 = n439 | n152;
  assign n144 = n441 | n152;
  assign n145 = n143 & n144;
  assign n146 = n434 | n152;
  assign n147 = n446 | n152;
  assign n148 = n146 & n147;
  assign n149 = n434 | n373;
  assign n150 = n434 | n369;
  assign n151 = n149 & n150;
  assign n152 = i_2_ | ~i_0_ | i_1_;
  assign n153 = n152 | ~n381;
  assign n154 = ~i_3_ | ~i_4_ | ~i_5_;
  assign n155 = i_0_ | i_1_ | ~i_2_;
  assign n156 = n154 | n155;
  assign n157 = i_0_ | i_1_ | i_2_;
  assign n158 = n157 | ~n366;
  assign n159 = n373 & n338;
  assign n160 = n514 & n505 & n363;
  assign n161 = n515 & n339 & n269 & n195 & n496;
  assign n162 = n179 & n458 & n408 & n461 & n374;
  assign n163 = n150 & n516 & n517 & n176 & n454;
  assign n164 = n159 & n160 & n161 & n162 & n163;
  assign n165 = n398 & n533 & n535;
  assign n166 = n523 & n524;
  assign n167 = n412 & n503;
  assign n168 = n504 & n363;
  assign n169 = n450 & n556;
  assign n170 = n372 & n555 & n180;
  assign n171 = n254 & n243 & n400;
  assign n172 = n518 & n192 & n554;
  assign n173 = n165 & n166 & n167 & n168 & n169 & n170 & n171 & n172;
  assign n174 = n208 & n309 & n563 & n421 & n254 & n518;
  assign n175 = n410 & n560 & n192 & n165 & n457 & n461 & n150 & n516;
  assign n176 = n452 & n451;
  assign n177 = n362 & n552 & n454;
  assign n178 = n369 | n462;
  assign n179 = n436 | n409;
  assign n180 = n436 | n270;
  assign n181 = n369 | n463;
  assign n182 = n174 & n175 & n176 & n177 & n178 & n179 & n180 & n181;
  assign n183 = n411 & (n157 | ~n382) & n412;
  assign n184 = n548 & n298;
  assign n185 = n418 & (n239 | n409);
  assign n186 = n569 & n570 & n310 & n345 & n169 & n334 & n255 & n163;
  assign n187 = n265 & n573 & n170 & n203;
  assign n188 = n594 & n493 & n487 & n483 & n408 & n397 & ~n383 & n387;
  assign n189 = n183 & n184 & n185 & n186 & n187 & n188;
  assign n190 = n576 & n575 & n532 & n451 & n414 & n140 & n297 & ~n367;
  assign n191 = n493 & ~n383 & n492;
  assign n192 = n405 & n550 & n404 & n145 & n551 & n549;
  assign n193 = n563 & n272;
  assign n194 = n421 & n485 & n487;
  assign n195 = n478 & n481 & n475 & n477;
  assign n196 = n351 & n158 & (n154 | n157);
  assign n197 = n190 & n191 & n192 & n193 & n194 & n195 & n138 & n196;
  assign n198 = n470 & n468;
  assign n199 = n150 & n536;
  assign n200 = n270 | n443;
  assign n201 = n261 & n471 & n394;
  assign n202 = n228 & n414 & (n339 | ~n382);
  assign n203 = n179 & n572;
  assign n204 = n221 & n215 & n422 & n185 & n423 & n300;
  assign n205 = n198 & n199 & n200 & n201 & n166 & n202 & n203 & n204;
  assign n206 = n578 & n579 & n554 & n169;
  assign n207 = n310 & n577;
  assign n208 = n496 & n562;
  assign n209 = n580 & ~n395 & n491;
  assign n210 = n149 & n378 & n370 & n419 & n306;
  assign n211 = n501 & n563;
  assign n212 = n180 & n518;
  assign n213 = n228 & n171 & n467 & n196 & n594 & n376 & n534 & n471;
  assign n214 = n206 & n207 & n208 & n209 & n210 & n211 & n212 & n213;
  assign n215 = n563 & n183;
  assign n216 = n537 & ~n367 & n451;
  assign n217 = n534 & n275 & n139 & n142;
  assign n218 = n570 & n571 & n184 & n581 & n337 & n582;
  assign n219 = n156 & n171 & n427 & n200;
  assign n220 = n215 & n216 & n180 & n166 & n217 & n218 & n219;
  assign n221 = n396 & n180 & n159;
  assign n222 = n474 & n247;
  assign n223 = n519 & n348 & n494;
  assign n224 = n472 & n470;
  assign n225 = n572 & n575 & n478 & n538 & n158 & n458 & n534 & n468;
  assign n226 = n209 & n219 & n193 & n221 & n222 & n223 & n224 & n225;
  assign n227 = n449 & n452;
  assign n228 = n525 & n526;
  assign n229 = n146 & n527 & n528 & n529 & n530;
  assign n230 = n391 & n392 & (n393 | n339);
  assign n231 = n476 & n583 & n537 & n137 & n141 & n534;
  assign n232 = n174 & n218 & n227 & n228 & n229 & n230 & n231;
  assign n233 = n351 & n215;
  assign n234 = n254 & n494 & n559 & n509 & n262 & n292 & n426;
  assign n235 = n387 & n491;
  assign n236 = n384 & n385 & (n373 | n386);
  assign n237 = n510 & n548;
  assign n238 = n233 & n234 & n224 & n235 & n236 & n186 & n162 & n237;
  assign n239 = ~n381 & ~n382;
  assign n240 = n155 | n239;
  assign n241 = n255 & n240 & n389 & n387 & n584 & n491;
  assign n242 = n488 & n489;
  assign n243 = n421 & n482;
  assign n244 = n254 & n494 & n453;
  assign n245 = n175 & n212 & n227 & n233 & n241 & n242 & n243 & n244;
  assign n246 = n560 & n203;
  assign n247 = n408 & ((~n381 & ~n382) | n409);
  assign n248 = n200 & n483 & n486;
  assign n249 = n540 & n539;
  assign n250 = n524 & n192 & n412 & n501 & n168 & n288 & n293;
  assign n251 = n535 & n543 & n546 & n477 & n380 & n533;
  assign n252 = n246 & n247 & n248 & n249 & n250 & n251;
  assign n253 = n288 & n248 & n342 & n586 & n266;
  assign n254 = n155 | n446;
  assign n255 = n155 | n443;
  assign n256 = n350 & n158 & n351 & n520;
  assign n257 = n193 & n235 & n253 & n254 & n255 & n256;
  assign n258 = n254 & n241 & n135 & n134;
  assign n259 = n258 & n253 & n242 & n160;
  assign n260 = n443 | n339;
  assign n261 = n434 | n339;
  assign n262 = n429 & n281 & n248;
  assign n263 = n417 & n224 & (n393 | n270);
  assign n264 = n260 & n190 & n139 & n261 & n262 & n250 & n263;
  assign n265 = n421 & n156 & n468 & n200;
  assign n266 = n210 & n585 & n345 & n207;
  assign n267 = n196 & n496 & n160 & n396 & n180 & n515;
  assign n268 = n265 & n191 & n206 & n263 & n266 & n267;
  assign n269 = n493 & n492 & n194 & n196 & ~n383;
  assign n270 = i_2_ | i_0_ | ~i_1_;
  assign n271 = n260 & n261;
  assign n272 = n500 & n330 & n420 & n411 & n497 & n498;
  assign n273 = n577 & n206 & n210;
  assign n274 = n269 & n168 & n270 & n271 & n272 & n217 & n273;
  assign n275 = n530 & n568 & n146 & n529;
  assign n276 = n211 & n273 & n161 & n275;
  assign n277 = n567 & n530 & n482 & ~n415 & n137 & n228 & ~n395;
  assign n278 = n196 & n330 & n451 & n431 & n254 & n491 & n588 & n589;
  assign n279 = n484 & n363 & n486 & n502;
  assign n280 = n180 & (n270 | n355);
  assign n281 = n476 & n583 & n468 & n396;
  assign n282 = n298 & n417 & n222;
  assign n283 = n511 & n405 & n499 & n508 & n374 & n377 & n179 & n595;
  assign n284 = n277 & n278 & n249 & n279 & n280 & n281 & n282 & n283;
  assign n285 = n477 & n394 & n471 & n378;
  assign n286 = n413 & n423 & n590 & n138 & n144 & n228;
  assign n287 = n179 & n553;
  assign n288 = n422 & n243;
  assign n289 = n419 & n420 & n579;
  assign n290 = n549 & n406 & n410 & n563 & n569 & n411 & n380 & n596;
  assign n291 = n285 & n286 & n248 & n278 & n287 & n288 & n289 & n290;
  assign n292 = n288 & n404 & (n152 | ~n366);
  assign n293 = n326 & n426 & n258;
  assign n294 = n585 & n586 & n345 & n248;
  assign n295 = n547 & n405 & n560 & n542 & n543 & n546;
  assign n296 = n292 & n293 & n294 & n193 & n207 & n223 & n295;
  assign n297 = n458 & n246 & n247;
  assign n298 = n402 & n547;
  assign n299 = n356 & n550 & n564;
  assign n300 = n254 & n400 & n543;
  assign n301 = n405 & n318 & n473 & n536 & n476 & n469 & n474 & n409;
  assign n302 = n482 & n411 & n153 & n339 & n380 & n330 & n523;
  assign n303 = n275 & n297 & n298 & n299 & n300 & n279 & n301 & n302;
  assign n304 = n573 & n185 & n581 & n587 & n315 & n167 & n203 & n591;
  assign n305 = n153 & n531;
  assign n306 = n356 & n564 & n184;
  assign n307 = n470 & n142 & n145 & n194 & n261 & ~n382;
  assign n308 = n277 & n285 & n304 & n305 & n306 & n258 & n307;
  assign n309 = n196 & n492 & n561;
  assign n310 = n142 & n275 & ~n415;
  assign n311 = n149 & n298 & n419;
  assign n312 = n147 & n370 & n508;
  assign n313 = n327 & n503 & n363;
  assign n314 = n309 & n310 & n206 & n294 & n311 & n312 & n208 & n313;
  assign n315 = n575 & n576 & n457 & n454;
  assign n316 = n448 & n513 & n459;
  assign n317 = n447 & n512 & n136 & n145 & n526 & n495 & n460;
  assign n318 = n525 & n478 & n481;
  assign n319 = n405 & n562 & n578 & n230 & n532 & n371;
  assign n320 = n541 & n556 & n147 & n449 & n510 & n551 & n565 & n597;
  assign n321 = n315 & n316 & n317 & n211 & n234 & n318 & n319 & n320;
  assign n322 = n477 & n550 & n342 & n318 & n311 & n471 & n470 & n592;
  assign n323 = n146 & n590;
  assign n324 = n561 & n548 & n531 & n491 & ~n382 & n387;
  assign n325 = n356 & n507;
  assign n326 = n242 & n256;
  assign n327 = n482 & n254;
  assign n328 = n322 & n323 & n193 & n324 & n325 & n326 & n327 & n194;
  assign n329 = n325 & n353 & (n152 | ~n381);
  assign n330 = n515 & n495;
  assign n331 = n531 & n486 & n485;
  assign n332 = n243 & n293 & n322 & n323 & n329 & n330 & n211 & n331;
  assign n333 = n143 & (n152 | ~n382);
  assign n334 = n416 & (n270 | ~n366) & n417;
  assign n335 = n518 & n398 & n243 & n180 & n254 & n508;
  assign n336 = n286 & n304 & n324 & n298 & n333 & n334 & n335;
  assign n337 = n572 & n578 & n287;
  assign n338 = n152 & n511 & n312 & n402 & n512 & n513;
  assign n339 = ~i_2_ | i_0_ | ~i_1_;
  assign n340 = n216 & n301 & n211 & n337 & n338 & n208 & n339 & n269;
  assign n341 = n550 & n311 & n329;
  assign n342 = n206 & n223;
  assign n343 = n180 & n482;
  assign n344 = n279 & n341 & n258 & n342 & n326 & n272 & n165 & n343;
  assign n345 = n202 & n413 & n567;
  assign n346 = n523 & n505 & n229 & n305 & n330 & n363 & ~n415;
  assign n347 = n345 & n206 & n171 & n334 & n224 & n262 & n341 & n346;
  assign n348 = n157 | n370;
  assign n349 = n519 & n520;
  assign n350 = n154 | n157;
  assign n351 = n445 | n157;
  assign n352 = n348 & n349 & n350 & n351;
  assign n353 = n152 | ~n366;
  assign n354 = n153 & n353;
  assign n355 = n435 | n442;
  assign n356 = n442 | n444;
  assign n357 = n355 & n356;
  assign n358 = n157 | n462;
  assign n359 = n488 & n515 & n178 & n552 & n316 & n396 & n486 & n593;
  assign n360 = (~n366 & ~n381) | n438;
  assign n361 = n143 & n358 & n134 & n140 & n359 & n360;
  assign n362 = n409 | n463;
  assign n363 = n358 & n506;
  assign n364 = n468 & n483 & n489 & n142 & n509 & n465;
  assign n365 = n181 & n362 & n363 & n317 & n359 & n364;
  assign n366 = i_3_ & i_4_ & ~i_5_;
  assign n367 = ~n369 & (~n154 | n366);
  assign n368 = n369 | (n356 & n378);
  assign n369 = ~i_0_ | ~i_1_ | ~i_2_;
  assign n370 = n438 | n444;
  assign n371 = n368 & (n369 | n370);
  assign n372 = n445 | n373;
  assign n373 = ~i_2_ | ~i_0_ | i_1_;
  assign n374 = n372 & ((n154 & ~n366) | n373);
  assign n375 = n339 | n239;
  assign n376 = n464 & n465;
  assign n377 = n376 & (n270 | n154);
  assign n378 = n440 | n444;
  assign n379 = n270 | (n356 & n378);
  assign n380 = n180 & (n270 | ~n381);
  assign n381 = ~i_5_ & ~i_3_ & i_4_;
  assign n382 = i_5_ & ~i_3_ & i_4_;
  assign n383 = ~n155 & (n381 | n382);
  assign n384 = n373 | n355;
  assign n385 = n436 | n373;
  assign n386 = n435 | n440;
  assign n387 = n155 | n436;
  assign n388 = n387 & (n155 | ~n381);
  assign n389 = n155 | (n355 & n386);
  assign n390 = ~n157 & (~n154 | n366);
  assign n391 = n378 | n339;
  assign n392 = n140 & n138 & n566;
  assign n393 = n154 & ~n366;
  assign n394 = n260 & n376 & (n393 | n270);
  assign n395 = ~n339 & (n381 | n382);
  assign n396 = n270 | n439;
  assign n397 = n396 & (n270 | ~n382);
  assign n398 = n198 & n397 & (n270 | ~n381);
  assign n399 = n155 | ~n382;
  assign n400 = n136 & (n239 | n155);
  assign n401 = n369 | (n355 & n386);
  assign n402 = n443 | n373;
  assign n403 = n435 | n438;
  assign n404 = n149 & n402 & (n373 | n403);
  assign n405 = n236 & (n239 | n373);
  assign n406 = n372 & (n393 | n373);
  assign n407 = n409 | n445;
  assign n408 = n459 & n460;
  assign n409 = ~i_0_ | ~i_1_ | i_2_;
  assign n410 = n407 & n408 & (n393 | n409);
  assign n411 = n436 | n157;
  assign n412 = n157 | ~n381;
  assign n413 = n137 & (n339 | ~n381);
  assign n414 = n391 & n565 & n534;
  assign n415 = ~n339 & (~n154 | n366);
  assign n416 = n271 & n377;
  assign n417 = n471 & n379;
  assign n418 = n407 & n455 & n456;
  assign n419 = n385 & (n373 | ~n381);
  assign n420 = n412 & (n157 | ~n382);
  assign n421 = n155 | ~n366;
  assign n422 = n421 & (n155 | n154);
  assign n423 = n339 | (n239 & n393);
  assign n424 = n373 | n393;
  assign n425 = n155 | (n356 & n378);
  assign n426 = n425 & (n155 | n370);
  assign n427 = n434 | n270;
  assign n428 = n270 | (n386 & n403);
  assign n429 = n280 & n427 & n428;
  assign n430 = n409 | (n434 & n443);
  assign n431 = n386 & n355 & n430;
  assign n432 = i_3_ | i_4_ | i_5_;
  assign n433 = ~i_6_ | ~i_7_;
  assign n434 = n432 | n433;
  assign n435 = i_3_ | i_4_ | ~i_5_;
  assign n436 = n433 | n435;
  assign n437 = i_5_ | ~i_3_ | i_4_;
  assign n438 = i_6_ | i_7_;
  assign n439 = n437 | n438;
  assign n440 = i_6_ | ~i_7_;
  assign n441 = n437 | n440;
  assign n442 = ~i_6_ | i_7_;
  assign n443 = n432 | n442;
  assign n444 = ~i_5_ | ~i_3_ | i_4_;
  assign n445 = n433 | n444;
  assign n446 = n433 | n437;
  assign n447 = n369 | n441;
  assign n448 = n369 | n439;
  assign n449 = n369 | n446;
  assign n450 = n437 | n442;
  assign n451 = n447 & n448 & n449 & n450;
  assign n452 = n436 | n369;
  assign n453 = n369 | n445;
  assign n454 = ~n367 & n453;
  assign n455 = n409 | n356;
  assign n456 = n409 | n378;
  assign n457 = n409 | n446;
  assign n458 = n457 & n418;
  assign n459 = n439 | n409;
  assign n460 = n441 | n409;
  assign n461 = n403 & n431;
  assign n462 = n432 | n438;
  assign n463 = n432 | n440;
  assign n464 = n339 | n462;
  assign n465 = n339 | n463;
  assign n466 = n403 | n339;
  assign n467 = n466 & n271;
  assign n468 = n270 | n441;
  assign n469 = n468 & n396;
  assign n470 = n270 | n446;
  assign n471 = n270 | n445;
  assign n472 = n270 | n370;
  assign n473 = n470 & n379 & n471 & n472;
  assign n474 = n270 | ~n366;
  assign n475 = n474 & n473;
  assign n476 = n270 | ~n382;
  assign n477 = n476 & n469;
  assign n478 = n377 & n467;
  assign n479 = n386 | n339;
  assign n480 = n355 | n339;
  assign n481 = n479 & n375 & n137 & n480;
  assign n482 = n155 | n445;
  assign n483 = n270 | n463;
  assign n484 = n427 & n200 & n483;
  assign n485 = n484 & n380;
  assign n486 = n270 | n462;
  assign n487 = n486 & n156;
  assign n488 = n155 | n462;
  assign n489 = n155 | n463;
  assign n490 = n255 & n242;
  assign n491 = n434 | n155;
  assign n492 = n387 & n491 & n490;
  assign n493 = n136 & n327;
  assign n494 = n446 | n157;
  assign n495 = n441 | n157;
  assign n496 = n494 & n495;
  assign n497 = n355 | n157;
  assign n498 = n386 | n157;
  assign n499 = n411 & n497 & n498;
  assign n500 = n403 | n157;
  assign n501 = n500 & n499;
  assign n502 = n434 | n157;
  assign n503 = n502 & n501;
  assign n504 = n443 | n157;
  assign n505 = n412 & n504 & n503;
  assign n506 = n157 | n463;
  assign n507 = n445 | n152;
  assign n508 = n378 & n325;
  assign n509 = n441 | n373;
  assign n510 = n439 | n373;
  assign n511 = n509 & n510;
  assign n512 = n373 | n463;
  assign n513 = n373 | n462;
  assign n514 = n157 | ~n382;
  assign n515 = n439 | n157;
  assign n516 = n369 | n443;
  assign n517 = n393 | n409;
  assign n518 = n486 & n156 & n484;
  assign n519 = n378 | n157;
  assign n520 = n356 | n157;
  assign n521 = n584 & n491 & n255;
  assign n522 = n521 & n489 & n488 & n349 & n351 & n388 & n389 & ~n390;
  assign n523 = n494 & n522;
  assign n524 = n514 & n330;
  assign n525 = n439 | n339;
  assign n526 = n441 | n339;
  assign n527 = n355 | n152;
  assign n528 = n386 | n152;
  assign n529 = n403 | n152;
  assign n530 = n443 | n152;
  assign n531 = n436 | n152;
  assign n532 = n141 & n229 & n305;
  assign n533 = n137 & n201 & ~n395;
  assign n534 = n446 | n339;
  assign n535 = n230 & n532 & n534 & n228;
  assign n536 = n516 & n181 & n178;
  assign n537 = n239 | n369;
  assign n538 = n537 & n451 & n454 & n401 & n371;
  assign n539 = n407 & n455;
  assign n540 = ~n366 | n409;
  assign n541 = n409 | n370;
  assign n542 = n540 & n408 & n539 & n456 & n541 & n457;
  assign n543 = n452 & n538;
  assign n544 = n369 | n403;
  assign n545 = n154 | n409;
  assign n546 = n544 & n545 & n199;
  assign n547 = n513 & n512;
  assign n548 = n154 | n152;
  assign n549 = n325 & n547 & n353 & n548;
  assign n550 = n147 & n378 & n370;
  assign n551 = n152 | ~n382;
  assign n552 = n409 | n462;
  assign n553 = n239 | n409;
  assign n554 = n543 & n546 & n461 & n542 & n552 & n553 & n179 & n362;
  assign n555 = n373 | ~n382;
  assign n556 = n446 | n373;
  assign n557 = n356 | n373;
  assign n558 = n378 | n373;
  assign n559 = n373 | n370;
  assign n560 = n511 & n169 & n406 & n557 & n558 & n559;
  assign n561 = n136 & ~n383;
  assign n562 = n515 & n514 & n412;
  assign n563 = n502 & n168;
  assign n564 = n507 & n353;
  assign n565 = n339 | n370;
  assign n566 = n356 | n339;
  assign n567 = n138 & n566;
  assign n568 = n531 & n527 & n528;
  assign n569 = n153 & n333;
  assign n570 = n144 & n299;
  assign n571 = n149 & n419;
  assign n572 = n362 & n552 & n461;
  assign n573 = n326 & n571 & n524 & n168;
  assign n574 = n452 & n537 & n401;
  assign n575 = n517 & n199;
  assign n576 = n544 & n574;
  assign n577 = n153 & n333 & n144 & n147;
  assign n578 = n558 & n424 & n372 & n557;
  assign n579 = n509 & n510 & n555;
  assign n580 = n350 & n490;
  assign n581 = n169 & n579;
  assign n582 = n473 & n536 & n569 & n150 & n458 & n271;
  assign n583 = n270 | ~n381;
  assign n584 = n155 | n403;
  assign n585 = n466 & n416 & n480 & n479;
  assign n586 = n429 & n281 & n263;
  assign n587 = n534 & n494;
  assign n588 = n457 & n261 & n470;
  assign n589 = n580 & n587 & n568 & n574 & n536 & n177 & n388 & n400;
  assign n590 = n142 & n530;
  assign n591 = n451 & n408 & n374;
  assign n592 = n145 & n339 & n474;
  assign n593 = n510 & n525 & n464;
  assign n594 = n239 | n270;
  assign n595 = n545 & n260;
  assign n596 = n151 & n402 & n427;
  assign n597 = n418 & n475 & n522 & n534 & n348 & n399;
endmodule


