//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog netlist for pre-configured FPGA fabric by design: and2
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Wed Jun 10 20:32:40 2020
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

module and2_top_formal_verification (
input [0:0] a_fm,
input [0:0] b_fm,
output [0:0] out_c_fm);

// ----- Local wires for FPGA fabric -----
wire [0:0] pReset;
wire [0:0] prog_clk;
wire [0:0] set;
wire [0:0] reset;
wire [0:0] clk;
wire [0:63] gfpga_pad_iopad_pad;
wire [0:0] enable;
wire [0:15] address;
wire [0:0] data_in;

// ----- FPGA top-level module to be capsulated -----
	fpga_top U0_formal_verification (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.set(set[0]),
		.reset(reset[0]),
		.clk(clk[0]),
		.gfpga_pad_iopad_pad(gfpga_pad_iopad_pad[0:63]),
		.enable(enable[0]),
		.address(address[0:15]),
		.data_in(data_in[0]));

// ----- Begin Connect Global ports of FPGA top module -----
	assign pReset[0] = {1{1'b0}};
	assign prog_clk[0] = {1{1'b0}};
	assign set[0] = {1{1'b0}};
	assign reset[0] = {1{1'b0}};
// ----- End Connect Global ports of FPGA top module -----

// ----- Link BLIF Benchmark I/Os to FPGA I/Os -----
// ----- Blif Benchmark input a is mapped to FPGA IOPAD gfpga_pad_iopad_pad[17] -----
	assign gfpga_pad_iopad_pad[17] = a_fm[0];
// ----- Blif Benchmark input b is mapped to FPGA IOPAD gfpga_pad_iopad_pad[40] -----
	assign gfpga_pad_iopad_pad[40] = b_fm[0];
// ----- Blif Benchmark output out_c is mapped to FPGA IOPAD gfpga_pad_iopad_pad[46] -----
	assign out_c_fm[0] = gfpga_pad_iopad_pad[46];

// ----- Wire unused FPGA I/Os to constants -----
	assign gfpga_pad_iopad_pad[0] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[1] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[2] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[3] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[4] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[5] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[6] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[7] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[8] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[9] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[10] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[11] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[12] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[13] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[14] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[15] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[16] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[18] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[19] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[20] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[21] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[22] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[23] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[24] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[25] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[26] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[27] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[28] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[29] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[30] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[31] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[32] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[33] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[34] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[35] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[36] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[37] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[38] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[39] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[41] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[42] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[43] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[44] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[45] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[47] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[48] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[49] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[50] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[51] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[52] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[53] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[54] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[55] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[56] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[57] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[58] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[59] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[60] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[61] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[62] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[63] = {1{1'b0}};

// ----- Begin load bitstream to configuration memories -----
`ifdef ICARUS_SIMULATOR
// ----- Begin assign bitstream to configuration memories -----
	assign U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15] = 16'b1010101000000000;
	assign U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b010;
	assign U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:7] = 8'b00100100;
	assign U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:7] = 8'b10001000;
	assign U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15] = {16{1'b0}};
	assign U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2] = 3'b001;
	assign U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:7] = 8'b00100001;
	assign U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b0}};
	assign U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0] = {1{1'b1}};
	assign U0_formal_verification.sb_0__0_.mem_top_track_0.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__0_.mem_top_track_2.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__0_.mem_top_track_4.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__0_.mem_top_track_6.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__0_.mem_top_track_8.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__0_.mem_top_track_10.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__0_.mem_top_track_12.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__0_.mem_top_track_14.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__0_.mem_top_track_16.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_0.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_2.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_4.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_6.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_8.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_10.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_12.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_14.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_16.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__1_.mem_top_track_0.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_0__1_.mem_top_track_8.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_0__1_.mem_top_track_16.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_0__1_.mem_right_track_2.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_4.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_6.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_8.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_10.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_12.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_14.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_0__1_.mem_bottom_track_9.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_0__1_.mem_bottom_track_17.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_0__2_.mem_right_track_0.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_2.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_4.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_6.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_8.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_10.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_12.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_14.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_16.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__2_.mem_bottom_track_3.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__2_.mem_bottom_track_5.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__2_.mem_bottom_track_7.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__2_.mem_bottom_track_9.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__2_.mem_bottom_track_11.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__2_.mem_bottom_track_13.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__2_.mem_bottom_track_15.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_0__2_.mem_bottom_track_17.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_0.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_1__0_.mem_top_track_2.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_8.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_14.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_16.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_1__0_.mem_right_track_0.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_1__0_.mem_right_track_8.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_1__0_.mem_right_track_16.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_1__0_.mem_left_track_1.mem_out[0:5] = 6'b010100;
	assign U0_formal_verification.sb_1__0_.mem_left_track_9.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_1__0_.mem_left_track_17.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_1__1_.mem_top_track_0.mem_out[0:7] = 8'b10001000;
	assign U0_formal_verification.sb_1__1_.mem_top_track_8.mem_out[0:7] = 8'b10001000;
	assign U0_formal_verification.sb_1__1_.mem_top_track_16.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_1__1_.mem_right_track_0.mem_out[0:7] = 8'b10001000;
	assign U0_formal_verification.sb_1__1_.mem_right_track_8.mem_out[0:7] = 8'b10001000;
	assign U0_formal_verification.sb_1__1_.mem_right_track_16.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_out[0:7] = 8'b00101000;
	assign U0_formal_verification.sb_1__1_.mem_bottom_track_9.mem_out[0:7] = 8'b10001000;
	assign U0_formal_verification.sb_1__1_.mem_bottom_track_17.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_1__1_.mem_left_track_1.mem_out[0:7] = 8'b10001000;
	assign U0_formal_verification.sb_1__1_.mem_left_track_9.mem_out[0:7] = 8'b10001000;
	assign U0_formal_verification.sb_1__1_.mem_left_track_17.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_1__2_.mem_right_track_0.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_1__2_.mem_right_track_8.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_1__2_.mem_right_track_16.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_3.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_5.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_7.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_9.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_11.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_13.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_15.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_17.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_1__2_.mem_left_track_1.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_1__2_.mem_left_track_9.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_1__2_.mem_left_track_17.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_2__0_.mem_top_track_0.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_2.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_4.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_6.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_8.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_10.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_12.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_14.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_16.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_1.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_3.mem_out[0:1] = 2'b01;
	assign U0_formal_verification.sb_2__0_.mem_left_track_5.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_7.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_9.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_11.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_13.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_15.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_17.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__1_.mem_top_track_0.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_2__1_.mem_top_track_8.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_2__1_.mem_top_track_16.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_2__1_.mem_bottom_track_9.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_2__1_.mem_bottom_track_17.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.sb_2__1_.mem_left_track_1.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_3.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_5.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_7.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_9.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_11.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_13.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_15.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_17.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_3.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_5.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_7.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_9.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_11.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_13.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_15.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_17.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__2_.mem_left_track_1.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__2_.mem_left_track_3.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__2_.mem_left_track_5.mem_out[0:1] = 2'b01;
	assign U0_formal_verification.sb_2__2_.mem_left_track_7.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__2_.mem_left_track_9.mem_out[0:1] = 2'b01;
	assign U0_formal_verification.sb_2__2_.mem_left_track_11.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__2_.mem_left_track_13.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__2_.mem_left_track_15.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.sb_2__2_.mem_left_track_17.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_1__0_.mem_top_ipin_1.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_1__0_.mem_top_ipin_2.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_1__0_.mem_top_ipin_3.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_1__0_.mem_top_ipin_4.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_1__0_.mem_top_ipin_5.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_1__0_.mem_top_ipin_6.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_1__0_.mem_top_ipin_7.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_1__1_.mem_top_ipin_0.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_1__1_.mem_top_ipin_1.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.cbx_1__1_.mem_top_ipin_2.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_1__2_.mem_bottom_ipin_3.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_1__2_.mem_bottom_ipin_4.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_1__2_.mem_bottom_ipin_5.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_1__2_.mem_bottom_ipin_6.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_1__2_.mem_bottom_ipin_7.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_1__2_.mem_top_ipin_0.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_1__2_.mem_top_ipin_1.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.cbx_1__2_.mem_top_ipin_2.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.mem_out[0:1] = 2'b01;
	assign U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_2__0_.mem_top_ipin_1.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_2__0_.mem_top_ipin_2.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_2__0_.mem_top_ipin_3.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_2__0_.mem_top_ipin_4.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_2__0_.mem_top_ipin_5.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_2__0_.mem_top_ipin_6.mem_out[0:5] = 6'b001100;
	assign U0_formal_verification.cbx_2__0_.mem_top_ipin_7.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_2__1_.mem_top_ipin_0.mem_out[0:5] = 6'b100010;
	assign U0_formal_verification.cbx_2__1_.mem_top_ipin_1.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.cbx_2__1_.mem_top_ipin_2.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_2__2_.mem_bottom_ipin_3.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_2__2_.mem_bottom_ipin_4.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_2__2_.mem_bottom_ipin_5.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_2__2_.mem_bottom_ipin_6.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_2__2_.mem_bottom_ipin_7.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_2__2_.mem_top_ipin_0.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cbx_2__2_.mem_top_ipin_1.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.cbx_2__2_.mem_top_ipin_2.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.cby_0__1_.mem_left_ipin_0.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_0__1_.mem_left_ipin_1.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_0__1_.mem_right_ipin_1.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_0__1_.mem_right_ipin_2.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_0__1_.mem_right_ipin_3.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_0__1_.mem_right_ipin_4.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_0__1_.mem_right_ipin_5.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_0__1_.mem_right_ipin_6.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_0__1_.mem_right_ipin_7.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_0__2_.mem_left_ipin_0.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_0__2_.mem_left_ipin_1.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_0__2_.mem_right_ipin_1.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_0__2_.mem_right_ipin_2.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_0__2_.mem_right_ipin_3.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_0__2_.mem_right_ipin_4.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_0__2_.mem_right_ipin_5.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_0__2_.mem_right_ipin_6.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_0__2_.mem_right_ipin_7.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_1__1_.mem_left_ipin_0.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_1__1_.mem_left_ipin_1.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.cby_1__2_.mem_left_ipin_0.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_1__2_.mem_left_ipin_1.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.cby_2__1_.mem_left_ipin_0.mem_out[0:5] = 6'b010100;
	assign U0_formal_verification.cby_2__1_.mem_left_ipin_1.mem_out[0:5] = 6'b010100;
	assign U0_formal_verification.cby_2__1_.mem_left_ipin_2.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_2__1_.mem_left_ipin_3.mem_out[0:5] = 6'b010100;
	assign U0_formal_verification.cby_2__1_.mem_left_ipin_4.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_2__1_.mem_left_ipin_5.mem_out[0:5] = 6'b010100;
	assign U0_formal_verification.cby_2__1_.mem_left_ipin_6.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_2__1_.mem_left_ipin_7.mem_out[0:5] = 6'b010100;
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_0.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_1.mem_out[0:1] = 2'b01;
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_2.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.cby_2__2_.mem_left_ipin_0.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_2__2_.mem_left_ipin_1.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_2__2_.mem_left_ipin_2.mem_out[0:5] = 6'b010100;
	assign U0_formal_verification.cby_2__2_.mem_left_ipin_3.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_2__2_.mem_left_ipin_4.mem_out[0:5] = 6'b010100;
	assign U0_formal_verification.cby_2__2_.mem_left_ipin_5.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_2__2_.mem_left_ipin_6.mem_out[0:5] = 6'b010100;
	assign U0_formal_verification.cby_2__2_.mem_left_ipin_7.mem_out[0:5] = 6'b100100;
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_0.mem_out[0:5] = 6'b010100;
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_1.mem_out[0:1] = {2{1'b1}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_2.mem_out[0:1] = 2'b01;
initial begin
	force U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15] = 16'b0101010111111111;
	force U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:7] = 8'b11011011;
	force U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:7] = 8'b11011110;
	force U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b1}};
	force U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0] = {1{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_0.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_2.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_4.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_6.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_10.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_12.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_14.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_16.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_0.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_2.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_4.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_6.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_8.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_10.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_12.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_14.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_16.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_0__1_.mem_top_track_8.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_0__1_.mem_top_track_16.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_0__1_.mem_right_track_2.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_4.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_6.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_8.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_10.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_12.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_14.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_9.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_17.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_0__2_.mem_right_track_0.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_2.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_4.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_6.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_8.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_10.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_12.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_14.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_16.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__0_.mem_top_track_2.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_14.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_16.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__0_.mem_right_track_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__0_.mem_right_track_8.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__0_.mem_right_track_16.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__0_.mem_left_track_1.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.sb_1__0_.mem_left_track_9.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__0_.mem_left_track_17.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__1_.mem_top_track_0.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.sb_1__1_.mem_top_track_8.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.sb_1__1_.mem_top_track_16.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__1_.mem_right_track_0.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.sb_1__1_.mem_right_track_8.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.sb_1__1_.mem_right_track_16.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_outb[0:7] = 8'b11010111;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_9.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_17.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__1_.mem_left_track_1.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.sb_1__1_.mem_left_track_9.mem_outb[0:7] = 8'b01110111;
	force U0_formal_verification.sb_1__1_.mem_left_track_17.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__2_.mem_right_track_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__2_.mem_right_track_8.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__2_.mem_right_track_16.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_1.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__2_.mem_left_track_9.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_1__2_.mem_left_track_17.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_2__0_.mem_top_track_0.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_2.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_4.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_6.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_10.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_12.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_14.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_16.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_1.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_3.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_left_track_5.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_7.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_9.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_11.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_13.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_15.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_17.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_2__1_.mem_top_track_8.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_2__1_.mem_top_track_16.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_9.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_17.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.sb_2__1_.mem_left_track_1.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_3.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_5.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_7.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_9.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_11.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_13.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_15.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_17.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_1.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_3.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_5.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__2_.mem_left_track_7.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_9.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__2_.mem_left_track_11.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_13.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_15.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_17.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_1.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_2.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_3.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_4.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_5.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_6.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_7.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_1.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_2.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_3.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_4.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_5.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_6.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_7.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_1.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_2.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_1.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_2.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_3.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_4.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_5.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_6.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_7.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_0.mem_outb[0:5] = 6'b011101;
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_1.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_2.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_3.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_4.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_5.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_6.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_7.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_1.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_2.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_1.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_1.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_2.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_3.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_4.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_5.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_6.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_7.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_1.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_1.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_2.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_3.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_4.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_5.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_6.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_7.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_1__1_.mem_left_ipin_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_1__1_.mem_left_ipin_1.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_left_ipin_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_1.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_left_ipin_0.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_1.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_2.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_3.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_4.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_5.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_6.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_7.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.cby_2__1_.mem_right_ipin_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_2__1_.mem_right_ipin_1.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.cby_2__1_.mem_right_ipin_2.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_left_ipin_0.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_1.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_2.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_3.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_4.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_5.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_6.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_7.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_0.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_1.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_2.mem_outb[0:1] = 2'b10;
end
// ----- End assign bitstream to configuration memories -----
`else
// ----- Begin deposit bitstream to configuration memories -----
initial begin
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_1_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15], 16'b1010101000000000);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15], 16'b0101010111111111);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b010);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b101);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:7], 8'b00100100);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:7], 8'b11011011);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:7], 8'b10001000);
	$deposit(U0_formal_verification.grid_clb_2_1.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:7], 8'b01110111);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_out[0:15], {16{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_config_latch_mem.mem_outb[0:15], {16{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:2], 3'b001);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:2], 3'b110);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:7], 8'b00100001);
	$deposit(U0_formal_verification.grid_clb_2_2.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:7], 8'b11011110);
	$deposit(U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_top_1_3.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_top_2_3.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_right_3_1.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_right_3_2.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_bottom_1_0.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_bottom_2_0.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_left_0_1.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_out[0], {1{1'b1}});
	$deposit(U0_formal_verification.grid_io_left_0_2.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.iopad_config_latch_mem.mem_outb[0], {1{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_0.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_0.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_2.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_2.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_4.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_4.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_6.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_6.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_8.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_8.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_10.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_10.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_12.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_12.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_14.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_14.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_16.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_16.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_0.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_0.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_2.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_2.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_4.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_4.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_6.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_6.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_8.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_8.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_10.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_10.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_12.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_12.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_14.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_14.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_16.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_16.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_0.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_0.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_8.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_8.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_16.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_16.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_2.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_2.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_4.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_4.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_6.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_6.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_8.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_8.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_10.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_10.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_12.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_12.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_14.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_14.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_9.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_9.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_17.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_17.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_0.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_0.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_2.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_2.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_4.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_4.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_6.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_6.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_8.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_8.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_10.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_10.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_12.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_12.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_14.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_14.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_16.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_16.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_3.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_3.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_5.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_5.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_7.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_7.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_9.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_9.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_11.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_11.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_13.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_13.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_15.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_15.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_17.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_17.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_0.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_0.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_2.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_2.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_8.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_8.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_14.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_14.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_16.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_16.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_0.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_0.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_8.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_8.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_16.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_16.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_1.mem_out[0:5], 6'b010100);
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_1.mem_outb[0:5], 6'b101011);
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_9.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_9.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_17.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_17.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_0.mem_out[0:7], 8'b10001000);
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_0.mem_outb[0:7], 8'b01110111);
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_8.mem_out[0:7], 8'b10001000);
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_8.mem_outb[0:7], 8'b01110111);
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_16.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_16.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_0.mem_out[0:7], 8'b10001000);
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_0.mem_outb[0:7], 8'b01110111);
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_8.mem_out[0:7], 8'b10001000);
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_8.mem_outb[0:7], 8'b01110111);
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_16.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_16.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_out[0:7], 8'b00101000);
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_outb[0:7], 8'b11010111);
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_9.mem_out[0:7], 8'b10001000);
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_9.mem_outb[0:7], 8'b01110111);
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_17.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_17.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_1.mem_out[0:7], 8'b10001000);
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_1.mem_outb[0:7], 8'b01110111);
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_9.mem_out[0:7], 8'b10001000);
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_9.mem_outb[0:7], 8'b01110111);
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_17.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_17.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_0.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_0.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_8.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_8.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_16.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_16.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_3.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_3.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_5.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_5.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_7.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_7.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_9.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_9.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_11.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_11.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_13.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_13.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_15.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_15.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_17.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_17.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_1.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_1.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_9.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_9.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_17.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_17.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_0.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_0.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_2.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_2.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_4.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_4.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_6.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_6.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_8.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_8.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_10.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_10.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_12.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_12.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_14.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_14.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_16.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_16.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_1.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_1.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_3.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_3.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_5.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_5.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_7.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_7.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_9.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_9.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_11.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_11.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_13.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_13.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_15.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_15.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_17.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_17.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_0.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_0.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_8.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_8.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_16.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_16.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_9.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_9.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_17.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_17.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_1.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_1.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_3.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_3.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_5.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_5.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_7.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_7.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_9.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_9.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_11.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_11.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_13.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_13.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_15.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_15.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_17.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_17.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_3.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_3.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_5.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_5.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_7.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_7.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_9.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_9.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_11.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_11.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_13.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_13.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_15.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_15.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_17.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_17.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_1.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_1.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_3.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_3.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_5.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_5.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_7.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_7.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_9.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_9.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_11.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_11.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_13.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_13.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_15.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_15.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_17.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_17.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_1.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_1.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_2.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_2.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_3.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_3.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_4.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_4.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_5.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_5.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_6.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_6.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_7.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_7.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_0.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_0.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_1.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_1.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_2.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_top_ipin_2.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_3.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_3.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_4.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_4.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_5.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_5.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_6.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_6.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_7.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_7.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_0.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_0.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_1.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_1.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_2.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_top_ipin_2.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_1.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_1.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_2.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_2.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_3.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_3.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_4.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_4.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_5.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_5.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_6.mem_out[0:5], 6'b001100);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_6.mem_outb[0:5], 6'b110011);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_7.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_7.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_0.mem_out[0:5], 6'b100010);
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_0.mem_outb[0:5], 6'b011101);
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_1.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_1.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_2.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_top_ipin_2.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_3.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_3.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_4.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_4.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_5.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_5.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_6.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_6.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_7.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_7.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_0.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_0.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_1.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_1.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_2.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_top_ipin_2.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_0__1_.mem_left_ipin_0.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_0__1_.mem_left_ipin_0.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_0__1_.mem_left_ipin_1.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_0__1_.mem_left_ipin_1.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_1.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_1.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_2.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_2.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_3.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_3.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_4.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_4.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_5.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_5.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_6.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_6.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_7.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_7.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_0__2_.mem_left_ipin_0.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_0__2_.mem_left_ipin_0.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_0__2_.mem_left_ipin_1.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_0__2_.mem_left_ipin_1.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_1.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_1.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_2.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_2.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_3.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_3.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_4.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_4.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_5.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_5.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_6.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_6.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_7.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_7.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_1__1_.mem_left_ipin_0.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_1__1_.mem_left_ipin_0.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_1__1_.mem_left_ipin_1.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_1__1_.mem_left_ipin_1.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_left_ipin_0.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_1__2_.mem_left_ipin_0.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_1__2_.mem_left_ipin_1.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_1__2_.mem_left_ipin_1.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_0.mem_out[0:5], 6'b010100);
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_0.mem_outb[0:5], 6'b101011);
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_1.mem_out[0:5], 6'b010100);
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_1.mem_outb[0:5], 6'b101011);
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_2.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_2.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_3.mem_out[0:5], 6'b010100);
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_3.mem_outb[0:5], 6'b101011);
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_4.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_4.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_5.mem_out[0:5], 6'b010100);
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_5.mem_outb[0:5], 6'b101011);
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_6.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_6.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_7.mem_out[0:5], 6'b010100);
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_7.mem_outb[0:5], 6'b101011);
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_0.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_0.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_1.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_1.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_2.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_2.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_0.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_0.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_1.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_1.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_2.mem_out[0:5], 6'b010100);
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_2.mem_outb[0:5], 6'b101011);
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_3.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_3.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_4.mem_out[0:5], 6'b010100);
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_4.mem_outb[0:5], 6'b101011);
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_5.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_5.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_6.mem_out[0:5], 6'b010100);
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_6.mem_outb[0:5], 6'b101011);
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_7.mem_out[0:5], 6'b100100);
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_7.mem_outb[0:5], 6'b011011);
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_0.mem_out[0:5], 6'b010100);
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_0.mem_outb[0:5], 6'b101011);
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_1.mem_out[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_1.mem_outb[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_2.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_2.mem_outb[0:1], 2'b10);
end
// ----- End deposit bitstream to configuration memories -----
`endif
// ----- End load bitstream to configuration memories -----
endmodule
// ----- END Verilog module for and2_top_formal_verification -----

