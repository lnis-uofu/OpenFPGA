// Benchmark "TOP" written by ABC on Tue Mar  5 09:55:52 2019

module clma ( clk, 
    Pi416, Pi415, Pi414, Pi413, Pi412, Pi411, Pi410, Pi409, Pi408, Pi407,
    Pi406, Pi405, Pi404, Pi403, Pi402, Pi401, Pi400, Pi399, Pi398, Pi397,
    Pi396, Pi395, Pi394, Pi393, Pi392, Pi391, Pi390, Pi389, Pi388, Pi387,
    Pi386, Pi385, Pi384, Pi383, Pi382, Pi381, Pi380, Pi379, Pi378, Pi377,
    Pi376, Pi375, Pi374, Pi373, Pi372, Pi371, Pi370, Pi369, Pi368, Pi367,
    Pi366, Pi365, Pi364, Pi363, Pi362, Pi361, Pi360, Pi359, Pi358, Pi357,
    Pi356, Pi355, Pi354, Pi353, Pi352, Pi351, Pi350, Pi349, Pi348, Pi347,
    Pi346, Pi345, Pi344, Pi343, Pi342, Pi341, Pi340, Pi339, Pi338, Pi337,
    Pi336, Pi335, Pi334, Pi333, Pi332, Pi331, Pi330, Pi329, Pi328, Pi327,
    Pi326, Pi325, Pi324, Pi323, Pi322, Pi321, Pi320, Pi319, Pi318, Pi317,
    Pi316, Pi315, Pi314, Pi313, Pi312, Pi311, Pi310, Pi309, Pi308, Pi307,
    Pi306, Pi305, Pi304, Pi303, Pi302, Pi301, Pi300, Pi299, Pi298, Pi297,
    Pi296, Pi295, Pi294, Pi293, Pi292, Pi291, Pi290, Pi289, Pi288, Pi287,
    Pi286, Pi285, Pi284, Pi283, Pi282, Pi281, Pi280, Pi279, Pi278, Pi277,
    Pi276, Pi275, Pi274, Pi273, Pi272, Pi271, Pi270, Pi269, Pi268, Pi267,
    Pi266, Pi265, Pi264, Pi263, Pi262, Pi261, Pi260, Pi259, Pi258, Pi257,
    Pi256, Pi255, Pi254, Pi253, Pi252, Pi251, Pi250, Pi249, Pi248, Pi247,
    Pi246, Pi245, Pi244, Pi243, Pi242, Pi241, Pi240, Pi239, Pi238, Pi237,
    Pi236, Pi235, Pi234, Pi233, Pi232, Pi231, Pi230, Pi229, Pi228, Pi227,
    Pi226, Pi225, Pi224, Pi223, Pi222, Pi221, Pi220, Pi219, Pi218, Pi217,
    Pi216, Pi215, Pi214, Pi213, Pi212, Pi211, Pi210, Pi209, Pi208, Pi207,
    Pi206, Pi205, Pi204, Pi203, Pi202, Pi201, Pi200, Pi199, Pi198, Pi197,
    Pi196, Pi195, Pi194, Pi193, Pi192, Pi191, Pi190, Pi189, Pi188, Pi187,
    Pi186, Pi185, Pi184, Pi183, Pi182, Pi181, Pi180, Pi179, Pi178, Pi177,
    Pi176, Pi175, Pi174, Pi173, Pi172, Pi171, Pi170, Pi169, Pi168, Pi167,
    Pi166, Pi165, Pi164, Pi163, Pi162, Pi161, Pi160, Pi159, Pi158, Pi157,
    Pi156, Pi155, Pi154, Pi153, Pi152, Pi151, Pi150, Pi149, Pi148, Pi147,
    Pi146, Pi145, Pi144, Pi143, Pi142, Pi141, Pi140, Pi139, Pi138, Pi137,
    Pi136, Pi135, Pi134, Pi133, Pi132, Pi131, Pi130, Pi129, Pi128, Pi127,
    Pi126, Pi125, Pi124, Pi123, Pi122, Pi121, Pi120, Pi119, Pi118, Pi117,
    Pi116, Pi115, Pi114, Pi113, Pi112, Pi111, Pi110, Pi109, Pi108, Pi107,
    Pi106, Pi105, Pi104, Pi103, Pi102, Pi101, Pi100, Pi99, Pi98, Pi97,
    Pi96, Pi95, Pi94, Pi93, Pi92, Pi91, Pi90, Pi89, Pi88, Pi87, Pi86, Pi85,
    Pi84, Pi83, Pi82, Pi81, Pi80, Pi79, Pi78, Pi77, Pi76, Pi75, Pi74, Pi73,
    Pi72, Pi71, Pi70, Pi69, Pi68, Pi67, Pi66, Pi65, Pi64, Pi63, Pi62, Pi61,
    Pi60, Pi59, Pi58, Pi57, Pi56, Pi55, Pi54, Pi53, Pi52, Pi51, Pi50, Pi49,
    Pi28, Pi27, Pi26, Pi25, Pi24, Pi23, Pi22, Pi21, Pi20, Pi19, Pi18, Pi17,
    Pi16, Pi15, 
    P__cmxir_1, P__cmxir_0, P__cmxig_1, P__cmxig_0, P__cmxcl_1, P__cmxcl_0,
    P__cmx1ad_35, P__cmx1ad_34, P__cmx1ad_33, P__cmx1ad_32, P__cmx1ad_31,
    P__cmx1ad_30, P__cmx1ad_29, P__cmx1ad_28, P__cmx1ad_27, P__cmx1ad_26,
    P__cmx1ad_25, P__cmx1ad_24, P__cmx1ad_23, P__cmx1ad_22, P__cmx1ad_21,
    P__cmx1ad_20, P__cmx1ad_19, P__cmx1ad_18, P__cmx1ad_17, P__cmx1ad_16,
    P__cmx1ad_15, P__cmx1ad_14, P__cmx1ad_13, P__cmx1ad_12, P__cmx1ad_11,
    P__cmx1ad_10, P__cmx1ad_9, P__cmx1ad_8, P__cmx1ad_7, P__cmx1ad_6,
    P__cmx1ad_5, P__cmx1ad_4, P__cmx1ad_3, P__cmx1ad_2, P__cmx1ad_1,
    P__cmx1ad_0, P__cmx0ad_35, P__cmx0ad_34, P__cmx0ad_33, P__cmx0ad_32,
    P__cmx0ad_31, P__cmx0ad_30, P__cmx0ad_29, P__cmx0ad_28, P__cmx0ad_27,
    P__cmx0ad_26, P__cmx0ad_25, P__cmx0ad_24, P__cmx0ad_23, P__cmx0ad_22,
    P__cmx0ad_21, P__cmx0ad_20, P__cmx0ad_19, P__cmx0ad_18, P__cmx0ad_17,
    P__cmx0ad_16, P__cmx0ad_15, P__cmx0ad_14, P__cmx0ad_13, P__cmx0ad_12,
    P__cmx0ad_11, P__cmx0ad_10, P__cmx0ad_9, P__cmx0ad_8, P__cmx0ad_7,
    P__cmx0ad_6, P__cmx0ad_5, P__cmx0ad_4, P__cmx0ad_3, P__cmx0ad_2,
    P__cmx0ad_1, P__cmx0ad_0, P__cmnxcp_1, P__cmnxcp_0, P__cmndst1p0,
    P__cmndst0p0  );
  input  Pi416, Pi415, Pi414, Pi413, Pi412, Pi411, Pi410, Pi409, Pi408,
    Pi407, Pi406, Pi405, Pi404, Pi403, Pi402, Pi401, Pi400, Pi399, Pi398,
    Pi397, Pi396, Pi395, Pi394, Pi393, Pi392, Pi391, Pi390, Pi389, Pi388,
    Pi387, Pi386, Pi385, Pi384, Pi383, Pi382, Pi381, Pi380, Pi379, Pi378,
    Pi377, Pi376, Pi375, Pi374, Pi373, Pi372, Pi371, Pi370, Pi369, Pi368,
    Pi367, Pi366, Pi365, Pi364, Pi363, Pi362, Pi361, Pi360, Pi359, Pi358,
    Pi357, Pi356, Pi355, Pi354, Pi353, Pi352, Pi351, Pi350, Pi349, Pi348,
    Pi347, Pi346, Pi345, Pi344, Pi343, Pi342, Pi341, Pi340, Pi339, Pi338,
    Pi337, Pi336, Pi335, Pi334, Pi333, Pi332, Pi331, Pi330, Pi329, Pi328,
    Pi327, Pi326, Pi325, Pi324, Pi323, Pi322, Pi321, Pi320, Pi319, Pi318,
    Pi317, Pi316, Pi315, Pi314, Pi313, Pi312, Pi311, Pi310, Pi309, Pi308,
    Pi307, Pi306, Pi305, Pi304, Pi303, Pi302, Pi301, Pi300, Pi299, Pi298,
    Pi297, Pi296, Pi295, Pi294, Pi293, Pi292, Pi291, Pi290, Pi289, Pi288,
    Pi287, Pi286, Pi285, Pi284, Pi283, Pi282, Pi281, Pi280, Pi279, Pi278,
    Pi277, Pi276, Pi275, Pi274, Pi273, Pi272, Pi271, Pi270, Pi269, Pi268,
    Pi267, Pi266, Pi265, Pi264, Pi263, Pi262, Pi261, Pi260, Pi259, Pi258,
    Pi257, Pi256, Pi255, Pi254, Pi253, Pi252, Pi251, Pi250, Pi249, Pi248,
    Pi247, Pi246, Pi245, Pi244, Pi243, Pi242, Pi241, Pi240, Pi239, Pi238,
    Pi237, Pi236, Pi235, Pi234, Pi233, Pi232, Pi231, Pi230, Pi229, Pi228,
    Pi227, Pi226, Pi225, Pi224, Pi223, Pi222, Pi221, Pi220, Pi219, Pi218,
    Pi217, Pi216, Pi215, Pi214, Pi213, Pi212, Pi211, Pi210, Pi209, Pi208,
    Pi207, Pi206, Pi205, Pi204, Pi203, Pi202, Pi201, Pi200, Pi199, Pi198,
    Pi197, Pi196, Pi195, Pi194, Pi193, Pi192, Pi191, Pi190, Pi189, Pi188,
    Pi187, Pi186, Pi185, Pi184, Pi183, Pi182, Pi181, Pi180, Pi179, Pi178,
    Pi177, Pi176, Pi175, Pi174, Pi173, Pi172, Pi171, Pi170, Pi169, Pi168,
    Pi167, Pi166, Pi165, Pi164, Pi163, Pi162, Pi161, Pi160, Pi159, Pi158,
    Pi157, Pi156, Pi155, Pi154, Pi153, Pi152, Pi151, Pi150, Pi149, Pi148,
    Pi147, Pi146, Pi145, Pi144, Pi143, Pi142, Pi141, Pi140, Pi139, Pi138,
    Pi137, Pi136, Pi135, Pi134, Pi133, Pi132, Pi131, Pi130, Pi129, Pi128,
    Pi127, Pi126, Pi125, Pi124, Pi123, Pi122, Pi121, Pi120, Pi119, Pi118,
    Pi117, Pi116, Pi115, Pi114, Pi113, Pi112, Pi111, Pi110, Pi109, Pi108,
    Pi107, Pi106, Pi105, Pi104, Pi103, Pi102, Pi101, Pi100, Pi99, Pi98,
    Pi97, Pi96, Pi95, Pi94, Pi93, Pi92, Pi91, Pi90, Pi89, Pi88, Pi87, Pi86,
    Pi85, Pi84, Pi83, Pi82, Pi81, Pi80, Pi79, Pi78, Pi77, Pi76, Pi75, Pi74,
    Pi73, Pi72, Pi71, Pi70, Pi69, Pi68, Pi67, Pi66, Pi65, Pi64, Pi63, Pi62,
    Pi61, Pi60, Pi59, Pi58, Pi57, Pi56, Pi55, Pi54, Pi53, Pi52, Pi51, Pi50,
    Pi49, Pi28, Pi27, Pi26, Pi25, Pi24, Pi23, Pi22, Pi21, Pi20, Pi19, Pi18,
    Pi17, Pi16, Pi15, clk;
  output P__cmxir_1, P__cmxir_0, P__cmxig_1, P__cmxig_0, P__cmxcl_1,
    P__cmxcl_0, P__cmx1ad_35, P__cmx1ad_34, P__cmx1ad_33, P__cmx1ad_32,
    P__cmx1ad_31, P__cmx1ad_30, P__cmx1ad_29, P__cmx1ad_28, P__cmx1ad_27,
    P__cmx1ad_26, P__cmx1ad_25, P__cmx1ad_24, P__cmx1ad_23, P__cmx1ad_22,
    P__cmx1ad_21, P__cmx1ad_20, P__cmx1ad_19, P__cmx1ad_18, P__cmx1ad_17,
    P__cmx1ad_16, P__cmx1ad_15, P__cmx1ad_14, P__cmx1ad_13, P__cmx1ad_12,
    P__cmx1ad_11, P__cmx1ad_10, P__cmx1ad_9, P__cmx1ad_8, P__cmx1ad_7,
    P__cmx1ad_6, P__cmx1ad_5, P__cmx1ad_4, P__cmx1ad_3, P__cmx1ad_2,
    P__cmx1ad_1, P__cmx1ad_0, P__cmx0ad_35, P__cmx0ad_34, P__cmx0ad_33,
    P__cmx0ad_32, P__cmx0ad_31, P__cmx0ad_30, P__cmx0ad_29, P__cmx0ad_28,
    P__cmx0ad_27, P__cmx0ad_26, P__cmx0ad_25, P__cmx0ad_24, P__cmx0ad_23,
    P__cmx0ad_22, P__cmx0ad_21, P__cmx0ad_20, P__cmx0ad_19, P__cmx0ad_18,
    P__cmx0ad_17, P__cmx0ad_16, P__cmx0ad_15, P__cmx0ad_14, P__cmx0ad_13,
    P__cmx0ad_12, P__cmx0ad_11, P__cmx0ad_10, P__cmx0ad_9, P__cmx0ad_8,
    P__cmx0ad_7, P__cmx0ad_6, P__cmx0ad_5, P__cmx0ad_4, P__cmx0ad_3,
    P__cmx0ad_2, P__cmx0ad_1, P__cmx0ad_0, P__cmnxcp_1, P__cmnxcp_0,
    P__cmndst1p0, P__cmndst0p0;
  reg Ni48, Ni47, Ni46, Ni45, Ni44, Ni43, Ni42, Ni41, Ni40, Ni39, Ni38,
    Ni37, Ni36, Ni35, Ni34, Ni33, Ni32, Ni31, Ni30, n18, Ni14, Ni13, Ni12,
    Ni11, Ni10, Ni9, Ni8, Ni7, Ni6, Ni5, Ni4, Ni3, Ni2;
  wire n646, n648, n649, n651, n653, n654, n655, n656, n658, n660, n662,
    n663, n664, n665, n666, n668, n670, n672, n674, n675, n676, n677, n678,
    n679, n681, n683, n684, n686, n688, n689, n690, n691, n692, n693, n694,
    n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
    n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
    n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
    n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
    n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
    n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
    n767, n768, n770, n772, n773, n774, n776, n778, n780, n781, n783, n784,
    n785, n786, n787, n788, n789, n790, n792, n793, n794, n795, n796, n797,
    n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
    n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
    n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
    n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
    n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
    n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
    n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936_1, n937, n938, n939, n940,
    n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
    n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
    n965, n966, n967, n968, n969, n970, n971_1, n972, n973, n974, n975,
    n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986_1,
    n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
    n999, n1000, n1001_1, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
    n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
    n1019, n1020, n1021_1, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
    n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036_1, n1037, n1038,
    n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
    n1049, n1050, n1051_1, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
    n1059, n1060, n1061_1, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
    n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076_1, n1077, n1078,
    n1079, n1080, n1081_1, n1082, n1083, n1084, n1085_1, n1086, n1087,
    n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
    n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
    n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
    n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
    n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
    n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
    n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
    n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
    n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
    n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
    n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
    n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
    n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
    n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
    n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
    n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
    n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
    n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
    n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
    n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
    n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
    n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
    n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
    n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
    n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
    n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
    n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
    n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
    n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
    n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
    n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
    n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
    n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
    n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
    n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
    n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
    n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
    n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
    n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
    n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
    n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
    n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
    n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
    n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
    n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
    n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
    n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
    n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
    n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
    n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
    n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
    n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
    n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
    n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
    n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
    n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
    n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
    n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
    n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
    n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
    n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
    n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
    n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
    n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
    n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
    n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
    n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
    n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
    n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
    n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
    n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
    n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
    n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
    n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
    n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
    n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
    n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
    n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
    n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
    n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
    n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
    n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
    n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
    n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
    n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
    n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
    n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
    n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
    n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
    n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
    n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
    n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
    n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
    n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
    n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
    n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
    n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
    n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
    n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
    n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
    n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
    n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
    n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
    n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
    n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
    n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
    n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
    n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
    n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
    n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
    n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
    n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
    n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
    n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
    n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
    n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
    n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
    n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
    n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
    n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
    n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
    n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
    n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
    n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
    n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
    n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
    n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
    n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
    n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
    n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
    n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
    n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
    n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
    n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
    n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
    n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
    n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
    n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
    n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
    n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
    n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
    n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
    n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
    n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
    n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
    n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
    n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
    n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
    n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
    n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
    n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
    n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
    n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
    n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
    n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
    n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
    n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
    n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
    n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
    n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
    n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
    n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
    n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
    n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
    n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
    n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
    n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
    n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
    n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
    n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
    n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
    n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
    n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
    n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
    n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
    n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
    n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
    n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
    n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
    n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
    n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
    n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
    n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
    n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
    n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
    n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
    n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
    n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
    n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
    n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
    n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
    n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
    n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
    n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
    n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
    n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
    n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
    n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
    n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
    n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
    n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
    n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
    n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
    n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
    n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
    n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
    n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
    n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
    n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
    n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
    n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
    n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
    n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
    n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
    n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
    n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
    n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
    n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
    n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
    n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
    n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
    n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
    n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
    n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
    n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
    n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
    n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
    n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
    n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
    n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
    n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
    n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
    n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
    n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
    n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
    n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
    n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
    n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
    n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
    n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
    n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
    n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
    n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
    n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
    n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
    n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
    n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
    n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
    n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
    n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
    n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
    n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
    n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
    n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
    n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
    n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
    n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
    n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
    n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
    n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
    n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
    n3758, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
    n3769, n3770, n3771, n3772, n3773, n3775, n3777, n3779, n3780, n3781,
    n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
    n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
    n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
    n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
    n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
    n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
    n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
    n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
    n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
    n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
    n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
    n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
    n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
    n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
    n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
    n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
    n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
    n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
    n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
    n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
    n3983, n3984, n3985, n3986, n3987, n3989, n3990, n3991, n3992, n3993,
    n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
    n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
    n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
    n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
    n4034, n4035, n4037, n4038, n4039, n4040, n4042, n4044, n4045, n4046,
    n4048, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
    n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
    n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
    n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
    n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
    n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
    n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
    n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
    n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
    n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
    n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
    n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
    n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
    n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
    n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
    n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
    n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
    n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
    n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
    n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
    n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
    n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
    n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
    n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
    n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
    n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
    n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
    n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
    n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
    n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
    n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
    n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
    n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
    n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
    n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
    n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
    n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
    n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
    n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
    n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
    n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
    n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
    n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
    n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
    n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
    n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
    n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
    n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
    n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
    n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
    n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
    n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
    n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
    n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
    n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
    n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
    n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
    n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
    n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
    n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
    n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
    n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
    n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
    n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
    n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
    n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
    n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
    n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
    n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
    n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
    n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
    n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
    n4769, n4770, n4771, n4772, n4773, n4774, n4775, n931_1, n936, n941_1,
    n946_1, n951_1, n956_1, n961_1, n966_1, n971, n976_1, n981_1, n986,
    n991_1, n996_1, n1001, n1006_1, n1011_1, n1016_1, n1021, n1026_1,
    n1031_1, n1036, n1041_1, n1046_1, n1051, n1056_1, n1061, n1066_1,
    n1071_1, n1076, n1081, n1085, n1090_1;
  assign P__cmxir_1 = n785 & ~n3327 & ~n3707;
  assign P__cmxir_0 = ~n773 & ~n3659;
  assign P__cmxig_1 = ~n785;
  assign P__cmxig_0 = ~n3950;
  assign P__cmxcl_1 = ~n3707;
  assign P__cmxcl_0 = ~n3707;
  assign P__cmx1ad_35 = 1'b0;
  assign P__cmx1ad_34 = 1'b0;
  assign P__cmx1ad_33 = 1'b0;
  assign P__cmx1ad_32 = 1'b0;
  assign P__cmx1ad_31 = Pi255 & ~n3985;
  assign P__cmx1ad_30 = Pi254 & ~n3985;
  assign P__cmx1ad_29 = Pi253 & ~n3985;
  assign P__cmx1ad_28 = Pi252 & ~n3985;
  assign P__cmx1ad_27 = Pi251 & ~n3985;
  assign P__cmx1ad_26 = Pi250 & ~n3985;
  assign P__cmx1ad_25 = Pi249 & ~n3985;
  assign P__cmx1ad_24 = Pi248 & ~n3985;
  assign P__cmx1ad_23 = Pi247 & ~n3985;
  assign P__cmx1ad_22 = Pi246 & ~n3985;
  assign P__cmx1ad_21 = Pi245 & ~n3985;
  assign P__cmx1ad_20 = Pi244 & ~n3985;
  assign P__cmx1ad_19 = Pi243 & ~n3985;
  assign P__cmx1ad_18 = Pi242 & ~n3985;
  assign P__cmx1ad_17 = Pi241 & ~n3985;
  assign P__cmx1ad_16 = Pi240 & ~n3985;
  assign P__cmx1ad_15 = ~n3985 & Pi27 & Pi26;
  assign P__cmx1ad_14 = ~n4051;
  assign P__cmx1ad_13 = n789 & ~n3985;
  assign P__cmx1ad_12 = ~n4760;
  assign P__cmx1ad_11 = 1'b0;
  assign P__cmx1ad_10 = 1'b0;
  assign P__cmx1ad_9 = ~n3985;
  assign P__cmx1ad_8 = 1'b0;
  assign P__cmx1ad_7 = Pi239 & ~n3985;
  assign P__cmx1ad_6 = Pi238 & ~n3985;
  assign P__cmx1ad_5 = Pi237 & ~n3985;
  assign P__cmx1ad_4 = Pi236 & ~n3985;
  assign P__cmx1ad_3 = Pi235 & ~n3985;
  assign P__cmx1ad_2 = Pi234 & ~n3985;
  assign P__cmx1ad_1 = Pi233 & ~n3985;
  assign P__cmx1ad_0 = Pi232 & ~n3985;
  assign P__cmx0ad_35 = 1'b0;
  assign P__cmx0ad_34 = 1'b0;
  assign P__cmx0ad_33 = 1'b0;
  assign P__cmx0ad_32 = 1'b0;
  assign P__cmx0ad_31 = Pi72 & ~n3986;
  assign P__cmx0ad_30 = Pi71 & ~n3986;
  assign P__cmx0ad_29 = Pi70 & ~n3986;
  assign P__cmx0ad_28 = Pi69 & ~n3986;
  assign P__cmx0ad_27 = Pi68 & ~n3986;
  assign P__cmx0ad_26 = Pi67 & ~n3986;
  assign P__cmx0ad_25 = Pi66 & ~n3986;
  assign P__cmx0ad_24 = Pi65 & ~n3986;
  assign P__cmx0ad_23 = Pi64 & ~n3986;
  assign P__cmx0ad_22 = Pi63 & ~n3986;
  assign P__cmx0ad_21 = Pi62 & ~n3986;
  assign P__cmx0ad_20 = Pi61 & ~n3986;
  assign P__cmx0ad_19 = Pi60 & ~n3986;
  assign P__cmx0ad_18 = Pi59 & ~n3986;
  assign P__cmx0ad_17 = Pi58 & ~n3986;
  assign P__cmx0ad_16 = Pi57 & ~n3986;
  assign P__cmx0ad_15 = ~n3986 & Pi24 & Pi23;
  assign P__cmx0ad_14 = ~n4052;
  assign P__cmx0ad_13 = n788 & ~n3986;
  assign P__cmx0ad_12 = ~n4762;
  assign P__cmx0ad_11 = 1'b0;
  assign P__cmx0ad_10 = 1'b0;
  assign P__cmx0ad_9 = ~n3986;
  assign P__cmx0ad_8 = 1'b0;
  assign P__cmx0ad_7 = Pi56 & ~n3986;
  assign P__cmx0ad_6 = Pi55 & ~n3986;
  assign P__cmx0ad_5 = Pi54 & ~n3986;
  assign P__cmx0ad_4 = Pi53 & ~n3986;
  assign P__cmx0ad_3 = Pi52 & ~n3986;
  assign P__cmx0ad_2 = Pi51 & ~n3986;
  assign P__cmx0ad_1 = Pi50 & ~n3986;
  assign P__cmx0ad_0 = Pi49 & ~n3986;
  assign P__cmnxcp_1 = ~n787;
  assign P__cmnxcp_0 = ~n786;
  assign P__cmndst1p0 = n784 & ~n3754;
  assign P__cmndst0p0 = n783 & ~n3984;
  assign n646 = ~n3662 & (~Ni48 | (~Pi22 & n3663));
  assign n931_1 = ~n646;
  assign n648 = ~n904 & n3185 & (Pi20 | n3186);
  assign n649 = Ni46 & (Pi21 | (~Ni32 & ~n2416));
  assign n941_1 = n648 | n649;
  assign n651 = ~n3829 & (~Ni44 | ~n3751);
  assign n951_1 = ~n651;
  assign n653 = Ni44 ^ ~Ni39;
  assign n654 = n653 & Ni38;
  assign n655 = n653 & Ni32 & (Ni37 | n654);
  assign n656 = n3190 & (n2398 | ~Ni41);
  assign n966_1 = ~n656;
  assign n658 = n3188 & (n2398 | ~Ni40);
  assign n971 = ~n658;
  assign n660 = n2391 & (n665 | ~Ni39);
  assign n976_1 = ~n660;
  assign n662 = ~n3183 & (~n1241 | ~n2389) & ~n3864;
  assign n663 = ~n1322 & ~n3183 & (n808 | ~n995);
  assign n664 = Pi15 & ~n741 & ~n3984;
  assign n665 = ~Ni32 & n2406;
  assign n666 = ~n3984 & ~n3183 & n3184;
  assign n981_1 = ~n4774 | n665 | n666 | n664 | n662 | n663;
  assign n668 = ~n2404 & (~Ni36 | n2398) & n2405;
  assign n991_1 = ~n668;
  assign n670 = ~n2396 & n2397 & (~Ni35 | n2398);
  assign n996_1 = ~n670;
  assign n672 = ~n2388 & ~n3806 & (~Ni34 | ~n3707);
  assign n1001 = ~n672;
  assign n674 = ~Ni42 & (~Ni44 | ~n738);
  assign n675 = ~Ni42 & (Ni44 | ~n738);
  assign n676 = ~Ni47 & ~Ni45;
  assign n677 = ~Ni42 | Ni43;
  assign n678 = n676 & n677;
  assign n679 = n3658 & (n3659 | (~n3657 & n3660));
  assign n1006_1 = ~n679;
  assign n681 = ~n3181 & n3182 & (~n2073 | ~n4431);
  assign n1011_1 = ~n681;
  assign n683 = n2078 & (~n678 | ~n814) & ~n3707;
  assign n684 = ~n3707 & n2254 & ~Ni32 & ~Ni30;
  assign n1016_1 = Ni31 | n683 | n684;
  assign n686 = n2076 & n2077 & (~Ni30 | ~n3707);
  assign n1021 = ~n686;
  assign n688 = n1393 & n1394 & (n689 | n1395);
  assign n689 = n4769 & n713;
  assign n690 = ~n814 | ~Ni36;
  assign n691 = n688 & ~n1539 & (n689 | n690);
  assign n692 = n1393 & n1394 & (n693 | n1398);
  assign n693 = n4770 & n713;
  assign n694 = n692 & ~n1539 & (n690 | n693);
  assign n695 = n985 & (n697 | ~Ni38);
  assign n696 = ~n1539 & (n744 | ~Ni35);
  assign n697 = n713 & (n689 | ~Ni40);
  assign n698 = Ni37 | ~Ni36;
  assign n699 = n695 & n696 & (n697 | n698);
  assign n700 = n985 & (n702 | ~Ni38);
  assign n701 = ~n1539 & (n746 | ~Ni35);
  assign n702 = n713 & (n693 | ~Ni40);
  assign n703 = n700 & n701 & (n702 | n698);
  assign n704 = n985 & (n706 | ~Ni38);
  assign n705 = ~n1539 & (Ni35 | n748);
  assign n706 = n713 & (Ni40 | n689);
  assign n707 = n704 & n705 & (n706 | n698);
  assign n708 = n985 & (n710 | ~Ni38);
  assign n709 = ~n1539 & (Ni35 | n750);
  assign n710 = n713 & (Ni40 | n693);
  assign n711 = n708 & n709 & (n710 | n698);
  assign n712 = n985 & (n713 | ~Ni38);
  assign n713 = n738 & (n1351 | ~Ni41);
  assign n714 = n712 & ~n1539 & (n698 | n713);
  assign n715 = n1393 & n1394 & (n716 | n1395);
  assign n716 = n738 & n4769;
  assign n717 = n715 & ~n1539 & (n690 | n716);
  assign n718 = n1393 & n1394 & (n719 | n1398);
  assign n719 = n738 & n4770;
  assign n720 = n718 & ~n1539 & (n690 | n719);
  assign n721 = n985 & (n723 | ~Ni38);
  assign n722 = (~Ni35 | n754) & ~n1539;
  assign n723 = n738 & (n716 | ~Ni40);
  assign n724 = n721 & n722 & (n723 | n698);
  assign n725 = n985 & (n727 | ~Ni38);
  assign n726 = (~Ni35 | n756) & ~n1539;
  assign n727 = n738 & (n719 | ~Ni40);
  assign n728 = n725 & n726 & (n727 | n698);
  assign n729 = n985 & (n731 | ~Ni38);
  assign n730 = ~n1539 & (Ni35 | n758);
  assign n731 = n738 & (Ni40 | n716);
  assign n732 = n729 & n730 & (n731 | n698);
  assign n733 = n985 & (n735 | ~Ni38);
  assign n734 = ~n1539 & (Ni35 | n760);
  assign n735 = n738 & (Ni40 | n719);
  assign n736 = n733 & n734 & (n735 | n698);
  assign n737 = n985 & (n738 | ~Ni38);
  assign n738 = n676 & ~Ni43;
  assign n739 = n737 & ~n1539 & (n698 | n738);
  assign n740 = n985 & ~n1539;
  assign n741 = ~Ni36 | ~Ni38;
  assign n742 = n688 & n740 & (n689 | n741);
  assign n743 = n692 & n740 & (n693 | n741);
  assign n744 = n697 | n817;
  assign n745 = n695 & ~n1539 & (n744 | ~Ni35);
  assign n746 = n702 | n853;
  assign n747 = n700 & ~n1539 & (n746 | ~Ni35);
  assign n748 = n706 | n817;
  assign n749 = n704 & ~n1539 & (Ni35 | n748);
  assign n750 = n710 | n853;
  assign n751 = n708 & ~n1539 & (Ni35 | n750);
  assign n752 = n740 & n715 & (n716 | n741);
  assign n753 = n740 & n718 & (n719 | n741);
  assign n754 = n723 | n817;
  assign n755 = n721 & ~n1539 & (~Ni35 | n754);
  assign n756 = n727 | n853;
  assign n757 = n725 & ~n1539 & (~Ni35 | n756);
  assign n758 = n731 | n817;
  assign n759 = n729 & ~n1539 & (Ni35 | n758);
  assign n760 = n735 | n853;
  assign n761 = n733 & ~n1539 & (Ni35 | n760);
  assign n762 = Ni47 | n923;
  assign n763 = (~Ni44 | n762) & ~Ni41;
  assign n764 = Ni45 | n923;
  assign n765 = (~Ni44 | n764) & ~Ni41;
  assign n766 = ~Ni41 & (Ni44 | n762);
  assign n767 = ~Ni41 & (Ni44 | n764);
  assign n768 = ~n3731 & (~Ni14 | (n3711 & ~Ni2));
  assign n1031_1 = ~n768;
  assign n770 = n3726 & (~Ni13 | (~n3707 & ~n3727));
  assign n1036 = ~n770;
  assign n772 = ~Pi25 | Ni10;
  assign n773 = n772 & ~Ni9 & (~Ni10 | ~n3950);
  assign n774 = n3718 & (~Ni9 | (~n3707 & ~n3957));
  assign n1056_1 = ~n774;
  assign n776 = (n2403 | n3707) & (~Ni8 | n3715);
  assign n1061 = ~n776;
  assign n778 = n3713 & (Ni6 | n3712) & ~n4756;
  assign n1071_1 = ~n778;
  assign n780 = Ni6 & ~n3843 & (~n3668 | ~n3982);
  assign n781 = n3709 & n3710 & (n2418 | n3708);
  assign n1076 = ~n781;
  assign n783 = ~Ni37 & Ni38;
  assign n784 = ~Ni32 | ~Ni30;
  assign n785 = ~n18 | ~Ni33;
  assign n786 = n3770 & n3771 & (n3769 | n3707);
  assign n787 = ~n3763 & (n3707 | n3762) & n3764;
  assign n788 = Pi23 | Pi24;
  assign n789 = Pi26 | Pi27;
  assign n790 = n3751 & (~n784 | (n3752 & n3753));
  assign n956_1 = ~n790;
  assign n792 = Ni34 & (Ni30 | Ni32 | Ni31);
  assign n793 = ~Pi21 | ~n2643;
  assign n794 = Ni30 & n793 & (n788 | ~n1463);
  assign n795 = Pi24 | ~Pi23;
  assign n796 = Ni30 & n793 & (n795 | ~n1463);
  assign n797 = ~n3795 | n3956 | n3973;
  assign n798 = ~n1919 & (n797 | ~n4771);
  assign n799 = ~n2254 & (n797 | ~n3539 | ~n4771);
  assign n800 = n3956 | n3751;
  assign n801 = ~Ni32 | ~Ni31;
  assign n802 = n800 & n801;
  assign n803 = n3811 & n2430;
  assign n804 = ~n2420 & (n803 | ~Ni33);
  assign n805 = ~n2420 & (n803 | Ni33);
  assign n806 = (~n655 | Ni31) & ~n784;
  assign n807 = n3283 & (~Pi20 | ~n3977);
  assign n808 = ~Ni35 & ~Ni30;
  assign n809 = n797 | ~n4771;
  assign n810 = Pi22 & (n809 | ~n3539);
  assign n811 = n2419 & (Ni45 | n2420);
  assign n812 = n801 & ~n3829;
  assign n813 = n811 & n812;
  assign n814 = ~Ni37 | Ni38;
  assign n815 = n881 & (Ni40 | n1048);
  assign n816 = n814 & (~Ni37 | n815);
  assign n817 = ~n3194 | n3852;
  assign n818 = n678 & (n815 | n817);
  assign n819 = n678 & n816 & (~n783 | n815);
  assign n820 = (n815 | n698) & (n819 | n2434);
  assign n821 = n816 & n820 & (Ni35 | n818);
  assign n822 = ~Ni37 & (Ni36 | (n676 & ~n3194));
  assign n823 = n1082 | n1083;
  assign n824 = ~Ni36 & n822;
  assign n825 = Ni35 | n2438;
  assign n826 = n823 & (n824 | n825);
  assign n827 = n883 & (Ni40 | n1051_1);
  assign n828 = n814 & (~Ni37 | n827);
  assign n829 = n3849 | n3854;
  assign n830 = n829 & n828 & (n827 | n817);
  assign n831 = Ni38 | n3849;
  assign n832 = n828 & (~n783 | n827) & n831;
  assign n833 = (n827 | n1052) & (n828 | n886);
  assign n834 = (n832 | n3856) & (n830 | n992);
  assign n835 = n833 & n834;
  assign n836 = n889 & (Ni40 | n1055);
  assign n837 = n814 & (~Ni37 | n836);
  assign n838 = n3874 | n3854;
  assign n839 = n838 & n837 & (n836 | n817);
  assign n840 = Ni38 | n3874;
  assign n841 = n837 & (~n783 | n836) & n840;
  assign n842 = (n839 | n995) & (n837 | n891);
  assign n843 = (n841 | n3851) & (n836 | n1056);
  assign n844 = n842 & n843;
  assign n845 = n835 & n844;
  assign n846 = (n845 | n3850) & (n821 | n896);
  assign n847 = Ni32 | n1355;
  assign n848 = n826 & n846 & (n815 | n847);
  assign n849 = n18 | ~n1539;
  assign n850 = n849 & n848 & (n18 | n821);
  assign n851 = n881 & (Ni40 | n1064);
  assign n852 = n814 & (~Ni37 | n851);
  assign n853 = ~n3195 | n3852;
  assign n854 = n678 & (n851 | n853);
  assign n855 = n678 & n852 & (~n783 | n851);
  assign n856 = (n851 | n698) & (n855 | n2434);
  assign n857 = n852 & n856 & (Ni35 | n854);
  assign n858 = ~Ni37 & (Ni36 | (n676 & ~n3195));
  assign n859 = ~Ni36 & n858;
  assign n860 = n823 & (n859 | n825);
  assign n861 = n883 & (Ni40 | n1067);
  assign n862 = n814 & (~Ni37 | n861);
  assign n863 = n3849 | n3855;
  assign n864 = n863 & n862 & (n861 | n853);
  assign n865 = n831 & n862 & (~n783 | n861);
  assign n866 = (n861 | n1052) & (n862 | n886);
  assign n867 = (n865 | n3856) & (n864 | n992);
  assign n868 = n866 & n867;
  assign n869 = n889 & (Ni40 | n1070);
  assign n870 = n814 & (~Ni37 | n869);
  assign n871 = n3874 | n3855;
  assign n872 = n871 & n870 & (n869 | n853);
  assign n873 = n840 & n870 & (~n783 | n869);
  assign n874 = (n872 | n995) & (n870 | n891);
  assign n875 = (n873 | n3851) & (n869 | n1056);
  assign n876 = n874 & n875;
  assign n877 = n868 & n876;
  assign n878 = (n877 | n3850) & (n857 | n896);
  assign n879 = n860 & n878 & (n851 | n847);
  assign n880 = n849 & n879 & (n18 | n857);
  assign n881 = n916 & ~Ni41;
  assign n882 = n678 & n814 & (n881 | ~Ni38);
  assign n883 = ~n762 & ~Ni41;
  assign n884 = n814 & n831 & (n883 | ~Ni38);
  assign n885 = n883 & n814;
  assign n886 = Ni32 | ~Ni36;
  assign n887 = Ni32 | Ni36;
  assign n888 = (n885 | n886) & (n884 | n887);
  assign n889 = ~n764 & ~Ni41;
  assign n890 = n814 & n840 & (n889 | ~Ni38);
  assign n891 = ~Ni32 | ~Ni36;
  assign n892 = (n889 | n891) & (~Ni32 | n890);
  assign n893 = ~n3850 & (~n888 | ~n892);
  assign n894 = (n881 | n847) & (n1082 | n2438);
  assign n895 = (~Ni36 | n881) & n882;
  assign n896 = ~n18 | n2420;
  assign n897 = ~n893 & n894 & (n895 | n896);
  assign n898 = n849 & n897 & (n18 | n895);
  assign n899 = Pi22 | ~Ni30;
  assign n900 = n899 & (Pi22 | ~n801);
  assign n901 = n900 & (Pi22 | n18);
  assign n902 = Pi21 | ~Ni30;
  assign n903 = n902 & (Ni31 | Pi21);
  assign n904 = n2421 & n903;
  assign n905 = n904 & (Pi21 | n18);
  assign n906 = Pi21 & ~Pi20;
  assign n907 = ~n844 & n906;
  assign n908 = Pi20 & Pi21;
  assign n909 = ~Pi22 & (n907 | (~n876 & n908));
  assign n910 = n901 & (Pi22 | n892);
  assign n911 = n905 & n910 & (Pi21 | n888);
  assign n912 = (n911 & (Pi19 | ~n3863)) | (~Pi19 & ~n3863);
  assign n913 = (n898 | n1702) & (n850 | n1408);
  assign n914 = Pi19 | n3859;
  assign n915 = n912 & n913 & (n880 | n914);
  assign n916 = n738 & ~Ni42;
  assign n917 = n916 & (Ni40 | n1134);
  assign n918 = n814 & (~Ni37 | n917);
  assign n919 = n678 & (n917 | n817);
  assign n920 = n678 & n918 & (~n783 | n917);
  assign n921 = (n917 | n698) & (n920 | n2434);
  assign n922 = n918 & n921 & (Ni35 | n919);
  assign n923 = Ni43 | Ni42;
  assign n924 = ~n762 & (n1137 | Ni40);
  assign n925 = n814 & (~Ni37 | n924);
  assign n926 = n829 & n925 & (n924 | n817);
  assign n927 = n831 & n925 & (~n783 | n924);
  assign n928 = (n924 | n1052) & (n925 | n886);
  assign n929 = (n927 | n3856) & (n926 | n992);
  assign n930 = n928 & n929;
  assign n931 = ~n764 & (n1140 | Ni40);
  assign n932 = n814 & (~Ni37 | n931);
  assign n933 = n838 & n932 & (n931 | n817);
  assign n934 = n840 & n932 & (~n783 | n931);
  assign n935 = (n933 | n995) & (n932 | n891);
  assign n936_1 = (n934 | n3851) & (n931 | n1056);
  assign n937 = n935 & n936_1;
  assign n938 = n930 & n937;
  assign n939 = (n938 | n3850) & (n922 | n896);
  assign n940 = n826 & n939 & (n917 | n847);
  assign n941 = n849 & n940 & (n18 | n922);
  assign n942 = n916 & (Ni40 | n1148);
  assign n943 = n814 & (~Ni37 | n942);
  assign n944 = n678 & (n942 | n853);
  assign n945 = n678 & n943 & (~n783 | n942);
  assign n946 = (n942 | n698) & (n945 | n2434);
  assign n947 = n943 & n946 & (Ni35 | n944);
  assign n948 = ~n762 & (n1151 | Ni40);
  assign n949 = n814 & (~Ni37 | n948);
  assign n950 = n863 & n949 & (n948 | n853);
  assign n951 = n831 & n949 & (~n783 | n948);
  assign n952 = (n948 | n1052) & (n949 | n886);
  assign n953 = (n951 | n3856) & (n950 | n992);
  assign n954 = n952 & n953;
  assign n955 = ~n764 & (n1154 | Ni40);
  assign n956 = n814 & (~Ni37 | n955);
  assign n957 = n871 & n956 & (n955 | n853);
  assign n958 = n840 & n956 & (~n783 | n955);
  assign n959 = (n957 | n995) & (n956 | n891);
  assign n960 = (n958 | n3851) & (n955 | n1056);
  assign n961 = n959 & n960;
  assign n962 = n954 & n961;
  assign n963 = (n962 | n3850) & (n947 | n896);
  assign n964 = n860 & n963 & (n942 | n847);
  assign n965 = n849 & n964 & (n18 | n947);
  assign n966 = n678 & n814 & (n916 | ~Ni38);
  assign n967 = n814 & n831 & (~n762 | ~Ni38);
  assign n968 = ~n762 & n814;
  assign n969 = (n968 | n886) & (n967 | n887);
  assign n970 = n814 & n840 & (~n764 | ~Ni38);
  assign n971_1 = (~Ni32 | n970) & (~n764 | n891);
  assign n972 = ~n3850 & (~n969 | ~n971_1);
  assign n973 = (n916 | n847) & (n1082 | n2438);
  assign n974 = (~Ni36 | n916) & n966;
  assign n975 = ~n972 & n973 & (n896 | n974);
  assign n976 = n849 & n975 & (n18 | n974);
  assign n977 = n906 & ~n937;
  assign n978 = ~Pi22 & (n977 | (n908 & ~n961));
  assign n979 = n901 & (Pi22 | n971_1);
  assign n980 = n905 & n979 & (Pi21 | n969);
  assign n981 = (n980 & (Pi19 | ~n3880)) | (~Pi19 & ~n3880);
  assign n982 = (n976 | n1702) & (n941 | n1408);
  assign n983 = n981 & n982 & (n965 | n914);
  assign n984 = n819 & (Ni35 | n818);
  assign n985 = Ni38 | n676;
  assign n986_1 = ~Ni37 & ~Ni38;
  assign n987 = n985 & n986_1;
  assign n988 = n987 | n1083;
  assign n989 = n987 & n822;
  assign n990 = n988 & (n989 | n825);
  assign n991 = Ni32 | ~n2530;
  assign n992 = Ni32 | Ni35;
  assign n993 = (n832 | n991) & (n830 | n992);
  assign n994 = n1241 & n891;
  assign n995 = ~Ni32 | Ni35;
  assign n996 = (n841 | n994) & (n839 | n995);
  assign n997 = n993 & n996;
  assign n998 = (n997 | n3850) & (n984 | n896);
  assign n999 = n990 & n998 & (n815 | n847);
  assign n1000 = n849 & n999 & (n18 | n984);
  assign n1001_1 = n855 & (Ni35 | n854);
  assign n1002 = n987 & n858;
  assign n1003 = n988 & (n1002 | n825);
  assign n1004 = (n865 | n991) & (n864 | n992);
  assign n1005 = (n873 | n994) & (n872 | n995);
  assign n1006 = n1004 & n1005;
  assign n1007 = (n1006 | n3850) & (n1001_1 | n896);
  assign n1008 = n1003 & n1007 & (n851 | n847);
  assign n1009 = n849 & n1008 & (n18 | n1001_1);
  assign n1010 = n4071 & (n890 | n3663);
  assign n1011 = (n881 | n847) & (n987 | n2438);
  assign n1012 = n1010 & n1011 & (n882 | n896);
  assign n1013 = n849 & n1012 & (n18 | n882);
  assign n1014 = n906 & ~n996;
  assign n1015 = ~Pi22 & (n1014 | (n908 & ~n1005));
  assign n1016 = n901 & (Pi22 | n890);
  assign n1017 = n905 & n1016 & (Pi21 | n884);
  assign n1018 = (n1017 & (Pi19 | ~n3873)) | (~Pi19 & ~n3873);
  assign n1019 = (n1013 | n1702) & (n1000 | n1408);
  assign n1020 = n1018 & n1019 & (n1009 | n914);
  assign n1021_1 = n920 & (Ni35 | n919);
  assign n1022 = (n927 | n991) & (n926 | n992);
  assign n1023 = (n934 | n994) & (n933 | n995);
  assign n1024 = n1022 & n1023;
  assign n1025 = (n1024 | n3850) & (n1021_1 | n896);
  assign n1026 = n990 & n1025 & (n917 | n847);
  assign n1027 = n849 & n1026 & (n18 | n1021_1);
  assign n1028 = n945 & (Ni35 | n944);
  assign n1029 = (n951 | n991) & (n950 | n992);
  assign n1030 = (n958 | n994) & (n957 | n995);
  assign n1031 = n1029 & n1030;
  assign n1032 = (n1031 | n3850) & (n1028 | n896);
  assign n1033 = n1003 & n1032 & (n942 | n847);
  assign n1034 = n849 & n1033 & (n18 | n1028);
  assign n1035 = n4072 & (n970 | n3663);
  assign n1036_1 = (n916 | n847) & (n987 | n2438);
  assign n1037 = n1035 & n1036_1 & (n966 | n896);
  assign n1038 = n849 & n1037 & (n18 | n966);
  assign n1039 = n906 & ~n1023;
  assign n1040 = ~Pi22 & (n1039 | (n908 & ~n1030));
  assign n1041 = n901 & (Pi22 | n970);
  assign n1042 = n905 & n1041 & (Pi21 | n967);
  assign n1043 = (n1042 & (Pi19 | ~n3887)) | (~Pi19 & ~n3887);
  assign n1044 = (n1038 | n1702) & (n1027 | n1408);
  assign n1045 = n1043 & n1044 & (n1034 | n914);
  assign n1046 = n1048 | (~Ni37 & n817);
  assign n1047 = n1046 & n814 & n678;
  assign n1048 = ~n674 & ~n2426;
  assign n1049 = n1047 & (n1048 | n698);
  assign n1050 = ~Ni32 & (~n814 | ~n829 | ~n4056);
  assign n1051_1 = ~n763 & ~Ni41;
  assign n1052 = Ni32 | n698;
  assign n1053 = ~n1050 & (n1051_1 | n1052);
  assign n1054 = Ni32 & (~n814 | ~n838 | ~n4055);
  assign n1055 = ~n765 & ~Ni41;
  assign n1056 = Ni37 | n891;
  assign n1057 = ~n1054 & (n1055 | n1056);
  assign n1058 = ~n3850 & (~n1053 | ~n1057);
  assign n1059 = (n1048 | n847) & (n824 | n2438);
  assign n1060 = ~n1058 & (n896 | n1049) & n1059;
  assign n1061_1 = n849 & n1060 & (n18 | n1049);
  assign n1062 = n1064 | (~Ni37 & n853);
  assign n1063 = n1062 & n814 & n678;
  assign n1064 = ~n675 & ~n2426;
  assign n1065 = n1063 & (n1064 | n698);
  assign n1066 = ~Ni32 & (~n814 | ~n863 | ~n4058);
  assign n1067 = ~n766 & ~Ni41;
  assign n1068 = ~n1066 & (n1052 | n1067);
  assign n1069 = Ni32 & (~n814 | ~n871 | ~n4057);
  assign n1070 = ~n767 & ~Ni41;
  assign n1071 = ~n1069 & (n1056 | n1070);
  assign n1072 = ~n3850 & (~n1068 | ~n1071);
  assign n1073 = (n1064 | n847) & (n859 | n2438);
  assign n1074 = ~n1072 & (n896 | n1065) & n1073;
  assign n1075 = n849 & n1074 & (n18 | n1065);
  assign n1076_1 = n881 & (n1048 | ~Ni40);
  assign n1077 = n814 & (~Ni37 | n1076_1);
  assign n1078 = n678 & n1077 & (~n783 | n1076_1);
  assign n1079 = n678 & (n1076_1 | n817);
  assign n1080 = (n1076_1 | n698) & (n1078 | n2530);
  assign n1081_1 = n1077 & n1080 & (~Ni35 | n1079);
  assign n1082 = ~Ni36 & n987;
  assign n1083 = ~Ni35 | n2438;
  assign n1084 = (n1082 | n825) & (n824 | n1083);
  assign n1085_1 = n883 & (n1051_1 | ~Ni40);
  assign n1086 = n814 & (~Ni37 | n1085_1);
  assign n1087 = n831 & n1086 & (~n783 | n1085_1);
  assign n1088 = n829 & n1086 & (n1085_1 | n817);
  assign n1089 = (n1085_1 | n1052) & (n1086 | n886);
  assign n1090 = (n1087 | n3869) & (n1088 | n1238);
  assign n1091 = n1089 & n1090;
  assign n1092 = n889 & (n1055 | ~Ni40);
  assign n1093 = n814 & (~Ni37 | n1092);
  assign n1094 = n840 & n1093 & (~n783 | n1092);
  assign n1095 = n838 & n1093 & (n1092 | n817);
  assign n1096 = (n1095 | n1241) & (n1093 | n891);
  assign n1097 = (n1094 | n3868) & (n1092 | n1056);
  assign n1098 = n1096 & n1097;
  assign n1099 = n1091 & n1098;
  assign n1100 = (n1099 | n3850) & (n1081_1 | n896);
  assign n1101 = n1084 & n1100 & (n1076_1 | n847);
  assign n1102 = n849 & n1101 & (n18 | n1081_1);
  assign n1103 = n881 & (n1064 | ~Ni40);
  assign n1104 = n814 & (~Ni37 | n1103);
  assign n1105 = n678 & n1104 & (~n783 | n1103);
  assign n1106 = n678 & (n1103 | n853);
  assign n1107 = (n1103 | n698) & (n1105 | n2530);
  assign n1108 = n1104 & n1107 & (~Ni35 | n1106);
  assign n1109 = (n1082 | n825) & (n859 | n1083);
  assign n1110 = n883 & (n1067 | ~Ni40);
  assign n1111 = n814 & (~Ni37 | n1110);
  assign n1112 = n831 & n1111 & (~n783 | n1110);
  assign n1113 = n863 & n1111 & (n1110 | n853);
  assign n1114 = (n1110 | n1052) & (n1111 | n886);
  assign n1115 = (n1112 | n3869) & (n1113 | n1238);
  assign n1116 = n1114 & n1115;
  assign n1117 = n889 & (n1070 | ~Ni40);
  assign n1118 = n814 & (~Ni37 | n1117);
  assign n1119 = n840 & n1118 & (~n783 | n1117);
  assign n1120 = n871 & n1118 & (n1117 | n853);
  assign n1121 = (n1120 | n1241) & (n1118 | n891);
  assign n1122 = (n1119 | n3868) & (n1117 | n1056);
  assign n1123 = n1121 & n1122;
  assign n1124 = n1116 & n1123;
  assign n1125 = (n1124 | n3850) & (n1108 | n896);
  assign n1126 = n1109 & n1125 & (n1103 | n847);
  assign n1127 = n849 & n1126 & (n18 | n1108);
  assign n1128 = n906 & ~n1098;
  assign n1129 = ~Pi22 & (n1128 | (n908 & ~n1123));
  assign n1130 = n906 & ~n1057;
  assign n1131 = ~Pi22 & (n1130 | (n908 & ~n1071));
  assign n1132 = n1134 | (~Ni37 & n817);
  assign n1133 = n1132 & n814 & n678;
  assign n1134 = n4769 & n916;
  assign n1135 = n1133 & (n1134 | n698);
  assign n1136 = ~Ni32 & (~n814 | ~n829 | ~n4062);
  assign n1137 = ~n762 & ~n763;
  assign n1138 = ~n1136 & (n1052 | n1137);
  assign n1139 = Ni32 & (~n814 | ~n838 | ~n4061);
  assign n1140 = ~n764 & ~n765;
  assign n1141 = ~n1139 & (n1056 | n1140);
  assign n1142 = ~n3850 & (~n1138 | ~n1141);
  assign n1143 = (n1134 | n847) & (n824 | n2438);
  assign n1144 = ~n1142 & (n896 | n1135) & n1143;
  assign n1145 = n849 & n1144 & (n18 | n1135);
  assign n1146 = n1148 | (~Ni37 & n853);
  assign n1147 = n1146 & n814 & n678;
  assign n1148 = n4770 & n916;
  assign n1149 = n1147 & (n1148 | n698);
  assign n1150 = ~Ni32 & (~n814 | ~n863 | ~n4064);
  assign n1151 = ~n762 & ~n766;
  assign n1152 = ~n1150 & (n1052 | n1151);
  assign n1153 = Ni32 & (~n814 | ~n871 | ~n4063);
  assign n1154 = ~n764 & ~n767;
  assign n1155 = ~n1153 & (n1056 | n1154);
  assign n1156 = ~n3850 & (~n1152 | ~n1155);
  assign n1157 = (n1148 | n847) & (n859 | n2438);
  assign n1158 = ~n1156 & (n896 | n1149) & n1157;
  assign n1159 = n849 & n1158 & (n18 | n1149);
  assign n1160 = n916 & (n1134 | ~Ni40);
  assign n1161 = n814 & (~Ni37 | n1160);
  assign n1162 = n678 & n1161 & (~n783 | n1160);
  assign n1163 = n678 & (n1160 | n817);
  assign n1164 = (n1160 | n698) & (n1162 | n2530);
  assign n1165 = n1161 & n1164 & (~Ni35 | n1163);
  assign n1166 = ~n762 & (n1137 | ~Ni40);
  assign n1167 = n814 & (~Ni37 | n1166);
  assign n1168 = n831 & n1167 & (~n783 | n1166);
  assign n1169 = n829 & n1167 & (n1166 | n817);
  assign n1170 = (n1166 | n1052) & (n1167 | n886);
  assign n1171 = (n1168 | n3869) & (n1169 | n1238);
  assign n1172 = n1170 & n1171;
  assign n1173 = ~n764 & (n1140 | ~Ni40);
  assign n1174 = n814 & (~Ni37 | n1173);
  assign n1175 = n840 & n1174 & (~n783 | n1173);
  assign n1176 = n838 & n1174 & (n1173 | n817);
  assign n1177 = (n1176 | n1241) & (n1174 | n891);
  assign n1178 = (n1175 | n3868) & (n1173 | n1056);
  assign n1179 = n1177 & n1178;
  assign n1180 = n1172 & n1179;
  assign n1181 = (n1180 | n3850) & (n1165 | n896);
  assign n1182 = n1084 & n1181 & (n1160 | n847);
  assign n1183 = n849 & n1182 & (n18 | n1165);
  assign n1184 = n916 & (n1148 | ~Ni40);
  assign n1185 = n814 & (~Ni37 | n1184);
  assign n1186 = n678 & n1185 & (~n783 | n1184);
  assign n1187 = n678 & (n1184 | n853);
  assign n1188 = (n1184 | n698) & (n1186 | n2530);
  assign n1189 = n1185 & n1188 & (~Ni35 | n1187);
  assign n1190 = ~n762 & (n1151 | ~Ni40);
  assign n1191 = n814 & (~Ni37 | n1190);
  assign n1192 = n831 & n1191 & (~n783 | n1190);
  assign n1193 = n863 & n1191 & (n1190 | n853);
  assign n1194 = (n1190 | n1052) & (n1191 | n886);
  assign n1195 = (n1192 | n3869) & (n1193 | n1238);
  assign n1196 = n1194 & n1195;
  assign n1197 = ~n764 & (n1154 | ~Ni40);
  assign n1198 = n814 & (~Ni37 | n1197);
  assign n1199 = n840 & n1198 & (~n783 | n1197);
  assign n1200 = n871 & n1198 & (n1197 | n853);
  assign n1201 = (n1200 | n1241) & (n1198 | n891);
  assign n1202 = (n1199 | n3868) & (n1197 | n1056);
  assign n1203 = n1201 & n1202;
  assign n1204 = n1196 & n1203;
  assign n1205 = (n1204 | n3850) & (n1189 | n896);
  assign n1206 = n1109 & n1205 & (n1184 | n847);
  assign n1207 = n849 & n1206 & (n18 | n1189);
  assign n1208 = n906 & ~n1179;
  assign n1209 = ~Pi22 & (n1208 | (n908 & ~n1203));
  assign n1210 = n906 & ~n1141;
  assign n1211 = ~Pi22 & (n1210 | (n908 & ~n1155));
  assign n1212 = (n914 | n1159) & (Pi19 | ~n3883);
  assign n1213 = (n1183 | n3893) & (n1207 | n2109);
  assign n1214 = n1145 | n1408;
  assign n1215 = ~n3789 & n1214 & n1212 & n1213;
  assign n1216 = n698 | ~Ni38;
  assign n1217 = n1047 & (n1048 | n1216);
  assign n1218 = n831 | n1052;
  assign n1219 = Ni32 | n1216;
  assign n1220 = ~n1050 & n1218 & (n1051_1 | n1219);
  assign n1221 = n891 | n840;
  assign n1222 = ~n783 | n891;
  assign n1223 = ~n1054 & n1221 & (n1055 | n1222);
  assign n1224 = ~n3850 & (~n1220 | ~n1223);
  assign n1225 = (n1048 | n847) & (n989 | n2438);
  assign n1226 = ~n1224 & (n896 | n1217) & n1225;
  assign n1227 = n849 & n1226 & (n18 | n1217);
  assign n1228 = n1063 & (n1064 | n1216);
  assign n1229 = ~n1066 & n1218 & (n1067 | n1219);
  assign n1230 = ~n1069 & n1221 & (n1070 | n1222);
  assign n1231 = ~n3850 & (~n1229 | ~n1230);
  assign n1232 = (n1064 | n847) & (n1002 | n2438);
  assign n1233 = ~n1231 & (n896 | n1228) & n1232;
  assign n1234 = n849 & n1233 & (n18 | n1228);
  assign n1235 = n1078 & (~Ni35 | n1079);
  assign n1236 = (n987 | n825) & (n989 | n1083);
  assign n1237 = Ni32 | ~n2434;
  assign n1238 = Ni32 | ~Ni35;
  assign n1239 = (n1087 | n1237) & (n1088 | n1238);
  assign n1240 = n995 & n891;
  assign n1241 = ~Ni32 | ~Ni35;
  assign n1242 = (n1094 | n1240) & (n1095 | n1241);
  assign n1243 = n1239 & n1242;
  assign n1244 = (n1243 | n3850) & (n1235 | n896);
  assign n1245 = n1236 & n1244 & (n1076_1 | n847);
  assign n1246 = n849 & n1245 & (n18 | n1235);
  assign n1247 = n1105 & (~Ni35 | n1106);
  assign n1248 = (n987 | n825) & (n1002 | n1083);
  assign n1249 = (n1112 | n1237) & (n1113 | n1238);
  assign n1250 = (n1119 | n1240) & (n1120 | n1241);
  assign n1251 = n1249 & n1250;
  assign n1252 = (n1251 | n3850) & (n1247 | n896);
  assign n1253 = n1248 & n1252 & (n1103 | n847);
  assign n1254 = n849 & n1253 & (n18 | n1247);
  assign n1255 = n906 & ~n1242;
  assign n1256 = ~Pi22 & (n1255 | (n908 & ~n1250));
  assign n1257 = n906 & ~n1223;
  assign n1258 = ~Pi22 & (n1257 | (n908 & ~n1230));
  assign n1259 = n1133 & (n1134 | n1216);
  assign n1260 = ~n1136 & n1218 & (n1137 | n1219);
  assign n1261 = ~n1139 & n1221 & (n1140 | n1222);
  assign n1262 = ~n3850 & (~n1260 | ~n1261);
  assign n1263 = (n1134 | n847) & (n989 | n2438);
  assign n1264 = ~n1262 & (n896 | n1259) & n1263;
  assign n1265 = n849 & n1264 & (n18 | n1259);
  assign n1266 = n1147 & (n1148 | n1216);
  assign n1267 = ~n1150 & n1218 & (n1151 | n1219);
  assign n1268 = ~n1153 & n1221 & (n1154 | n1222);
  assign n1269 = ~n3850 & (~n1267 | ~n1268);
  assign n1270 = (n1148 | n847) & (n1002 | n2438);
  assign n1271 = ~n1269 & (n896 | n1266) & n1270;
  assign n1272 = n849 & n1271 & (n18 | n1266);
  assign n1273 = n1162 & (~Ni35 | n1163);
  assign n1274 = (n1168 | n1237) & (n1169 | n1238);
  assign n1275 = (n1175 | n1240) & (n1176 | n1241);
  assign n1276 = n1274 & n1275;
  assign n1277 = (n1276 | n3850) & (n1273 | n896);
  assign n1278 = n1236 & n1277 & (n1160 | n847);
  assign n1279 = n849 & n1278 & (n18 | n1273);
  assign n1280 = n1186 & (~Ni35 | n1187);
  assign n1281 = (n1192 | n1237) & (n1193 | n1238);
  assign n1282 = (n1199 | n1240) & (n1200 | n1241);
  assign n1283 = n1281 & n1282;
  assign n1284 = (n1283 | n3850) & (n1280 | n896);
  assign n1285 = n1248 & n1284 & (n1184 | n847);
  assign n1286 = n849 & n1285 & (n18 | n1280);
  assign n1287 = n906 & ~n1275;
  assign n1288 = ~Pi22 & (n1287 | (n908 & ~n1282));
  assign n1289 = n906 & ~n1261;
  assign n1290 = ~Pi22 & (n1289 | (n908 & ~n1268));
  assign n1291 = (n914 | n1272) & (Pi19 | ~n3890);
  assign n1292 = (n1279 | n3893) & (n1286 | n2109);
  assign n1293 = n1265 | n1408;
  assign n1294 = ~n3792 & n1293 & n1291 & n1292;
  assign n1295 = ~n901 | n1129 | n3783 | n3784;
  assign n1296 = ~n3870 & (n1295 | ~n4084 | ~n4085);
  assign n1297 = ~n901 | n1256 | n3785 | n3786;
  assign n1298 = ~n3877 & (n1297 | ~n4087 | ~n4088);
  assign n1299 = ~n901 | n1258 | n3875 | n3876;
  assign n1300 = ~n2272 & (n1299 | ~n4075);
  assign n1301 = n18 & (n3737 | (~n3792 & n4078));
  assign n1302 = n4082 & (n3743 | (~n3890 & n4077));
  assign n1303 = n4081 & (n3740 | (~n3887 & n4074));
  assign n1304 = n4079 & (n1012 | n1495);
  assign n1305 = n1304 & n1303 & n1301 & n1302;
  assign n1306 = ~n901 | n1131 | n3865 | n3866;
  assign n1307 = ~n2272 & (n1306 | ~n4059);
  assign n1308 = n18 & (n3737 | (~n3789 & n4066));
  assign n1309 = n4070 & (n3743 | (~n3883 & n4065));
  assign n1310 = n4069 & (n3740 | (~n3880 & n4054));
  assign n1311 = n4067 & (n897 | n1495);
  assign n1312 = n1311 & n1310 & n1308 & n1309;
  assign n1313 = n4103 & (n1183 | n2372);
  assign n1314 = ~Pi25 | n3859;
  assign n1315 = n1313 & ~n3789 & (n1207 | n1314);
  assign n1316 = n4102 & (n1145 | n2372);
  assign n1317 = n1316 & (n1159 | n1314) & ~n3883;
  assign n1318 = n4101 & (n941 | n2372);
  assign n1319 = n1318 & (n965 | n1314) & ~n3880;
  assign n1320 = (n1319 | n3864) & (n1317 | n3867);
  assign n1321 = n4096 & n4104 & (n975 | n3848);
  assign n1322 = ~Pi19 | Pi17;
  assign n1323 = n1320 & n1321 & (n1315 | n1322);
  assign n1324 = n4094 & (n1102 | n2372);
  assign n1325 = ~n1295 & n1324 & (n1127 | n1314);
  assign n1326 = n4093 & (n1061_1 | n2372);
  assign n1327 = ~n1306 & n1326 & (n1075 | n1314);
  assign n1328 = n4092 & (n850 | n2372);
  assign n1329 = n1328 & (n880 | n1314) & ~n3863;
  assign n1330 = (n1329 | n3864) & (n1327 | n3867);
  assign n1331 = n4096 & n4095 & (n897 | n3848);
  assign n1332 = n1330 & n1331 & (n1325 | n1322);
  assign n1333 = n4107 & (n1279 | n2372);
  assign n1334 = n1333 & (n1286 | n1314) & ~n3792;
  assign n1335 = n4106 & (n1265 | n2372);
  assign n1336 = n1335 & (n1272 | n1314) & ~n3890;
  assign n1337 = n4105 & (n1027 | n2372);
  assign n1338 = n1337 & (n1034 | n1314) & ~n3887;
  assign n1339 = (n1338 | n3864) & (n1336 | n3867);
  assign n1340 = n4096 & n4108 & (n1037 | n3848);
  assign n1341 = n1339 & n1340 & (n1334 | n1322);
  assign n1342 = n4099 & (n1246 | n2372);
  assign n1343 = ~n1297 & n1342 & (n1254 | n1314);
  assign n1344 = n4098 & (n1227 | n2372);
  assign n1345 = ~n1299 & n1344 & (n1234 | n1314);
  assign n1346 = n4097 & (n1000 | n2372);
  assign n1347 = n1346 & (n1009 | n1314) & ~n3873;
  assign n1348 = (n1347 | n3864) & (n1345 | n3867);
  assign n1349 = n4096 & n4100 & (n1012 | n3848);
  assign n1350 = n1348 & n1349 & (n1343 | n1322);
  assign n1351 = n738 & Ni42;
  assign n1352 = n985 & (~n814 | n1351);
  assign n1353 = ~Ni31 | ~Ni30;
  assign n1354 = (~Ni30 | Ni33) & n1353;
  assign n1355 = ~n18 | ~Ni30;
  assign n1356 = ~n707 & ~Ni30;
  assign n1357 = n1355 & (n18 | n1356);
  assign n1358 = ~n711 & ~Ni30;
  assign n1359 = n1355 & (n18 | n1358);
  assign n1360 = ~n714 & ~Ni30;
  assign n1361 = n1355 & (n18 | n1360);
  assign n1362 = n899 & n902;
  assign n1363 = (n1534 | n1702) & (n4135 | n1408);
  assign n1364 = n1520 & n1359;
  assign n1365 = n1362 & n1363 & (n1364 | n914);
  assign n1366 = ~n732 & ~Ni30;
  assign n1367 = n1355 & (n18 | n1366);
  assign n1368 = ~n736 & ~Ni30;
  assign n1369 = n1355 & (n18 | n1368);
  assign n1370 = ~n739 & ~Ni30;
  assign n1371 = n1355 & (n18 | n1370);
  assign n1372 = (n1535 | n1702) & (n4136 | n1408);
  assign n1373 = n1532 & n1369;
  assign n1374 = n1362 & n1372 & (n1373 | n914);
  assign n1375 = ~n749 & ~Ni30;
  assign n1376 = n1355 & (n18 | n1375);
  assign n1377 = ~n751 & ~Ni30;
  assign n1378 = n1355 & (n18 | n1377);
  assign n1379 = ~Ni30 & n1465;
  assign n1380 = n1355 & (n18 | n1379);
  assign n1381 = (n1494 | n1702) & (n4149 | n1408);
  assign n1382 = n1480 & n1378;
  assign n1383 = n1362 & n1381 & (n1382 | n914);
  assign n1384 = ~n759 & ~Ni30;
  assign n1385 = n1355 & (n18 | n1384);
  assign n1386 = ~n761 & ~Ni30;
  assign n1387 = n1355 & (n18 | n1386);
  assign n1388 = ~Ni30 & n1468;
  assign n1389 = n1355 & (n18 | n1388);
  assign n1390 = (n1496 | n1702) & (n4150 | n1408);
  assign n1391 = n1492 & n1387;
  assign n1392 = n1362 & n1390 & (n1391 | n914);
  assign n1393 = ~Ni37 | n985;
  assign n1394 = n676 | n3853;
  assign n1395 = n3959 & n3183;
  assign n1396 = ~n691 & ~Ni30;
  assign n1397 = n1355 & (n18 | n1396);
  assign n1398 = n3961 & n3183;
  assign n1399 = ~n694 & ~Ni30;
  assign n1400 = n1355 & (n18 | n1399);
  assign n1401 = ~n699 & ~Ni30;
  assign n1402 = n1355 & (n18 | n1401);
  assign n1403 = ~n703 & ~Ni30;
  assign n1404 = n1355 & (n18 | n1403);
  assign n1405 = (n4140 | n3893) & (n4141 | n2109);
  assign n1406 = n1362 & (n4138 | n914);
  assign n1407 = n1514 & n1397;
  assign n1408 = Pi19 | n3857;
  assign n1409 = n1405 & n1406 & (n1407 | n1408);
  assign n1410 = ~n717 & ~Ni30;
  assign n1411 = n1355 & (n18 | n1410);
  assign n1412 = ~n720 & ~Ni30;
  assign n1413 = n1355 & (n18 | n1412);
  assign n1414 = ~n724 & ~Ni30;
  assign n1415 = n1355 & (n18 | n1414);
  assign n1416 = ~n728 & ~Ni30;
  assign n1417 = n1355 & (n18 | n1416);
  assign n1418 = (n4145 | n3893) & (n4146 | n2109);
  assign n1419 = n1362 & (n4143 | n914);
  assign n1420 = n1526 & n1411;
  assign n1421 = n1418 & n1419 & (n1420 | n1408);
  assign n1422 = ~n742 & ~Ni30;
  assign n1423 = n1355 & (n18 | n1422);
  assign n1424 = ~n743 & ~Ni30;
  assign n1425 = n1355 & (n18 | n1424);
  assign n1426 = ~n745 & ~Ni30;
  assign n1427 = n1355 & (n18 | n1426);
  assign n1428 = ~n747 & ~Ni30;
  assign n1429 = n1355 & (n18 | n1428);
  assign n1430 = (n4154 | n3893) & (n4155 | n2109);
  assign n1431 = n1362 & (n4152 | n914);
  assign n1432 = n1474 & n1423;
  assign n1433 = n1430 & n1431 & (n1432 | n1408);
  assign n1434 = ~n752 & ~Ni30;
  assign n1435 = n1355 & (n18 | n1434);
  assign n1436 = ~n753 & ~Ni30;
  assign n1437 = n1355 & (n18 | n1436);
  assign n1438 = ~n755 & ~Ni30;
  assign n1439 = n1355 & (n18 | n1438);
  assign n1440 = ~n757 & ~Ni30;
  assign n1441 = n1355 & (n18 | n1440);
  assign n1442 = (n4159 | n3893) & (n4160 | n2109);
  assign n1443 = n1362 & (n4157 | n914);
  assign n1444 = n1486 & n1435;
  assign n1445 = n1442 & n1443 & (n1444 | n1408);
  assign n1446 = Ni12 | n2750;
  assign n1447 = n1461 & n1362;
  assign n1448 = Ni12 | ~n2750;
  assign n1449 = (n1447 | n1448) & (n1446 | ~n3991);
  assign n1450 = ~n3696 & (~n1552 | (~n1986 & ~n2254));
  assign n1451 = ~n1450 & (n2632 | (~n3918 & n4300));
  assign n1452 = ~Ni12 | ~Ni13;
  assign n1453 = n1449 & n1451 & (n1447 | n1452);
  assign n1454 = n1354 & (~Ni30 | ~n3761);
  assign n1455 = n1454 | (Pi22 & Pi21);
  assign n1456 = n1455 | n3677;
  assign n1457 = (n1541 | n1610) & (n1447 | ~n3898);
  assign n1458 = n1456 & n1457 & (Ni11 | n1453);
  assign n1459 = n4772 | n2254;
  assign n1460 = (Pi24 | n1362) & (~n793 | n1463);
  assign n1461 = n1918 | n2254;
  assign n1462 = n1459 & n1460 & (Pi24 | n1461);
  assign n1463 = n1353 & n3795;
  assign n1464 = n4766 | n1465;
  assign n1465 = ~n712 | n1539;
  assign n1466 = n1463 & n1464 & (n18 | n1465);
  assign n1467 = n4766 | n1468;
  assign n1468 = ~n737 | n1539;
  assign n1469 = n1463 & n1467 & (n18 | n1468);
  assign n1470 = ~n745 | n4766;
  assign n1471 = n1463 & n1470 & (n18 | ~n745);
  assign n1472 = ~n747 | n4766;
  assign n1473 = n1463 & n1472 & (n18 | ~n747);
  assign n1474 = ~n742 | n4766;
  assign n1475 = n1463 & n1474 & (n18 | ~n742);
  assign n1476 = ~n743 | n4766;
  assign n1477 = n1463 & n1476 & (n18 | ~n743);
  assign n1478 = ~n749 | n4766;
  assign n1479 = n1463 & n1478 & (n18 | ~n749);
  assign n1480 = ~n751 | n4766;
  assign n1481 = n1463 & n1480 & (n18 | ~n751);
  assign n1482 = ~n755 | n4766;
  assign n1483 = n1463 & n1482 & (n18 | ~n755);
  assign n1484 = ~n757 | n4766;
  assign n1485 = n1463 & n1484 & (n18 | ~n757);
  assign n1486 = ~n752 | n4766;
  assign n1487 = n1463 & n1486 & (n18 | ~n752);
  assign n1488 = ~n753 | n4766;
  assign n1489 = n1463 & n1488 & (n18 | ~n753);
  assign n1490 = ~n759 | n4766;
  assign n1491 = n1463 & n1490 & (n18 | ~n759);
  assign n1492 = ~n761 | n4766;
  assign n1493 = n1463 & n1492 & (n18 | ~n761);
  assign n1494 = n1464 & n1380;
  assign n1495 = Pi16 | n3848;
  assign n1496 = n1467 & n1389;
  assign n1497 = ~Pi16 | n3848;
  assign n1498 = (n1494 | n1495) & (n1496 | n1497);
  assign n1499 = ~n3894 & (~n4277 | ~n4278);
  assign n1500 = ~n2272 & (~n4281 | ~n4282);
  assign n1501 = n1460 & (n3737 | (n4288 & n4287));
  assign n1502 = n4290 & (n3743 | (n4286 & n4285));
  assign n1503 = ~n1499 & (n3740 | (n4279 & n4280));
  assign n1504 = n4289 & (Pi24 | n1498);
  assign n1505 = n1504 & n1503 & n1501 & n1502;
  assign n1506 = ~n714 | n4766;
  assign n1507 = n1463 & n1506 & (n18 | ~n714);
  assign n1508 = ~n739 | n4766;
  assign n1509 = n1463 & n1508 & (n18 | ~n739);
  assign n1510 = ~n699 | n4766;
  assign n1511 = n1463 & n1510 & (n18 | ~n699);
  assign n1512 = ~n703 | n4766;
  assign n1513 = n1463 & n1512 & (n18 | ~n703);
  assign n1514 = ~n691 | n4766;
  assign n1515 = n1463 & n1514 & (n18 | ~n691);
  assign n1516 = ~n694 | n4766;
  assign n1517 = n1463 & n1516 & (n18 | ~n694);
  assign n1518 = ~n707 | n4766;
  assign n1519 = n1463 & n1518 & (n18 | ~n707);
  assign n1520 = ~n711 | n4766;
  assign n1521 = n1463 & n1520 & (n18 | ~n711);
  assign n1522 = ~n724 | n4766;
  assign n1523 = n1463 & n1522 & (n18 | ~n724);
  assign n1524 = ~n728 | n4766;
  assign n1525 = n1463 & n1524 & (n18 | ~n728);
  assign n1526 = ~n717 | n4766;
  assign n1527 = n1463 & n1526 & (n18 | ~n717);
  assign n1528 = ~n720 | n4766;
  assign n1529 = n1463 & n1528 & (n18 | ~n720);
  assign n1530 = ~n732 | n4766;
  assign n1531 = n1463 & n1530 & (n18 | ~n732);
  assign n1532 = ~n736 | n4766;
  assign n1533 = n1463 & n1532 & (n18 | ~n736);
  assign n1534 = n1506 & n1361;
  assign n1535 = n1508 & n1371;
  assign n1536 = (n1534 | n1495) & (n1535 | n1497);
  assign n1537 = ~n3894 & (~n4259 | ~n4260);
  assign n1538 = ~n2272 & (~n4263 | ~n4264);
  assign n1539 = Ni32 | n2420;
  assign n1540 = ~n1352 | n1539;
  assign n1541 = n3794 & (Pi26 | n1918);
  assign n1542 = ~Ni11 | ~Ni12;
  assign n1543 = Ni12 | Ni11;
  assign n1544 = n1542 & ~Ni13 & (Ni14 | n1543);
  assign n1545 = Ni11 & ~Ni12;
  assign n1546 = ~n1462 & n1545 & (~n1541 | ~Ni14);
  assign n1547 = ~n3928 & ~n4674 & (Ni14 | ~n3993);
  assign n1548 = ~n3944 & (~n4273 | ~n4275 | ~n4276);
  assign n1549 = ~n794 & n1459 & (~n788 | n1461);
  assign n1550 = Pi21 | n3801;
  assign n1551 = Pi22 | n3801;
  assign n1552 = n1550 & n1551;
  assign n1553 = ~Ni13 & (Ni14 | Ni12);
  assign n1554 = ~n794 & (n1523 | n3935);
  assign n1555 = (n4145 | n3936) & (n4146 | n2707);
  assign n1556 = n3859 | n788;
  assign n1557 = n1554 & n1555 & (n1525 | n1556);
  assign n1558 = ~n794 & (n1527 | n3935);
  assign n1559 = (n1420 | n3936) & (n4143 | n2707);
  assign n1560 = n1558 & n1559 & (n1529 | n1556);
  assign n1561 = ~n794 & (n1531 | n3935);
  assign n1562 = (n4136 | n3936) & (n1373 | n2707);
  assign n1563 = n1561 & n1562 & (n1533 | n1556);
  assign n1564 = (n1563 | n3864) & (n1560 | n3867);
  assign n1565 = n4254 & n4252 & (n1535 | n3934);
  assign n1566 = n1564 & n1565 & (n1557 | n1322);
  assign n1567 = ~n794 & (n1511 | n3935);
  assign n1568 = (n4140 | n3936) & (n4141 | n2707);
  assign n1569 = n1567 & n1568 & (n1513 | n1556);
  assign n1570 = ~n794 & (n1515 | n3935);
  assign n1571 = (n1407 | n3936) & (n4138 | n2707);
  assign n1572 = n1570 & n1571 & (n1517 | n1556);
  assign n1573 = ~n794 & (n1519 | n3935);
  assign n1574 = (n4135 | n3936) & (n1364 | n2707);
  assign n1575 = n1573 & n1574 & (n1521 | n1556);
  assign n1576 = (n1575 | n3864) & (n1572 | n3867);
  assign n1577 = n4251 & n4252 & (n1534 | n3934);
  assign n1578 = n1576 & n1577 & (n1569 | n1322);
  assign n1579 = ~n794 & (n1483 | n3935);
  assign n1580 = (n4159 | n3936) & (n4160 | n2707);
  assign n1581 = n1579 & n1580 & (n1485 | n1556);
  assign n1582 = ~n794 & (n1487 | n3935);
  assign n1583 = (n1444 | n3936) & (n4157 | n2707);
  assign n1584 = n1582 & n1583 & (n1489 | n1556);
  assign n1585 = ~n794 & (n1491 | n3935);
  assign n1586 = (n4150 | n3936) & (n1391 | n2707);
  assign n1587 = n1585 & n1586 & (n1493 | n1556);
  assign n1588 = (n1587 | n3864) & (n1584 | n3867);
  assign n1589 = n4255 & n4252 & (n1496 | n3934);
  assign n1590 = n1588 & n1589 & (n1581 | n1322);
  assign n1591 = ~n794 & (n1471 | n3935);
  assign n1592 = (n4154 | n3936) & (n4155 | n2707);
  assign n1593 = n1591 & n1592 & (n1473 | n1556);
  assign n1594 = ~n794 & (n1475 | n3935);
  assign n1595 = (n1432 | n3936) & (n4152 | n2707);
  assign n1596 = n1594 & n1595 & (n1477 | n1556);
  assign n1597 = ~n794 & (n1479 | n3935);
  assign n1598 = (n4149 | n3936) & (n1382 | n2707);
  assign n1599 = n1597 & n1598 & (n1481 | n1556);
  assign n1600 = (n1599 | n3864) & (n1596 | n3867);
  assign n1601 = n4253 & n4252 & (n1494 | n3934);
  assign n1602 = n1600 & n1601 & (n1593 | n1322);
  assign n1603 = ~Ni14 & ~n3796 & (n788 | ~n3797);
  assign n1604 = ~n1986 & n788 & Ni14 & ~n2254;
  assign n1605 = Ni12 & (n1603 | n1604 | ~n4250);
  assign n1606 = ~n1605 & (n1446 | (n4256 & n4257));
  assign n1607 = n1606 & (n1549 | n1553);
  assign n1608 = ~n1454 & ~n3677 & (n788 | ~n1463);
  assign n1609 = (Ni11 | n1607) & (n1549 | ~n3898);
  assign n1610 = n2254 | n3677;
  assign n1611 = ~n1608 & n1609 & (n1540 | n1610);
  assign n1612 = ~n796 & n1459 & (~n795 | n1461);
  assign n1613 = ~n796 & (n1523 | n3947);
  assign n1614 = (n4145 | n3948) & (n4146 | n2757);
  assign n1615 = n3859 | n795;
  assign n1616 = n1613 & n1614 & (n1525 | n1615);
  assign n1617 = ~n796 & (n1527 | n3947);
  assign n1618 = (n1420 | n3948) & (n4143 | n2757);
  assign n1619 = n1617 & n1618 & (n1529 | n1615);
  assign n1620 = ~n796 & (n1531 | n3947);
  assign n1621 = (n4136 | n3948) & (n1373 | n2757);
  assign n1622 = n1620 & n1621 & (n1533 | n1615);
  assign n1623 = (n1622 | n3864) & (n1619 | n3867);
  assign n1624 = n4296 & n4294 & (n1535 | n3946);
  assign n1625 = n1623 & n1624 & (n1616 | n1322);
  assign n1626 = ~n796 & (n1511 | n3947);
  assign n1627 = (n4140 | n3948) & (n4141 | n2757);
  assign n1628 = n1626 & n1627 & (n1513 | n1615);
  assign n1629 = ~n796 & (n1515 | n3947);
  assign n1630 = (n1407 | n3948) & (n4138 | n2757);
  assign n1631 = n1629 & n1630 & (n1517 | n1615);
  assign n1632 = ~n796 & (n1519 | n3947);
  assign n1633 = (n4135 | n3948) & (n1364 | n2757);
  assign n1634 = n1632 & n1633 & (n1521 | n1615);
  assign n1635 = (n1634 | n3864) & (n1631 | n3867);
  assign n1636 = n4293 & n4294 & (n1534 | n3946);
  assign n1637 = n1635 & n1636 & (n1628 | n1322);
  assign n1638 = ~n796 & (n1483 | n3947);
  assign n1639 = (n4159 | n3948) & (n4160 | n2757);
  assign n1640 = n1638 & n1639 & (n1485 | n1615);
  assign n1641 = ~n796 & (n1487 | n3947);
  assign n1642 = (n1444 | n3948) & (n4157 | n2757);
  assign n1643 = n1641 & n1642 & (n1489 | n1615);
  assign n1644 = ~n796 & (n1491 | n3947);
  assign n1645 = (n4150 | n3948) & (n1391 | n2757);
  assign n1646 = n1644 & n1645 & (n1493 | n1615);
  assign n1647 = (n1646 | n3864) & (n1643 | n3867);
  assign n1648 = n4297 & n4294 & (n1496 | n3946);
  assign n1649 = n1647 & n1648 & (n1640 | n1322);
  assign n1650 = ~n796 & (n1471 | n3947);
  assign n1651 = (n4154 | n3948) & (n4155 | n2757);
  assign n1652 = n1650 & n1651 & (n1473 | n1615);
  assign n1653 = ~n796 & (n1475 | n3947);
  assign n1654 = (n1432 | n3948) & (n4152 | n2757);
  assign n1655 = n1653 & n1654 & (n1477 | n1615);
  assign n1656 = ~n796 & (n1479 | n3947);
  assign n1657 = (n4149 | n3948) & (n1382 | n2757);
  assign n1658 = n1656 & n1657 & (n1481 | n1615);
  assign n1659 = (n1658 | n3864) & (n1655 | n3867);
  assign n1660 = n4295 & n4294 & (n1494 | n3946);
  assign n1661 = n1659 & n1660 & (n1652 | n1322);
  assign n1662 = ~Ni14 & ~n3796 & (n795 | ~n3797);
  assign n1663 = ~n1986 & n795 & Ni14 & ~n2254;
  assign n1664 = Ni12 & (n1662 | n1663 | ~n4292);
  assign n1665 = ~n1664 & (n1446 | (n4298 & n4299));
  assign n1666 = n1665 & (n1553 | n1612);
  assign n1667 = ~n1454 & ~n3677 & (n795 | ~n1463);
  assign n1668 = (Ni11 | n1666) & (n1612 | ~n3898);
  assign n1669 = ~n1667 & (n1540 | n1610) & n1668;
  assign n1670 = ~Ni9 & (~Ni8 | ~Ni7);
  assign n1671 = n1670 & (Ni10 | ~Ni7);
  assign n1672 = (n4129 | n1702) & (n1783 | n1408);
  assign n1673 = n1778 & n1359;
  assign n1674 = n1362 & n1672 & (n1673 | n914);
  assign n1675 = (n4131 | n1702) & (n1748 | n1408);
  assign n1676 = n1743 & n1369;
  assign n1677 = n1362 & n1675 & (n1676 | n914);
  assign n1678 = (n4130 | n1702) & (n1853 | n1408);
  assign n1679 = n1848 & n1378;
  assign n1680 = n1362 & n1678 & (n1679 | n914);
  assign n1681 = (n4132 | n1702) & (n1818 | n1408);
  assign n1682 = n1813 & n1387;
  assign n1683 = n1362 & n1681 & (n1682 | n914);
  assign n1684 = (n1764 | n3893) & (n4119 | n2109);
  assign n1685 = n1362 & (n4120 | n914);
  assign n1686 = n1766 & n1397;
  assign n1687 = n1684 & n1685 & (n1686 | n1408);
  assign n1688 = (n1728 | n3893) & (n4123 | n2109);
  assign n1689 = n1362 & (n4124 | n914);
  assign n1690 = n1731 & n1411;
  assign n1691 = n1688 & n1689 & (n1690 | n1408);
  assign n1692 = (n1834 | n3893) & (n4121 | n2109);
  assign n1693 = n1362 & (n4122 | n914);
  assign n1694 = n1836 & n1423;
  assign n1695 = n1692 & n1693 & (n1694 | n1408);
  assign n1696 = (n1799 | n3893) & (n4125 | n2109);
  assign n1697 = n1362 & (n4126 | n914);
  assign n1698 = n1801 & n1435;
  assign n1699 = n1696 & n1697 & (n1698 | n1408);
  assign n1700 = (Pi20 & n1368) | (n1366 & (~Pi20 | n1368));
  assign n1701 = Pi19 | n2254;
  assign n1702 = ~Pi19 | n2254;
  assign n1703 = (n1700 | n1701) & (n1370 | n1702);
  assign n1704 = (Pi20 & n1377) | (n1375 & (~Pi20 | n1377));
  assign n1705 = (n1704 | n1701) & (n1379 | n1702);
  assign n1706 = (Pi20 & n1386) | (n1384 & (~Pi20 | n1386));
  assign n1707 = (n1706 | n1701) & (n1388 | n1702);
  assign n1708 = (Pi20 & n1412) | (n1410 & (~Pi20 | n1412));
  assign n1709 = (Pi20 & n1416) | (n1414 & (~Pi20 | n1416));
  assign n1710 = (n1708 | n1701) & (n1709 | n1702);
  assign n1711 = (Pi20 & n1424) | (n1422 & (~Pi20 | n1424));
  assign n1712 = (Pi20 & n1428) | (n1426 & (~Pi20 | n1428));
  assign n1713 = (n1711 | n1701) & (n1712 | n1702);
  assign n1714 = (Pi20 & n1436) | (n1434 & (~Pi20 | n1436));
  assign n1715 = (Pi20 & n1440) | (n1438 & (~Pi20 | n1440));
  assign n1716 = (n1714 | n1701) & (n1715 | n1702);
  assign n1717 = n1446 | n4684 | n4685;
  assign n1718 = ~n4683 & (Pi17 | (n4127 & n4128));
  assign n1719 = n1717 & (n1718 | n1448);
  assign n1720 = ~n724 | n4767;
  assign n1721 = ~n724 & n1354;
  assign n1722 = n1354 & n1720 & (n18 | n1721);
  assign n1723 = ~n728 | n4767;
  assign n1724 = ~n728 & n1354;
  assign n1725 = n1354 & n1723 & (n18 | n1724);
  assign n1726 = (n1722 | n3915) & (n1725 | n3916);
  assign n1727 = ~n3918 & (n3917 | n4123);
  assign n1728 = n1720 & n1415;
  assign n1729 = ~n789 | n3857;
  assign n1730 = n1726 & n1727 & (n1728 | n1729);
  assign n1731 = ~n717 | n4767;
  assign n1732 = ~n717 & n1354;
  assign n1733 = n1354 & n1731 & (n18 | n1732);
  assign n1734 = ~n720 | n4767;
  assign n1735 = ~n720 & n1354;
  assign n1736 = n1354 & n1734 & (n18 | n1735);
  assign n1737 = (n1733 | n3915) & (n1736 | n3916);
  assign n1738 = ~n3918 & (n3917 | n4124);
  assign n1739 = n1737 & n1738 & (n1690 | n1729);
  assign n1740 = ~n732 | n4767;
  assign n1741 = ~n732 & n1354;
  assign n1742 = n1354 & n1740 & (n18 | n1741);
  assign n1743 = ~n736 | n4767;
  assign n1744 = ~n736 & n1354;
  assign n1745 = n1354 & n1743 & (n18 | n1744);
  assign n1746 = (n1742 | n3915) & (n1745 | n3916);
  assign n1747 = ~n3918 & (n1676 | n3917);
  assign n1748 = n1740 & n1367;
  assign n1749 = n1746 & n1747 & (n1748 | n1729);
  assign n1750 = ~n739 | n4767;
  assign n1751 = ~n739 & n1354;
  assign n1752 = n1354 & n1750 & (n18 | n1751);
  assign n1753 = (n1749 | n3864) & (n1739 | n3867);
  assign n1754 = n4244 & n4242 & (n4131 | n3914);
  assign n1755 = n1753 & n1754 & (n1730 | n1322);
  assign n1756 = ~n699 | n4767;
  assign n1757 = ~n699 & n1354;
  assign n1758 = n1354 & n1756 & (n18 | n1757);
  assign n1759 = ~n703 | n4767;
  assign n1760 = ~n703 & n1354;
  assign n1761 = n1354 & n1759 & (n18 | n1760);
  assign n1762 = (n1758 | n3915) & (n1761 | n3916);
  assign n1763 = ~n3918 & (n3917 | n4119);
  assign n1764 = n1756 & n1402;
  assign n1765 = n1762 & n1763 & (n1764 | n1729);
  assign n1766 = ~n691 | n4767;
  assign n1767 = ~n691 & n1354;
  assign n1768 = n1354 & n1766 & (n18 | n1767);
  assign n1769 = ~n694 | n4767;
  assign n1770 = ~n694 & n1354;
  assign n1771 = n1354 & n1769 & (n18 | n1770);
  assign n1772 = (n1768 | n3915) & (n1771 | n3916);
  assign n1773 = ~n3918 & (n3917 | n4120);
  assign n1774 = n1772 & n1773 & (n1686 | n1729);
  assign n1775 = ~n707 | n4767;
  assign n1776 = ~n707 & n1354;
  assign n1777 = n1354 & n1775 & (n18 | n1776);
  assign n1778 = ~n711 | n4767;
  assign n1779 = ~n711 & n1354;
  assign n1780 = n1354 & n1778 & (n18 | n1779);
  assign n1781 = (n1777 | n3915) & (n1780 | n3916);
  assign n1782 = ~n3918 & (n1673 | n3917);
  assign n1783 = n1775 & n1357;
  assign n1784 = n1781 & n1782 & (n1783 | n1729);
  assign n1785 = ~n714 | n4767;
  assign n1786 = ~n714 & n1354;
  assign n1787 = n1354 & n1785 & (n18 | n1786);
  assign n1788 = (n1784 | n3864) & (n1774 | n3867);
  assign n1789 = n4241 & n4242 & (n4129 | n3914);
  assign n1790 = n1788 & n1789 & (n1765 | n1322);
  assign n1791 = ~n755 | n4767;
  assign n1792 = ~n755 & n1354;
  assign n1793 = n1354 & n1791 & (n18 | n1792);
  assign n1794 = ~n757 | n4767;
  assign n1795 = ~n757 & n1354;
  assign n1796 = n1354 & n1794 & (n18 | n1795);
  assign n1797 = (n1793 | n3915) & (n1796 | n3916);
  assign n1798 = ~n3918 & (n3917 | n4125);
  assign n1799 = n1791 & n1439;
  assign n1800 = n1797 & n1798 & (n1799 | n1729);
  assign n1801 = ~n752 | n4767;
  assign n1802 = ~n752 & n1354;
  assign n1803 = n1354 & n1801 & (n18 | n1802);
  assign n1804 = ~n753 | n4767;
  assign n1805 = ~n753 & n1354;
  assign n1806 = n1354 & n1804 & (n18 | n1805);
  assign n1807 = (n1803 | n3915) & (n1806 | n3916);
  assign n1808 = ~n3918 & (n3917 | n4126);
  assign n1809 = n1807 & n1808 & (n1698 | n1729);
  assign n1810 = ~n759 | n4767;
  assign n1811 = ~n759 & n1354;
  assign n1812 = n1354 & n1810 & (n18 | n1811);
  assign n1813 = ~n761 | n4767;
  assign n1814 = ~n761 & n1354;
  assign n1815 = n1354 & n1813 & (n18 | n1814);
  assign n1816 = (n1812 | n3915) & (n1815 | n3916);
  assign n1817 = ~n3918 & (n1682 | n3917);
  assign n1818 = n1810 & n1385;
  assign n1819 = n1816 & n1817 & (n1818 | n1729);
  assign n1820 = n4767 | n1468;
  assign n1821 = n1468 & n1354;
  assign n1822 = n1354 & n1820 & (n18 | n1821);
  assign n1823 = (n1819 | n3864) & (n1809 | n3867);
  assign n1824 = n4245 & n4242 & (n4132 | n3914);
  assign n1825 = n1823 & n1824 & (n1800 | n1322);
  assign n1826 = ~n745 | n4767;
  assign n1827 = ~n745 & n1354;
  assign n1828 = n1354 & n1826 & (n18 | n1827);
  assign n1829 = ~n747 | n4767;
  assign n1830 = ~n747 & n1354;
  assign n1831 = n1354 & n1829 & (n18 | n1830);
  assign n1832 = (n1828 | n3915) & (n1831 | n3916);
  assign n1833 = ~n3918 & (n3917 | n4121);
  assign n1834 = n1826 & n1427;
  assign n1835 = n1832 & n1833 & (n1834 | n1729);
  assign n1836 = ~n742 | n4767;
  assign n1837 = ~n742 & n1354;
  assign n1838 = n1354 & n1836 & (n18 | n1837);
  assign n1839 = ~n743 | n4767;
  assign n1840 = ~n743 & n1354;
  assign n1841 = n1354 & n1839 & (n18 | n1840);
  assign n1842 = (n1838 | n3915) & (n1841 | n3916);
  assign n1843 = ~n3918 & (n3917 | n4122);
  assign n1844 = n1842 & n1843 & (n1694 | n1729);
  assign n1845 = ~n749 | n4767;
  assign n1846 = ~n749 & n1354;
  assign n1847 = n1354 & n1845 & (n18 | n1846);
  assign n1848 = ~n751 | n4767;
  assign n1849 = ~n751 & n1354;
  assign n1850 = n1354 & n1848 & (n18 | n1849);
  assign n1851 = (n1847 | n3915) & (n1850 | n3916);
  assign n1852 = ~n3918 & (n1679 | n3917);
  assign n1853 = n1845 & n1376;
  assign n1854 = n1851 & n1852 & (n1853 | n1729);
  assign n1855 = n4767 | n1465;
  assign n1856 = n1465 & n1354;
  assign n1857 = n1354 & n1855 & (n18 | n1856);
  assign n1858 = (n1854 | n3864) & (n1844 | n3867);
  assign n1859 = n4243 & n4242 & (n4130 | n3914);
  assign n1860 = n1858 & n1859 & (n1835 | n1322);
  assign n1861 = ~n2272 & (~n4226 | ~n4227);
  assign n1862 = ~n2272 & (~n4207 | ~n4208);
  assign n1863 = n3696 | n4680 | n4682;
  assign n1864 = n1719 & (n2632 | (n4247 & n4246));
  assign n1865 = n1863 & n1864 & (n1718 | n1452);
  assign n1866 = (n1722 | n3901) & (n1725 | n3902);
  assign n1867 = n1455 & (n4123 | n3903);
  assign n1868 = ~n3761 | n3857;
  assign n1869 = n1866 & n1867 & (n1728 | n1868);
  assign n1870 = (n1733 | n3901) & (n1736 | n3902);
  assign n1871 = n1455 & (n4124 | n3903);
  assign n1872 = n1870 & n1871 & (n1690 | n1868);
  assign n1873 = (n1742 | n3901) & (n1745 | n3902);
  assign n1874 = n1455 & (n1676 | n3903);
  assign n1875 = n1873 & n1874 & (n1748 | n1868);
  assign n1876 = (n1875 | n3864) & (n1872 | n3867);
  assign n1877 = n4201 & n4199 & (n4131 | n3900);
  assign n1878 = n1876 & n1877 & (n1869 | n1322);
  assign n1879 = (n1758 | n3901) & (n1761 | n3902);
  assign n1880 = n1455 & (n4119 | n3903);
  assign n1881 = n1879 & n1880 & (n1764 | n1868);
  assign n1882 = (n1768 | n3901) & (n1771 | n3902);
  assign n1883 = n1455 & (n4120 | n3903);
  assign n1884 = n1882 & n1883 & (n1686 | n1868);
  assign n1885 = (n1777 | n3901) & (n1780 | n3902);
  assign n1886 = n1455 & (n1673 | n3903);
  assign n1887 = n1885 & n1886 & (n1783 | n1868);
  assign n1888 = (n1887 | n3864) & (n1884 | n3867);
  assign n1889 = n4198 & n4199 & (n4129 | n3900);
  assign n1890 = n1888 & n1889 & (n1881 | n1322);
  assign n1891 = (n1793 | n3901) & (n1796 | n3902);
  assign n1892 = n1455 & (n4125 | n3903);
  assign n1893 = n1891 & n1892 & (n1799 | n1868);
  assign n1894 = (n1803 | n3901) & (n1806 | n3902);
  assign n1895 = n1455 & (n4126 | n3903);
  assign n1896 = n1894 & n1895 & (n1698 | n1868);
  assign n1897 = (n1812 | n3901) & (n1815 | n3902);
  assign n1898 = n1455 & (n1682 | n3903);
  assign n1899 = n1897 & n1898 & (n1818 | n1868);
  assign n1900 = (n1899 | n3864) & (n1896 | n3867);
  assign n1901 = n4202 & n4199 & (n4132 | n3900);
  assign n1902 = n1900 & n1901 & (n1893 | n1322);
  assign n1903 = (n1828 | n3901) & (n1831 | n3902);
  assign n1904 = n1455 & (n4121 | n3903);
  assign n1905 = n1903 & n1904 & (n1834 | n1868);
  assign n1906 = (n1838 | n3901) & (n1841 | n3902);
  assign n1907 = n1455 & (n4122 | n3903);
  assign n1908 = n1906 & n1907 & (n1694 | n1868);
  assign n1909 = (n1847 | n3901) & (n1850 | n3902);
  assign n1910 = n1455 & (n1679 | n3903);
  assign n1911 = n1909 & n1910 & (n1853 | n1868);
  assign n1912 = (n1911 | n3864) & (n1908 | n3867);
  assign n1913 = n4200 & n4199 & (n4130 | n3900);
  assign n1914 = n1912 & n1913 & (n1905 | n1322);
  assign n1915 = (n1878 | n3884) & (n1902 | n3891);
  assign n1916 = (n1890 | n3870) & (n1914 | n3877);
  assign n1917 = n1915 & n1916;
  assign n1918 = ~Ni30 & n1540;
  assign n1919 = Pi25 | n2254;
  assign n1920 = n1362 & (n1918 | n1919);
  assign n1921 = n1920 & (n1929 | (n4118 & n4116));
  assign n1922 = n1379 & (~Pi16 | n1388);
  assign n1923 = ~Pi25 | n3848;
  assign n1924 = n1921 & (n1922 | n1923);
  assign n1925 = n1920 & (n1929 | (n4114 & n4112));
  assign n1926 = n1360 & (~Pi16 | n1370);
  assign n1927 = n1925 & (n1926 | n1923);
  assign n1928 = (n4149 | n3858) & (n1382 | n3860);
  assign n1929 = ~Pi25 | n2254;
  assign n1930 = n1928 & (n1704 | n1929);
  assign n1931 = ~n3740 & ((~n1706 & ~n1929) | ~n4151);
  assign n1932 = ~n2272 & ((~n1711 & ~n1929) | ~n4153);
  assign n1933 = ~n3895 & ((~n1712 & ~n1929) | ~n4156);
  assign n1934 = ~n3743 & ((~n1714 & ~n1929) | ~n4158);
  assign n1935 = ~n3737 & ((~n1715 & ~n1929) | ~n4161);
  assign n1936 = (n4135 | n3858) & (n1364 | n3860);
  assign n1937 = (Pi20 & n1358) | (n1356 & (~Pi20 | n1358));
  assign n1938 = n1936 & (n1937 | n1929);
  assign n1939 = ~n3740 & ((~n1700 & ~n1929) | ~n4137);
  assign n1940 = ~n2272 & ((~n1929 & ~n1961) | ~n4139);
  assign n1941 = ~n3895 & ((~n1929 & ~n1958) | ~n4142);
  assign n1942 = ~n3743 & ((~n1708 & ~n1929) | ~n4144);
  assign n1943 = ~n3737 & ((~n1709 & ~n1929) | ~n4147);
  assign n1944 = (~Pi15 & n1927) | (n1924 & (Pi15 | n1927));
  assign n1945 = (n1448 | n1944) & (n1446 | ~n3990);
  assign n1946 = n1455 & (n1541 | n1919);
  assign n1947 = (n1721 | n3931) & (n1724 | n3932);
  assign n1948 = n1929 | ~n3761;
  assign n1949 = n1946 & n1947 & (n1709 | n1948);
  assign n1950 = (n1732 | n3931) & (n1735 | n3932);
  assign n1951 = n1946 & n1950 & (n1708 | n1948);
  assign n1952 = (n1741 | n3931) & (n1744 | n3932);
  assign n1953 = n1946 & n1952 & (n1700 | n1948);
  assign n1954 = (n1953 | n3864) & (n1951 | n3867);
  assign n1955 = n4190 & n4188 & (n1370 | n3930);
  assign n1956 = n1954 & n1955 & (n1949 | n1322);
  assign n1957 = (n1757 | n3931) & (n1760 | n3932);
  assign n1958 = (Pi20 & n1403) | (n1401 & (~Pi20 | n1403));
  assign n1959 = n1946 & n1957 & (n1958 | n1948);
  assign n1960 = (n1767 | n3931) & (n1770 | n3932);
  assign n1961 = (Pi20 & n1399) | (n1396 & (~Pi20 | n1399));
  assign n1962 = n1946 & n1960 & (n1961 | n1948);
  assign n1963 = (n1776 | n3931) & (n1779 | n3932);
  assign n1964 = n1946 & n1963 & (n1937 | n1948);
  assign n1965 = (n1964 | n3864) & (n1962 | n3867);
  assign n1966 = n4187 & n4188 & (n1360 | n3930);
  assign n1967 = n1965 & n1966 & (n1959 | n1322);
  assign n1968 = (n1792 | n3931) & (n1795 | n3932);
  assign n1969 = n1946 & n1968 & (n1715 | n1948);
  assign n1970 = (n1802 | n3931) & (n1805 | n3932);
  assign n1971 = n1946 & n1970 & (n1714 | n1948);
  assign n1972 = (n1811 | n3931) & (n1814 | n3932);
  assign n1973 = n1946 & n1972 & (n1706 | n1948);
  assign n1974 = (n1973 | n3864) & (n1971 | n3867);
  assign n1975 = n4191 & n4188 & (n1388 | n3930);
  assign n1976 = n1974 & n1975 & (n1969 | n1322);
  assign n1977 = (n1827 | n3931) & (n1830 | n3932);
  assign n1978 = n1946 & n1977 & (n1712 | n1948);
  assign n1979 = (n1837 | n3931) & (n1840 | n3932);
  assign n1980 = n1946 & n1979 & (n1711 | n1948);
  assign n1981 = (n1846 | n3931) & (n1849 | n3932);
  assign n1982 = n1946 & n1981 & (n1704 | n1948);
  assign n1983 = (n1982 | n3864) & (n1980 | n3867);
  assign n1984 = n4189 & n4188 & (n1379 | n3930);
  assign n1985 = n1983 & n1984 & (n1978 | n1322);
  assign n1986 = n3793 & (Pi27 | n1918);
  assign n1987 = n1552 & (n1986 | n1919);
  assign n1988 = (n1709 | n3922) & (n1721 | n3923);
  assign n1989 = ~Pi27 | n1314;
  assign n1990 = n1987 & n1988 & (n1724 | n1989);
  assign n1991 = (n1708 | n3922) & (n1732 | n3923);
  assign n1992 = n1987 & n1991 & (n1735 | n1989);
  assign n1993 = (n1700 | n3922) & (n1741 | n3923);
  assign n1994 = n1987 & n1993 & (n1744 | n1989);
  assign n1995 = (n1994 | n3864) & (n1992 | n3867);
  assign n1996 = n4183 & n4181 & (n1751 | n3921);
  assign n1997 = n1995 & n1996 & (n1990 | n1322);
  assign n1998 = (n1958 | n3922) & (n1757 | n3923);
  assign n1999 = n1987 & n1998 & (n1760 | n1989);
  assign n2000 = (n1961 | n3922) & (n1767 | n3923);
  assign n2001 = n1987 & n2000 & (n1770 | n1989);
  assign n2002 = (n1937 | n3922) & (n1776 | n3923);
  assign n2003 = n1987 & n2002 & (n1779 | n1989);
  assign n2004 = (n2003 | n3864) & (n2001 | n3867);
  assign n2005 = n4180 & n4181 & (n1786 | n3921);
  assign n2006 = n2004 & n2005 & (n1999 | n1322);
  assign n2007 = (n1715 | n3922) & (n1792 | n3923);
  assign n2008 = n1987 & n2007 & (n1795 | n1989);
  assign n2009 = (n1714 | n3922) & (n1802 | n3923);
  assign n2010 = n1987 & n2009 & (n1805 | n1989);
  assign n2011 = (n1706 | n3922) & (n1811 | n3923);
  assign n2012 = n1987 & n2011 & (n1814 | n1989);
  assign n2013 = (n2012 | n3864) & (n2010 | n3867);
  assign n2014 = n4184 & n4181 & (n1821 | n3921);
  assign n2015 = n2013 & n2014 & (n2008 | n1322);
  assign n2016 = (n1712 | n3922) & (n1827 | n3923);
  assign n2017 = n1987 & n2016 & (n1830 | n1989);
  assign n2018 = (n1711 | n3922) & (n1837 | n3923);
  assign n2019 = n1987 & n2018 & (n1840 | n1989);
  assign n2020 = (n1704 | n3922) & (n1846 | n3923);
  assign n2021 = n1987 & n2020 & (n1849 | n1989);
  assign n2022 = (n2021 | n3864) & (n2019 | n3867);
  assign n2023 = n4182 & n4181 & (n1856 | n3921);
  assign n2024 = n2022 & n2023 & (n2017 | n1322);
  assign n2025 = (~Pi26 | n1918) & n3794;
  assign n2026 = ~n3918 & (n1919 | n2025);
  assign n2027 = (n1721 | n3926) & (n1724 | n3927);
  assign n2028 = ~n789 | n1929;
  assign n2029 = n2026 & n2027 & (n1709 | n2028);
  assign n2030 = (n1732 | n3926) & (n1735 | n3927);
  assign n2031 = n2026 & n2030 & (n1708 | n2028);
  assign n2032 = (n1741 | n3926) & (n1744 | n3927);
  assign n2033 = n2026 & n2032 & (n1700 | n2028);
  assign n2034 = (n2033 | n3864) & (n2031 | n3867);
  assign n2035 = n4176 & n4174 & (n1370 | n3925);
  assign n2036 = n2034 & n2035 & (n2029 | n1322);
  assign n2037 = (n1757 | n3926) & (n1760 | n3927);
  assign n2038 = n2026 & n2037 & (n1958 | n2028);
  assign n2039 = (n1767 | n3926) & (n1770 | n3927);
  assign n2040 = n2026 & n2039 & (n1961 | n2028);
  assign n2041 = (n1776 | n3926) & (n1779 | n3927);
  assign n2042 = n2026 & n2041 & (n1937 | n2028);
  assign n2043 = (n2042 | n3864) & (n2040 | n3867);
  assign n2044 = n4173 & n4174 & (n1360 | n3925);
  assign n2045 = n2043 & n2044 & (n2038 | n1322);
  assign n2046 = (n1792 | n3926) & (n1795 | n3927);
  assign n2047 = n2026 & n2046 & (n1715 | n2028);
  assign n2048 = (n1802 | n3926) & (n1805 | n3927);
  assign n2049 = n2026 & n2048 & (n1714 | n2028);
  assign n2050 = (n1811 | n3926) & (n1814 | n3927);
  assign n2051 = n2026 & n2050 & (n1706 | n2028);
  assign n2052 = (n2051 | n3864) & (n2049 | n3867);
  assign n2053 = n4177 & n4174 & (n1388 | n3925);
  assign n2054 = n2052 & n2053 & (n2047 | n1322);
  assign n2055 = (n1827 | n3926) & (n1830 | n3927);
  assign n2056 = n2026 & n2055 & (n1712 | n2028);
  assign n2057 = (n1837 | n3926) & (n1840 | n3927);
  assign n2058 = n2026 & n2057 & (n1711 | n2028);
  assign n2059 = (n1846 | n3926) & (n1849 | n3927);
  assign n2060 = n2026 & n2059 & (n1704 | n2028);
  assign n2061 = (n2060 | n3864) & (n2058 | n3867);
  assign n2062 = n4175 & n4174 & (n1379 | n3925);
  assign n2063 = n2061 & n2062 & (n2056 | n1322);
  assign n2064 = (n1611 | n3937) & (n3805 | ~n3992);
  assign n2065 = (n1669 | n3766) & (n1458 | n1671);
  assign n2066 = ~Ni10 | n3768;
  assign n2067 = n2064 & n2065 & (n2066 | ~n4773);
  assign n2068 = (n1449 | Ni11) & (n1447 | ~n1543);
  assign n2069 = (n1945 | n3897) & (~n1543 | ~n3989);
  assign n2070 = Ni11 | ~Ni10;
  assign n2071 = n2069 & (n1719 | n2070);
  assign n2072 = Ni7 & n2398;
  assign n2073 = n2398 & ~Ni7;
  assign n2074 = Ni9 | Ni8;
  assign n2075 = ~n2068 & (n2072 | (n2073 & n2074));
  assign n2076 = ~n3896 | n2067 | n3707;
  assign n2077 = ~n2075 & (n2071 | ~n2073 | n2074);
  assign n2078 = ~Ni32 & ~Ni30;
  assign n2079 = ~n18 | n1539;
  assign n2080 = ~Ni34 | ~Ni33;
  assign n2081 = ~n792 & (n2079 | n2080);
  assign n2082 = (~Ni34 | n821) & n2081;
  assign n2083 = (~Ni34 | n857) & n2081;
  assign n2084 = (~Ni34 | n895) & n2081;
  assign n2085 = ~Ni34 | ~n793;
  assign n2086 = (n2082 | n1408) & (n2083 | n914);
  assign n2087 = n2085 & n2086 & (n2084 | n1702);
  assign n2088 = (~Ni34 | n922) & n2081;
  assign n2089 = (~Ni34 | n947) & n2081;
  assign n2090 = (~Ni34 | n974) & n2081;
  assign n2091 = (n2088 | n1408) & (n2089 | n914);
  assign n2092 = n2085 & n2091 & (n2090 | n1702);
  assign n2093 = (~Ni34 | n984) & n2081;
  assign n2094 = (~Ni34 | n1001_1) & n2081;
  assign n2095 = (~Ni34 | n882) & n2081;
  assign n2096 = (n2093 | n1408) & (n2094 | n914);
  assign n2097 = n2085 & n2096 & (n2095 | n1702);
  assign n2098 = (~Ni34 | n1021_1) & n2081;
  assign n2099 = (~Ni34 | n1028) & n2081;
  assign n2100 = (~Ni34 | n966) & n2081;
  assign n2101 = (n2098 | n1408) & (n2099 | n914);
  assign n2102 = n2085 & n2101 & (n2100 | n1702);
  assign n2103 = (~Ni34 | n1049) & n2081;
  assign n2104 = (~Ni34 | n1065) & n2081;
  assign n2105 = (~Ni34 | n1081_1) & n2081;
  assign n2106 = (~Ni34 | n1108) & n2081;
  assign n2107 = n2085 & (n2105 | n3893);
  assign n2108 = (n2103 | n1408) & (n2104 | n914);
  assign n2109 = ~Pi19 | n3859;
  assign n2110 = n2107 & n2108 & (n2106 | n2109);
  assign n2111 = (~Ni34 | n1135) & n2081;
  assign n2112 = (~Ni34 | n1149) & n2081;
  assign n2113 = (~Ni34 | n1165) & n2081;
  assign n2114 = (~Ni34 | n1189) & n2081;
  assign n2115 = n2085 & (n2113 | n3893);
  assign n2116 = (n2111 | n1408) & (n2112 | n914);
  assign n2117 = n2115 & n2116 & (n2114 | n2109);
  assign n2118 = (~Ni34 | n1217) & n2081;
  assign n2119 = (~Ni34 | n1228) & n2081;
  assign n2120 = (~Ni34 | n1235) & n2081;
  assign n2121 = (~Ni34 | n1247) & n2081;
  assign n2122 = n2085 & (n2120 | n3893);
  assign n2123 = (n2118 | n1408) & (n2119 | n914);
  assign n2124 = n2122 & n2123 & (n2121 | n2109);
  assign n2125 = (~Ni34 | n1259) & n2081;
  assign n2126 = (~Ni34 | n1266) & n2081;
  assign n2127 = (~Ni34 | n1273) & n2081;
  assign n2128 = (~Ni34 | n1280) & n2081;
  assign n2129 = n2085 & (n2127 | n3893);
  assign n2130 = (n2125 | n1408) & (n2126 | n914);
  assign n2131 = n2129 & n2130 & (n2128 | n2109);
  assign n2132 = n2080 & (~Ni33 | ~n821);
  assign n2133 = (n2132 | n3949) & (~n821 | n3951);
  assign n2134 = (n821 & n4691) | (n4690 & (~n821 | n4691));
  assign n2135 = n2082 & n2133 & (~Pi25 | n2134);
  assign n2136 = n2080 & (~Ni33 | ~n857);
  assign n2137 = (n2136 | n3949) & (~n857 | n3951);
  assign n2138 = (n857 & n4691) | (n4690 & (~n857 | n4691));
  assign n2139 = n2083 & n2137 & (~Pi25 | n2138);
  assign n2140 = n2080 & (~Ni33 | ~n895);
  assign n2141 = (n2140 | n3949) & (~n895 | n3951);
  assign n2142 = (n895 & n4691) | (n4690 & (~n895 | n4691));
  assign n2143 = n2084 & n2141 & (~Pi25 | n2142);
  assign n2144 = (n2135 | n1408) & (n2139 | n914);
  assign n2145 = n2085 & n2144 & (n2143 | n1702);
  assign n2146 = n2080 & (~Ni33 | ~n922);
  assign n2147 = (n2146 | n3949) & (~n922 | n3951);
  assign n2148 = (n922 & n4691) | (n4690 & (~n922 | n4691));
  assign n2149 = n2088 & n2147 & (~Pi25 | n2148);
  assign n2150 = n2080 & (~Ni33 | ~n947);
  assign n2151 = (n2150 | n3949) & (~n947 | n3951);
  assign n2152 = (n947 & n4691) | (n4690 & (~n947 | n4691));
  assign n2153 = n2089 & n2151 & (~Pi25 | n2152);
  assign n2154 = n2080 & (~Ni33 | ~n974);
  assign n2155 = (n2154 | n3949) & (~n974 | n3951);
  assign n2156 = (n974 & n4691) | (n4690 & (~n974 | n4691));
  assign n2157 = n2090 & n2155 & (~Pi25 | n2156);
  assign n2158 = (n2149 | n1408) & (n2153 | n914);
  assign n2159 = n2085 & n2158 & (n2157 | n1702);
  assign n2160 = n2080 & (~Ni33 | ~n984);
  assign n2161 = (n2160 | n3949) & (~n984 | n3951);
  assign n2162 = (n984 & n4691) | (n4690 & (~n984 | n4691));
  assign n2163 = n2093 & n2161 & (~Pi25 | n2162);
  assign n2164 = n2080 & (~Ni33 | ~n1001_1);
  assign n2165 = (n2164 | n3949) & (~n1001_1 | n3951);
  assign n2166 = (n1001_1 & n4691) | (n4690 & (~n1001_1 | n4691));
  assign n2167 = n2094 & n2165 & (~Pi25 | n2166);
  assign n2168 = n2080 & (~Ni33 | ~n882);
  assign n2169 = (n2168 | n3949) & (~n882 | n3951);
  assign n2170 = (n882 & n4691) | (n4690 & (~n882 | n4691));
  assign n2171 = n2095 & n2169 & (~Pi25 | n2170);
  assign n2172 = (n2163 | n1408) & (n2167 | n914);
  assign n2173 = n2085 & n2172 & (n2171 | n1702);
  assign n2174 = n2080 & (~Ni33 | ~n1021_1);
  assign n2175 = (n2174 | n3949) & (~n1021_1 | n3951);
  assign n2176 = (n1021_1 & n4691) | (n4690 & (~n1021_1 | n4691));
  assign n2177 = n2098 & n2175 & (~Pi25 | n2176);
  assign n2178 = n2080 & (~Ni33 | ~n1028);
  assign n2179 = (n2178 | n3949) & (~n1028 | n3951);
  assign n2180 = (n1028 & n4691) | (n4690 & (~n1028 | n4691));
  assign n2181 = n2099 & n2179 & (~Pi25 | n2180);
  assign n2182 = n2080 & (~Ni33 | ~n966);
  assign n2183 = (n2182 | n3949) & (~n966 | n3951);
  assign n2184 = (n966 & n4691) | (n4690 & (~n966 | n4691));
  assign n2185 = n2100 & n2183 & (~Pi25 | n2184);
  assign n2186 = (n2177 | n1408) & (n2181 | n914);
  assign n2187 = n2085 & n2186 & (n2185 | n1702);
  assign n2188 = n2080 & (~Ni33 | ~n1049);
  assign n2189 = (n2188 | n3949) & (~n1049 | n3951);
  assign n2190 = (n1049 & n4691) | (n4690 & (~n1049 | n4691));
  assign n2191 = n2103 & n2189 & (~Pi25 | n2190);
  assign n2192 = n2080 & (~Ni33 | ~n1065);
  assign n2193 = (n2192 | n3949) & (~n1065 | n3951);
  assign n2194 = (n1065 & n4691) | (n4690 & (~n1065 | n4691));
  assign n2195 = n2104 & n2193 & (~Pi25 | n2194);
  assign n2196 = n2080 & (~Ni33 | ~n1081_1);
  assign n2197 = n2080 & (~Ni33 | ~n1108);
  assign n2198 = (n2197 | n3949) & (~n1108 | n3951);
  assign n2199 = (n1108 & n4691) | (n4690 & (~n1108 | n4691));
  assign n2200 = n2106 & n2198 & (~Pi25 | n2199);
  assign n2201 = n2085 & (n3893 | (n4309 & n4308));
  assign n2202 = (n2191 | n1408) & (n2195 | n914);
  assign n2203 = n2201 & n2202 & (n2200 | n2109);
  assign n2204 = n2080 & (~Ni33 | ~n1135);
  assign n2205 = (n2204 | n3949) & (~n1135 | n3951);
  assign n2206 = (n1135 & n4691) | (n4690 & (~n1135 | n4691));
  assign n2207 = n2111 & n2205 & (~Pi25 | n2206);
  assign n2208 = n2080 & (~Ni33 | ~n1149);
  assign n2209 = (n2208 | n3949) & (~n1149 | n3951);
  assign n2210 = (n1149 & n4691) | (n4690 & (~n1149 | n4691));
  assign n2211 = n2112 & n2209 & (~Pi25 | n2210);
  assign n2212 = n2080 & (~Ni33 | ~n1165);
  assign n2213 = n2080 & (~Ni33 | ~n1189);
  assign n2214 = (n2213 | n3949) & (~n1189 | n3951);
  assign n2215 = (n1189 & n4691) | (n4690 & (~n1189 | n4691));
  assign n2216 = n2114 & n2214 & (~Pi25 | n2215);
  assign n2217 = n2085 & (n3893 | (n4313 & n4312));
  assign n2218 = (n2207 | n1408) & (n2211 | n914);
  assign n2219 = n2217 & n2218 & (n2216 | n2109);
  assign n2220 = n2080 & (~Ni33 | ~n1217);
  assign n2221 = (n2220 | n3949) & (~n1217 | n3951);
  assign n2222 = (n1217 & n4691) | (n4690 & (~n1217 | n4691));
  assign n2223 = n2118 & n2221 & (~Pi25 | n2222);
  assign n2224 = n2080 & (~Ni33 | ~n1228);
  assign n2225 = (n2224 | n3949) & (~n1228 | n3951);
  assign n2226 = (n1228 & n4691) | (n4690 & (~n1228 | n4691));
  assign n2227 = n2119 & n2225 & (~Pi25 | n2226);
  assign n2228 = n2080 & (~Ni33 | ~n1235);
  assign n2229 = n2080 & (~Ni33 | ~n1247);
  assign n2230 = (n2229 | n3949) & (~n1247 | n3951);
  assign n2231 = (n1247 & n4691) | (n4690 & (~n1247 | n4691));
  assign n2232 = n2121 & n2230 & (~Pi25 | n2231);
  assign n2233 = n2085 & (n3893 | (n4311 & n4310));
  assign n2234 = (n2223 | n1408) & (n2227 | n914);
  assign n2235 = n2233 & n2234 & (n2232 | n2109);
  assign n2236 = n2080 & (~Ni33 | ~n1259);
  assign n2237 = (n2236 | n3949) & (~n1259 | n3951);
  assign n2238 = (n1259 & n4691) | (n4690 & (~n1259 | n4691));
  assign n2239 = n2125 & n2237 & (~Pi25 | n2238);
  assign n2240 = n2080 & (~Ni33 | ~n1266);
  assign n2241 = (n2240 | n3949) & (~n1266 | n3951);
  assign n2242 = (n1266 & n4691) | (n4690 & (~n1266 | n4691));
  assign n2243 = n2126 & n2241 & (~Pi25 | n2242);
  assign n2244 = n2080 & (~Ni33 | ~n1273);
  assign n2245 = n2080 & (~Ni33 | ~n1280);
  assign n2246 = (n2245 | n3949) & (~n1280 | n3951);
  assign n2247 = (n1280 & n4691) | (n4690 & (~n1280 | n4691));
  assign n2248 = n2128 & n2246 & (~Pi25 | n2247);
  assign n2249 = n2085 & (n3893 | (n4315 & n4314));
  assign n2250 = (n2239 | n1408) & (n2243 | n914);
  assign n2251 = n2249 & n2250 & (n2248 | n2109);
  assign n2252 = ~n792 & n2085;
  assign n2253 = (n882 | n3954) & (n2168 | n3952);
  assign n2254 = ~Pi22 | ~Pi21;
  assign n2255 = n2252 & n2253 & (n2170 | n2254);
  assign n2256 = (n966 | n3954) & (n2182 | n3952);
  assign n2257 = n2252 & n2256 & (n2184 | n2254);
  assign n2258 = (n1228 | n3954) & (n2224 | n3952);
  assign n2259 = n2252 & n2258 & (n2226 | n2254);
  assign n2260 = (n1247 | n3954) & (n2229 | n3952);
  assign n2261 = n2252 & n2260 & (n2231 | n2254);
  assign n2262 = (n1001_1 | n3954) & (n2164 | n3952);
  assign n2263 = n2252 & n2262 & (n2166 | n2254);
  assign n2264 = (n1266 | n3954) & (n2240 | n3952);
  assign n2265 = n2252 & n2264 & (n2242 | n2254);
  assign n2266 = (n1280 | n3954) & (n2245 | n3952);
  assign n2267 = n2252 & n2266 & (n2247 | n2254);
  assign n2268 = (n1028 | n3954) & (n2178 | n3952);
  assign n2269 = n2252 & n2268 & (n2180 | n2254);
  assign n2270 = (n2263 | n3894) & (n2269 | n3740);
  assign n2271 = n4370 & (n2267 | n3737);
  assign n2272 = Pi16 | n3867;
  assign n2273 = n2270 & n2271 & (n2259 | n2272);
  assign n2274 = (n1217 | n3954) & (n2220 | n3952);
  assign n2275 = n2252 & n2274 & (n2222 | n2254);
  assign n2276 = (n1235 | n3954) & (n2228 | n3952);
  assign n2277 = (n1235 & n4691) | (n4690 & (~n1235 | n4691));
  assign n2278 = n2252 & n2276 & (n2277 | n2254);
  assign n2279 = (n984 | n3954) & (n2160 | n3952);
  assign n2280 = n2252 & n2279 & (n2162 | n2254);
  assign n2281 = (n1259 | n3954) & (n2236 | n3952);
  assign n2282 = n2252 & n2281 & (n2238 | n2254);
  assign n2283 = (n1273 | n3954) & (n2244 | n3952);
  assign n2284 = (n1273 & n4691) | (n4690 & (~n1273 | n4691));
  assign n2285 = n2252 & n2283 & (n2284 | n2254);
  assign n2286 = (n1021_1 | n3954) & (n2174 | n3952);
  assign n2287 = n2252 & n2286 & (n2176 | n2254);
  assign n2288 = (n2280 | n3894) & (n2287 | n3740);
  assign n2289 = n4369 & (n2285 | n3737);
  assign n2290 = n2288 & n2289 & (n2275 | n2272);
  assign n2291 = (n895 | n3954) & (n2140 | n3952);
  assign n2292 = n2252 & n2291 & (n2142 | n2254);
  assign n2293 = (n974 | n3954) & (n2154 | n3952);
  assign n2294 = n2252 & n2293 & (n2156 | n2254);
  assign n2295 = (n1065 | n3954) & (n2192 | n3952);
  assign n2296 = n2252 & n2295 & (n2194 | n2254);
  assign n2297 = (n1108 | n3954) & (n2197 | n3952);
  assign n2298 = n2252 & n2297 & (n2199 | n2254);
  assign n2299 = (n857 | n3954) & (n2136 | n3952);
  assign n2300 = n2252 & n2299 & (n2138 | n2254);
  assign n2301 = (n1149 | n3954) & (n2208 | n3952);
  assign n2302 = n2252 & n2301 & (n2210 | n2254);
  assign n2303 = (n1189 | n3954) & (n2213 | n3952);
  assign n2304 = n2252 & n2303 & (n2215 | n2254);
  assign n2305 = (n947 | n3954) & (n2150 | n3952);
  assign n2306 = n2252 & n2305 & (n2152 | n2254);
  assign n2307 = (n2300 | n3894) & (n2306 | n3740);
  assign n2308 = n4367 & (n2304 | n3737);
  assign n2309 = n2307 & n2308 & (n2296 | n2272);
  assign n2310 = (n1049 | n3954) & (n2188 | n3952);
  assign n2311 = n2252 & n2310 & (n2190 | n2254);
  assign n2312 = (n1081_1 | n3954) & (n2196 | n3952);
  assign n2313 = (n1081_1 & n4691) | (n4690 & (~n1081_1 | n4691));
  assign n2314 = n2252 & n2312 & (n2313 | n2254);
  assign n2315 = (n821 | n3954) & (n2132 | n3952);
  assign n2316 = n2252 & n2315 & (n2134 | n2254);
  assign n2317 = (n1135 | n3954) & (n2204 | n3952);
  assign n2318 = n2252 & n2317 & (n2206 | n2254);
  assign n2319 = (n1165 | n3954) & (n2212 | n3952);
  assign n2320 = (n1165 & n4691) | (n4690 & (~n1165 | n4691));
  assign n2321 = n2252 & n2319 & (n2320 | n2254);
  assign n2322 = (n922 | n3954) & (n2146 | n3952);
  assign n2323 = n2252 & n2322 & (n2148 | n2254);
  assign n2324 = (n2316 | n3894) & (n2323 | n3740);
  assign n2325 = n4366 & (n2321 | n3737);
  assign n2326 = n2324 & n2325 & (n2311 | n2272);
  assign n2327 = ~Ni34 & (~n882 | n1539);
  assign n2328 = ~Ni34 & (~n966 | n1539);
  assign n2329 = ~Ni34 & (~n1228 | n1539);
  assign n2330 = ~Ni34 & (~n1247 | n1539);
  assign n2331 = ~Ni34 & (~n1001_1 | n1539);
  assign n2332 = ~Ni34 & (~n1266 | n1539);
  assign n2333 = ~Ni34 & (~n1280 | n1539);
  assign n2334 = ~Ni34 & (~n1028 | n1539);
  assign n2335 = ~n3894 & (~n3955 | ~n4355);
  assign n2336 = ~n3743 & (~n3955 | ~n4359);
  assign n2337 = ~Ni34 & (~n1217 | n1539);
  assign n2338 = ~Ni34 & (~n1235 | n1539);
  assign n2339 = ~Ni34 & (~n984 | n1539);
  assign n2340 = ~Ni34 & (~n1259 | n1539);
  assign n2341 = ~Ni34 & (~n1273 | n1539);
  assign n2342 = ~Ni34 & (~n1021_1 | n1539);
  assign n2343 = ~n3894 & (~n3955 | ~n4345);
  assign n2344 = ~n3743 & (~n3955 | ~n4349);
  assign n2345 = n3184 & Pi16;
  assign n2346 = n2345 & (~n3955 | ~n4344);
  assign n2347 = ~Ni34 & (~n895 | n1539);
  assign n2348 = ~Ni34 & (~n974 | n1539);
  assign n2349 = ~Ni34 & (~n1065 | n1539);
  assign n2350 = ~Ni34 & (~n1108 | n1539);
  assign n2351 = ~Ni34 & (~n857 | n1539);
  assign n2352 = ~Ni34 & (~n1149 | n1539);
  assign n2353 = ~Ni34 & (~n1189 | n1539);
  assign n2354 = ~Ni34 & (~n947 | n1539);
  assign n2355 = ~n3894 & (~n3955 | ~n4332);
  assign n2356 = ~n3743 & (~n3955 | ~n4336);
  assign n2357 = ~Ni34 & (~n1049 | n1539);
  assign n2358 = ~Ni34 & (~n1081_1 | n1539);
  assign n2359 = ~Ni34 & (~n821 | n1539);
  assign n2360 = ~Ni34 & (~n1135 | n1539);
  assign n2361 = ~Ni34 & (~n1165 | n1539);
  assign n2362 = ~Ni34 & (~n922 | n1539);
  assign n2363 = ~n3894 & (~n3955 | ~n4322);
  assign n2364 = ~n3743 & (~n3955 | ~n4326);
  assign n2365 = n2345 & (~n3955 | ~n4321);
  assign n2366 = n4371 & (n3944 | (n4368 & n4372));
  assign n2367 = ~Pi15 | n3327;
  assign n2368 = (n2255 | ~n3772) & (n2257 | ~n2345);
  assign n2369 = (~Pi20 & n2290) | (n2273 & (Pi20 | n2290));
  assign n2370 = n2366 & (n2367 | (n2368 & n2369));
  assign n2371 = (~Ni34 | n1919) & n2085;
  assign n2372 = ~Pi25 | n3857;
  assign n2373 = (n2338 | n2372) & (n2330 | n1314);
  assign n2374 = (n2337 | n2372) & (n2329 | n1314);
  assign n2375 = (n2339 | n2372) & (n2331 | n1314);
  assign n2376 = (n2341 | n2372) & (n2333 | n1314);
  assign n2377 = (n2340 | n2372) & (n2332 | n1314);
  assign n2378 = (n2342 | n2372) & (n2334 | n1314);
  assign n2379 = ~n1923 & ~n2328 & (Pi16 | ~n2327);
  assign n2380 = (n2358 | n2372) & (n2350 | n1314);
  assign n2381 = (n2357 | n2372) & (n2349 | n1314);
  assign n2382 = (n2359 | n2372) & (n2351 | n1314);
  assign n2383 = (n2361 | n2372) & (n2353 | n1314);
  assign n2384 = (n2360 | n2372) & (n2352 | n1314);
  assign n2385 = (n2362 | n2372) & (n2354 | n1314);
  assign n2386 = ~n1923 & ~n2348 & (Pi16 | ~n2347);
  assign n2387 = ~n4689 & (~Pi15 | ~n4305 | ~n4307);
  assign n2388 = ~n3659 & (~n3994 | (n2387 & ~n3892));
  assign n2389 = ~Ni35 | Ni30;
  assign n2390 = n1241 & n2389 & (~Ni35 | n1353);
  assign n2391 = Ni32 | n3958;
  assign n2392 = n2390 & (~Pi26 | n2391);
  assign n2393 = n1543 | n3727;
  assign n2394 = Ni35 & (n2393 | ~n3807);
  assign n2395 = ~n2072 & (~n2073 | ~n2403);
  assign n2396 = ~n2395 & (n2394 | (~n2392 & ~n2393));
  assign n2397 = ~n2073 | n2403 | n4702 | n4703;
  assign n2398 = ~n3707 & ~n3896;
  assign n2399 = ~Ni31 | ~Ni36;
  assign n2400 = n891 & n2399 & (Ni30 | ~Ni36);
  assign n2401 = (~Pi27 | n2391) & n2400;
  assign n2402 = ~n4706 & (Ni36 | ~n2393);
  assign n2403 = Ni8 | n3957;
  assign n2404 = n2402 & (n2072 | (n2073 & n2403));
  assign n2405 = ~n2073 | n2403 | n4704 | n4705;
  assign n2406 = ~Ni31 & Ni30;
  assign n2407 = ~n4708 & ~Ni32 & n2406;
  assign n2408 = ~Ni30 & (~n814 | (Ni37 & ~n4708));
  assign n2409 = ~Pi20 | n3961 | n3962;
  assign n2410 = Pi20 | n3959 | n3962;
  assign n2411 = Pi20 | n3959 | n3960;
  assign n2412 = ~Pi20 | n3960 | n3961;
  assign n2413 = n2412 & n2411 & n2409 & n2410;
  assign n2414 = n1216 | (n784 & Ni30);
  assign n2415 = ~n784 & ((Ni37 & n654) | ~n814);
  assign n2416 = ~Ni31 | Ni30;
  assign n2417 = Ni45 & (Ni32 | n2416);
  assign n2418 = ~Ni6 | Ni5;
  assign n2419 = ~Ni32 | Ni30;
  assign n2420 = Ni30 | Ni31;
  assign n2421 = Pi21 | ~Ni32;
  assign n2422 = Pi22 | n3812;
  assign n2423 = n2421 & (~Pi21 | n2422);
  assign n2424 = n2419 & (~n803 | n2420);
  assign n2425 = ~Ni45 & (Ni47 | ~Ni43);
  assign n2426 = Ni41 | Ni42;
  assign n2427 = n2425 & (Ni47 | n2426 | ~n3331);
  assign n2428 = n2425 & n2451;
  assign n2429 = n2518 | Ni40;
  assign n2430 = ~Ni37 | Ni47 | Ni38;
  assign n2431 = n3811 | n3854;
  assign n2432 = n2431 & n2430 & n2428 & n2429;
  assign n2433 = Ni38 | n3811;
  assign n2434 = ~Ni35 | Ni36;
  assign n2435 = n2432 & (n2433 | n2434);
  assign n2436 = n2419 & (~n804 | ~n2435);
  assign n2437 = n2419 & (n2420 | ~n2435);
  assign n2438 = ~n18 | n784;
  assign n2439 = n784 & n2437;
  assign n2440 = n2438 & (n18 | n2439);
  assign n2441 = ~Ni44 & ~Ni43;
  assign n2442 = n2425 & (Ni47 | n2441 | n2426);
  assign n2443 = n2523 | Ni40;
  assign n2444 = n3811 | n3855;
  assign n2445 = n2444 & n2430 & n2428 & n2443;
  assign n2446 = n2445 & (n2433 | n2434);
  assign n2447 = n2419 & (~n804 | ~n2446);
  assign n2448 = n2419 & (n2420 | ~n2446);
  assign n2449 = n784 & n2448;
  assign n2450 = n2438 & (n18 | n2449);
  assign n2451 = ~Ni41 | n3811;
  assign n2452 = n2428 & n2433 & n2430;
  assign n2453 = n2428 & n2430 & (Ni36 | n2452);
  assign n2454 = n2419 & (~n804 | ~n2453);
  assign n2455 = n2419 & (n2420 | ~n2453);
  assign n2456 = n784 & n2455;
  assign n2457 = n2438 & (n18 | n2456);
  assign n2458 = (n2689 | n1702) & (n4404 | n1408);
  assign n2459 = n2447 & n2450;
  assign n2460 = n2423 & n2458 & (n2459 | n914);
  assign n2461 = n2427 | Ni40;
  assign n2462 = n2431 & n2430 & n2425 & n2461;
  assign n2463 = n2462 & (n2433 | n2434);
  assign n2464 = n2419 & (~n804 | ~n2463);
  assign n2465 = n2419 & (n2420 | ~n2463);
  assign n2466 = n784 & n2465;
  assign n2467 = n2438 & (n18 | n2466);
  assign n2468 = n2442 | Ni40;
  assign n2469 = n2444 & n2430 & n2425 & n2468;
  assign n2470 = n2469 & (n2433 | n2434);
  assign n2471 = n2419 & (~n804 | ~n2470);
  assign n2472 = n2419 & (n2420 | ~n2470);
  assign n2473 = n784 & n2472;
  assign n2474 = n2438 & (n18 | n2473);
  assign n2475 = n2425 & n2433 & n2430;
  assign n2476 = n2425 & n2430 & (Ni36 | n2475);
  assign n2477 = n2419 & (~n804 | ~n2476);
  assign n2478 = n2419 & (n2420 | ~n2476);
  assign n2479 = n784 & n2478;
  assign n2480 = n2438 & (n18 | n2479);
  assign n2481 = (n2690 | n1702) & (n4405 | n1408);
  assign n2482 = n2471 & n2474;
  assign n2483 = n2423 & n2481 & (n2482 | n914);
  assign n2484 = n2432 & (n2433 | ~n2530);
  assign n2485 = n2419 & (~n804 | ~n2484);
  assign n2486 = n2419 & (n2420 | ~n2484);
  assign n2487 = n784 & n2486;
  assign n2488 = n2438 & (n18 | n2487);
  assign n2489 = n2445 & (n2433 | ~n2530);
  assign n2490 = n2419 & (~n804 | ~n2489);
  assign n2491 = n2419 & (n2420 | ~n2489);
  assign n2492 = n784 & n2491;
  assign n2493 = n2438 & (n18 | n2492);
  assign n2494 = n2419 & (~n804 | ~n2452);
  assign n2495 = n2419 & (n2420 | ~n2452);
  assign n2496 = n784 & n2495;
  assign n2497 = n2438 & (n18 | n2496);
  assign n2498 = (n2666 | n1702) & (n4414 | n1408);
  assign n2499 = n2490 & n2493;
  assign n2500 = n2423 & n2498 & (n2499 | n914);
  assign n2501 = n2462 & (n2433 | ~n2530);
  assign n2502 = n2419 & (~n804 | ~n2501);
  assign n2503 = n2419 & (n2420 | ~n2501);
  assign n2504 = n784 & n2503;
  assign n2505 = n2438 & (n18 | n2504);
  assign n2506 = n2469 & (n2433 | ~n2530);
  assign n2507 = n2419 & (~n804 | ~n2506);
  assign n2508 = n2419 & (n2420 | ~n2506);
  assign n2509 = n784 & n2508;
  assign n2510 = n2438 & (n18 | n2509);
  assign n2511 = n2419 & (~n804 | ~n2475);
  assign n2512 = n2419 & (n2420 | ~n2475);
  assign n2513 = n784 & n2512;
  assign n2514 = n2438 & (n18 | n2513);
  assign n2515 = (n2667 | n1702) & (n4415 | n1408);
  assign n2516 = n2507 & n2510;
  assign n2517 = n2423 & n2515 & (n2516 | n914);
  assign n2518 = n2451 & n2427;
  assign n2519 = n2419 & (~n804 | ~n3963);
  assign n2520 = n2419 & (n2420 | ~n3963);
  assign n2521 = n784 & n2520;
  assign n2522 = n2438 & (n18 | n2521);
  assign n2523 = n2451 & n2442;
  assign n2524 = n2419 & (~n804 | ~n3964);
  assign n2525 = n2419 & (n2420 | ~n3964);
  assign n2526 = n784 & n2525;
  assign n2527 = n2438 & (n18 | n2526);
  assign n2528 = n2518 | ~Ni40;
  assign n2529 = n2431 & n2430 & n2428 & n2528;
  assign n2530 = Ni35 | Ni36;
  assign n2531 = n2529 & (n2433 | n2530);
  assign n2532 = n2419 & (~n804 | ~n2531);
  assign n2533 = n2419 & (n2420 | ~n2531);
  assign n2534 = n784 & n2533;
  assign n2535 = n2438 & (n18 | n2534);
  assign n2536 = n2523 | ~Ni40;
  assign n2537 = n2444 & n2430 & n2428 & n2536;
  assign n2538 = n2537 & (n2433 | n2530);
  assign n2539 = n2419 & (~n804 | ~n2538);
  assign n2540 = n2419 & (n2420 | ~n2538);
  assign n2541 = n784 & n2540;
  assign n2542 = n2438 & (n18 | n2541);
  assign n2543 = (n4408 | n3893) & (n2718 | n2109);
  assign n2544 = n2423 & (n2721 | n914);
  assign n2545 = n2519 & n2522;
  assign n2546 = n2543 & n2544 & (n2545 | n1408);
  assign n2547 = n2419 & (~n804 | ~n3965);
  assign n2548 = n2419 & (n2420 | ~n3965);
  assign n2549 = n784 & n2548;
  assign n2550 = n2438 & (n18 | n2549);
  assign n2551 = n2419 & (~n804 | ~n3966);
  assign n2552 = n2419 & (n2420 | ~n3966);
  assign n2553 = n784 & n2552;
  assign n2554 = n2438 & (n18 | n2553);
  assign n2555 = n2427 | ~Ni40;
  assign n2556 = n2431 & n2430 & n2425 & n2555;
  assign n2557 = n2556 & (n2433 | n2530);
  assign n2558 = n2419 & (~n804 | ~n2557);
  assign n2559 = n2419 & (n2420 | ~n2557);
  assign n2560 = n784 & n2559;
  assign n2561 = n2438 & (n18 | n2560);
  assign n2562 = n2442 | ~Ni40;
  assign n2563 = n2444 & n2430 & n2425 & n2562;
  assign n2564 = n2563 & (n2433 | n2530);
  assign n2565 = n2419 & (~n804 | ~n2564);
  assign n2566 = n2419 & (n2420 | ~n2564);
  assign n2567 = n784 & n2566;
  assign n2568 = n2438 & (n18 | n2567);
  assign n2569 = (n4411 | n3893) & (n2706 | n2109);
  assign n2570 = n2423 & (n2710 | n914);
  assign n2571 = n2547 & n2550;
  assign n2572 = n2569 & n2570 & (n2571 | n1408);
  assign n2573 = ~n3963 | ~n4768;
  assign n2574 = n2419 & (~n804 | n2573);
  assign n2575 = n2419 & (n2420 | n2573);
  assign n2576 = n784 & n2575;
  assign n2577 = n2438 & (n18 | n2576);
  assign n2578 = ~n3964 | ~n4768;
  assign n2579 = n2419 & (~n804 | n2578);
  assign n2580 = n2419 & (n2420 | n2578);
  assign n2581 = n784 & n2580;
  assign n2582 = n2438 & (n18 | n2581);
  assign n2583 = n2529 & (n2433 | ~n2434);
  assign n2584 = n2419 & (~n804 | ~n2583);
  assign n2585 = n2419 & (n2420 | ~n2583);
  assign n2586 = n784 & n2585;
  assign n2587 = n2438 & (n18 | n2586);
  assign n2588 = n2537 & (n2433 | ~n2434);
  assign n2589 = n2419 & (~n804 | ~n2588);
  assign n2590 = n2419 & (n2420 | ~n2588);
  assign n2591 = n784 & n2590;
  assign n2592 = n2438 & (n18 | n2591);
  assign n2593 = (n4418 | n3893) & (n2740 | n2109);
  assign n2594 = n2423 & (n2743 | n914);
  assign n2595 = n2574 & n2577;
  assign n2596 = n2593 & n2594 & (n2595 | n1408);
  assign n2597 = ~n3965 | ~n4768;
  assign n2598 = n2419 & (~n804 | n2597);
  assign n2599 = n2419 & (n2420 | n2597);
  assign n2600 = n784 & n2599;
  assign n2601 = n2438 & (n18 | n2600);
  assign n2602 = ~n3966 | ~n4768;
  assign n2603 = n2419 & (~n804 | n2602);
  assign n2604 = n2419 & (n2420 | n2602);
  assign n2605 = n784 & n2604;
  assign n2606 = n2438 & (n18 | n2605);
  assign n2607 = n2556 & (n2433 | ~n2434);
  assign n2608 = n2419 & (~n804 | ~n2607);
  assign n2609 = n2419 & (n2420 | ~n2607);
  assign n2610 = n784 & n2609;
  assign n2611 = n2438 & (n18 | n2610);
  assign n2612 = n2563 & (n2433 | ~n2434);
  assign n2613 = n2419 & (~n804 | ~n2612);
  assign n2614 = n2419 & (n2420 | ~n2612);
  assign n2615 = n784 & n2614;
  assign n2616 = n2438 & (n18 | n2615);
  assign n2617 = (n4421 | n3893) & (n2729 | n2109);
  assign n2618 = n2423 & (n2732 | n914);
  assign n2619 = n2598 & n2601;
  assign n2620 = n2617 & n2618 & (n2619 | n1408);
  assign n2621 = n2641 & n2423;
  assign n2622 = (n1448 | n2621) & (n1446 | ~n3998);
  assign n2623 = n802 & (~Pi27 | ~Ni32) & n2419;
  assign n2624 = n4709 & (Pi22 | ~Pi21 | n3821);
  assign n2625 = (~Pi26 | n3037) & n3817;
  assign n2626 = n2624 & (n2625 | n2254);
  assign n2627 = n802 & n2419 & (Pi27 | ~Ni32);
  assign n2628 = (n2627 & (~Pi21 | ~n3999)) | (Pi21 & ~n3999);
  assign n2629 = n3813 & (Pi27 | n3037);
  assign n2630 = n2628 & (n2629 | n2254);
  assign n2631 = (n2621 | n1452) & (n2630 | n3696);
  assign n2632 = ~Ni12 | n3912;
  assign n2633 = n2622 & n2631 & (n2626 | n2632);
  assign n2634 = ~n4711 & (Pi22 | ~Pi21 | n3826);
  assign n2635 = n3817 & (Pi26 | n3037);
  assign n2636 = n2634 & (n2635 | n2254);
  assign n2637 = Pi21 & ~n2422 & (~Pi24 | ~n813);
  assign n2638 = Pi21 | n3822;
  assign n2639 = ~n2637 & (Pi24 | n2421) & n2638;
  assign n2640 = n3825 | n2254;
  assign n2641 = n3037 | n2254;
  assign n2642 = n2640 & n2639 & (Pi24 | n2641);
  assign n2643 = Pi22 | ~Pi21;
  assign n2644 = n2640 & n2638 & (n813 | n2643);
  assign n2645 = n3823 | n2643;
  assign n2646 = n2649 & (~Pi27 | n3822);
  assign n2647 = n3824 & (~Pi27 | n3825);
  assign n2648 = n2645 & n2646 & (n2647 | n2254);
  assign n2649 = n2419 & n801;
  assign n2650 = (n2750 | ~n4005) & (n3912 | ~n4006);
  assign n2651 = n2650 & (n2642 | ~Ni13);
  assign n2652 = n812 & n2494 & (n18 | n2495);
  assign n2653 = n812 & n2511 & (n18 | n2512);
  assign n2654 = n812 & n2584 & (n18 | n2585);
  assign n2655 = n812 & n2589 & (n18 | n2590);
  assign n2656 = n812 & n2574 & (n18 | n2575);
  assign n2657 = n812 & n2579 & (n18 | n2580);
  assign n2658 = n812 & n2485 & (n18 | n2486);
  assign n2659 = n812 & n2490 & (n18 | n2491);
  assign n2660 = n812 & n2608 & (n18 | n2609);
  assign n2661 = n812 & n2613 & (n18 | n2614);
  assign n2662 = n812 & n2598 & (n18 | n2599);
  assign n2663 = n812 & n2603 & (n18 | n2604);
  assign n2664 = n812 & n2502 & (n18 | n2503);
  assign n2665 = n812 & n2507 & (n18 | n2508);
  assign n2666 = n2494 & n2497;
  assign n2667 = n2511 & n2514;
  assign n2668 = (n2666 | n1495) & (n2667 | n1497);
  assign n2669 = ~n3740 & (~n4553 | ~n4554);
  assign n2670 = ~n2272 & (~n4555 | ~n4556);
  assign n2671 = n2639 & (n3737 | (n4562 & n4561));
  assign n2672 = n4565 & (n3743 | (n4560 & n4559));
  assign n2673 = n4563 & n4564 & (Pi24 | n2668);
  assign n2674 = n2673 & n2671 & n2672;
  assign n2675 = n812 & n2454 & (n18 | n2455);
  assign n2676 = n812 & n2477 & (n18 | n2478);
  assign n2677 = n812 & n2532 & (n18 | n2533);
  assign n2678 = n812 & n2539 & (n18 | n2540);
  assign n2679 = n812 & n2519 & (n18 | n2520);
  assign n2680 = n812 & n2524 & (n18 | n2525);
  assign n2681 = n812 & n2436 & (n18 | n2437);
  assign n2682 = n812 & n2447 & (n18 | n2448);
  assign n2683 = n812 & n2558 & (n18 | n2559);
  assign n2684 = n812 & n2565 & (n18 | n2566);
  assign n2685 = n812 & n2547 & (n18 | n2548);
  assign n2686 = n812 & n2551 & (n18 | n2552);
  assign n2687 = n812 & n2464 & (n18 | n2465);
  assign n2688 = n812 & n2471 & (n18 | n2472);
  assign n2689 = n2454 & n2457;
  assign n2690 = n2477 & n2480;
  assign n2691 = (n2689 | n1495) & (n2690 | n1497);
  assign n2692 = ~n3740 & (~n4535 | ~n4536);
  assign n2693 = ~n2272 & (~n4537 | ~n4538);
  assign n2694 = ~n3944 & (~n4547 | ~n4549 | ~n4550);
  assign n2695 = ~n2694 & (n2642 | (n1448 & n1542));
  assign n2696 = (n2651 | n3919) & (n3677 | ~n4007);
  assign n2697 = n2695 & n2696 & (n2674 | n2367);
  assign n2698 = Pi21 & ~n2422 & (n788 | ~n813);
  assign n2699 = n2638 & (~n788 | n2421) & ~n2698;
  assign n2700 = n2640 & n2699 & (~n788 | n2641);
  assign n2701 = ~n2643 & (~n4508 | (Pi24 & ~n3821));
  assign n2702 = ~n2254 & (~n4509 | (Pi24 & ~n2625));
  assign n2703 = ~Pi21 & (~n4510 | (Pi24 & ~n3818));
  assign n2704 = n1542 & (n1543 | ~n2750);
  assign n2705 = n4523 & (n4411 | n3936);
  assign n2706 = n2565 & n2568;
  assign n2707 = ~n788 | n3859;
  assign n2708 = n2699 & n2705 & (n2706 | n2707);
  assign n2709 = n4522 & (n2571 | n3936);
  assign n2710 = n2551 & n2554;
  assign n2711 = n2699 & n2709 & (n2710 | n2707);
  assign n2712 = n4521 & (n4405 | n3936);
  assign n2713 = n2699 & n2712 & (n2482 | n2707);
  assign n2714 = (n2713 | n3864) & (n2711 | n3867);
  assign n2715 = n4524 & (n2690 | n3934);
  assign n2716 = n2714 & n2715 & (n2708 | n1322);
  assign n2717 = n4514 & (n4408 | n3936);
  assign n2718 = n2539 & n2542;
  assign n2719 = n2699 & n2717 & (n2718 | n2707);
  assign n2720 = n4513 & (n2545 | n3936);
  assign n2721 = n2524 & n2527;
  assign n2722 = n2699 & n2720 & (n2721 | n2707);
  assign n2723 = n4512 & (n4404 | n3936);
  assign n2724 = n2699 & n2723 & (n2459 | n2707);
  assign n2725 = (n2724 | n3864) & (n2722 | n3867);
  assign n2726 = n4516 & (n2689 | n3934);
  assign n2727 = n2725 & n2726 & (n2719 | n1322);
  assign n2728 = n4527 & (n4421 | n3936);
  assign n2729 = n2613 & n2616;
  assign n2730 = n2699 & n2728 & (n2729 | n2707);
  assign n2731 = n4526 & (n2619 | n3936);
  assign n2732 = n2603 & n2606;
  assign n2733 = n2699 & n2731 & (n2732 | n2707);
  assign n2734 = n4525 & (n4415 | n3936);
  assign n2735 = n2699 & n2734 & (n2516 | n2707);
  assign n2736 = (n2735 | n3864) & (n2733 | n3867);
  assign n2737 = n4528 & n4515 & (n2667 | n3934);
  assign n2738 = n2736 & n2737 & (n2730 | n1322);
  assign n2739 = n4519 & (n4418 | n3936);
  assign n2740 = n2589 & n2592;
  assign n2741 = n2699 & n2739 & (n2740 | n2707);
  assign n2742 = n4518 & (n2595 | n3936);
  assign n2743 = n2579 & n2582;
  assign n2744 = n2699 & n2742 & (n2743 | n2707);
  assign n2745 = n4517 & (n4414 | n3936);
  assign n2746 = n2699 & n2745 & (n2499 | n2707);
  assign n2747 = (n2746 | n3864) & (n2744 | n3867);
  assign n2748 = n4520 & (n2666 | n3934);
  assign n2749 = n2747 & n2748 & (n2741 | n1322);
  assign n2750 = ~Ni14 | Ni13;
  assign n2751 = n1545 & ~n2700 & (~n2636 | n2750);
  assign n2752 = ~n3919 & (~n4511 | (~n2700 & Ni13));
  assign n2753 = Pi21 & ~n2422 & (n795 | ~n813);
  assign n2754 = n2638 & (~n795 | n2421) & ~n2753;
  assign n2755 = n2640 & n2754 & (~n795 | n2641);
  assign n2756 = n4578 & (n4411 | n3948);
  assign n2757 = ~n795 | n3859;
  assign n2758 = n2754 & n2756 & (n2706 | n2757);
  assign n2759 = n4577 & (n2571 | n3948);
  assign n2760 = n2754 & n2759 & (n2710 | n2757);
  assign n2761 = n4576 & (n4405 | n3948);
  assign n2762 = n2754 & n2761 & (n2482 | n2757);
  assign n2763 = (n2762 | n3864) & (n2760 | n3867);
  assign n2764 = n4579 & (n2690 | n3946);
  assign n2765 = n2763 & n2764 & (n2758 | n1322);
  assign n2766 = n4569 & (n4408 | n3948);
  assign n2767 = n2754 & n2766 & (n2718 | n2757);
  assign n2768 = n4568 & (n2545 | n3948);
  assign n2769 = n2754 & n2768 & (n2721 | n2757);
  assign n2770 = n4567 & (n4404 | n3948);
  assign n2771 = n2754 & n2770 & (n2459 | n2757);
  assign n2772 = (n2771 | n3864) & (n2769 | n3867);
  assign n2773 = n4571 & (n2689 | n3946);
  assign n2774 = n2772 & n2773 & (n2767 | n1322);
  assign n2775 = n4582 & (n4421 | n3948);
  assign n2776 = n2754 & n2775 & (n2729 | n2757);
  assign n2777 = n4581 & (n2619 | n3948);
  assign n2778 = n2754 & n2777 & (n2732 | n2757);
  assign n2779 = n4580 & (n4415 | n3948);
  assign n2780 = n2754 & n2779 & (n2516 | n2757);
  assign n2781 = (n2780 | n3864) & (n2778 | n3867);
  assign n2782 = n4583 & n4570 & (n2667 | n3946);
  assign n2783 = n2781 & n2782 & (n2776 | n1322);
  assign n2784 = n4574 & (n4418 | n3948);
  assign n2785 = n2754 & n2784 & (n2740 | n2757);
  assign n2786 = n4573 & (n2595 | n3948);
  assign n2787 = n2754 & n2786 & (n2743 | n2757);
  assign n2788 = n4572 & (n4414 | n3948);
  assign n2789 = n2754 & n2788 & (n2499 | n2757);
  assign n2790 = (n2789 | n3864) & (n2787 | n3867);
  assign n2791 = n4575 & (n2666 | n3946);
  assign n2792 = n2790 & n2791 & (n2785 | n1322);
  assign n2793 = n1545 & ~n2755 & (~n2636 | n2750);
  assign n2794 = ~n3919 & ((Ni13 & ~n2755) | ~n4566);
  assign n2795 = n2419 & (~n805 | ~n2435);
  assign n2796 = n2419 & (~n805 | ~n2446);
  assign n2797 = n2419 & (~n805 | ~n2453);
  assign n2798 = (n4398 | n1702) & (n2918 | n1408);
  assign n2799 = n2796 & n2450;
  assign n2800 = n2423 & n2798 & (n2799 | n914);
  assign n2801 = n2419 & (~n805 | ~n2463);
  assign n2802 = n2419 & (~n805 | ~n2470);
  assign n2803 = n2419 & (~n805 | ~n2476);
  assign n2804 = (n4400 | n1702) & (n2890 | n1408);
  assign n2805 = n2802 & n2474;
  assign n2806 = n2423 & n2804 & (n2805 | n914);
  assign n2807 = n2419 & (~n805 | ~n2484);
  assign n2808 = n2419 & (~n805 | ~n2489);
  assign n2809 = n2419 & (~n805 | ~n2452);
  assign n2810 = (n4399 | n1702) & (n2974 | n1408);
  assign n2811 = n2808 & n2493;
  assign n2812 = n2423 & n2810 & (n2811 | n914);
  assign n2813 = n2419 & (~n805 | ~n2501);
  assign n2814 = n2419 & (~n805 | ~n2506);
  assign n2815 = n2419 & (~n805 | ~n2475);
  assign n2816 = (n4401 | n1702) & (n2946 | n1408);
  assign n2817 = n2814 & n2510;
  assign n2818 = n2423 & n2816 & (n2817 | n914);
  assign n2819 = n2419 & (~n805 | ~n3963);
  assign n2820 = n2419 & (~n805 | ~n3964);
  assign n2821 = n2419 & (~n805 | ~n2531);
  assign n2822 = n2419 & (~n805 | ~n2538);
  assign n2823 = (n2903 | n3893) & (n4388 | n2109);
  assign n2824 = n2423 & (n4389 | n914);
  assign n2825 = n2819 & n2522;
  assign n2826 = n2823 & n2824 & (n2825 | n1408);
  assign n2827 = n2419 & (~n805 | ~n3965);
  assign n2828 = n2419 & (~n805 | ~n3966);
  assign n2829 = n2419 & (~n805 | ~n2557);
  assign n2830 = n2419 & (~n805 | ~n2564);
  assign n2831 = (n2875 | n3893) & (n4392 | n2109);
  assign n2832 = n2423 & (n4393 | n914);
  assign n2833 = n2827 & n2550;
  assign n2834 = n2831 & n2832 & (n2833 | n1408);
  assign n2835 = n2419 & (~n805 | n2573);
  assign n2836 = n2419 & (~n805 | n2578);
  assign n2837 = n2419 & (~n805 | ~n2583);
  assign n2838 = n2419 & (~n805 | ~n2588);
  assign n2839 = (n2959 | n3893) & (n4390 | n2109);
  assign n2840 = n2423 & (n4391 | n914);
  assign n2841 = n2835 & n2577;
  assign n2842 = n2839 & n2840 & (n2841 | n1408);
  assign n2843 = n2419 & (~n805 | n2597);
  assign n2844 = n2419 & (~n805 | n2602);
  assign n2845 = n2419 & (~n805 | ~n2607);
  assign n2846 = n2419 & (~n805 | ~n2612);
  assign n2847 = (n2931 | n3893) & (n4394 | n2109);
  assign n2848 = n2423 & (n4395 | n914);
  assign n2849 = n2843 & n2601;
  assign n2850 = n2847 & n2848 & (n2849 | n1408);
  assign n2851 = (Pi20 & n2449) | (n2439 & (~Pi20 | n2449));
  assign n2852 = (n2851 | n1701) & (n2456 | n1702);
  assign n2853 = (Pi20 & n2473) | (n2466 & (~Pi20 | n2473));
  assign n2854 = (n2853 | n1701) & (n2479 | n1702);
  assign n2855 = (Pi20 & n2509) | (n2504 & (~Pi20 | n2509));
  assign n2856 = (n2855 | n1701) & (n2513 | n1702);
  assign n2857 = (Pi20 & n2526) | (n2521 & (~Pi20 | n2526));
  assign n2858 = (Pi20 & n2541) | (n2534 & (~Pi20 | n2541));
  assign n2859 = (n2857 | n1701) & (n2858 | n1702);
  assign n2860 = (Pi20 & n2553) | (n2549 & (~Pi20 | n2553));
  assign n2861 = (Pi20 & n2567) | (n2560 & (~Pi20 | n2567));
  assign n2862 = (n2860 | n1701) & (n2861 | n1702);
  assign n2863 = (Pi20 & n2605) | (n2600 & (~Pi20 | n2605));
  assign n2864 = (Pi20 & n2615) | (n2610 & (~Pi20 | n2615));
  assign n2865 = (n2863 | n1701) & (n2864 | n1702);
  assign n2866 = n1446 | n4721 | n4722;
  assign n2867 = ~n4720 & (Pi17 | (n4396 & n4397));
  assign n2868 = n2866 & (n2867 | n1448);
  assign n2869 = n802 & n2559;
  assign n2870 = n802 & n2829 & (n18 | n2869);
  assign n2871 = n802 & n2566;
  assign n2872 = n802 & n2830 & (n18 | n2871);
  assign n2873 = (n2870 | n3915) & (n2872 | n3916);
  assign n2874 = n2624 & (n4392 | n3917);
  assign n2875 = n2829 & n2561;
  assign n2876 = n2873 & n2874 & (n2875 | n1729);
  assign n2877 = n802 & n2548;
  assign n2878 = n802 & n2827 & (n18 | n2877);
  assign n2879 = n802 & n2552;
  assign n2880 = n802 & n2828 & (n18 | n2879);
  assign n2881 = (n2878 | n3915) & (n2880 | n3916);
  assign n2882 = n2624 & (n4393 | n3917);
  assign n2883 = n2881 & n2882 & (n2833 | n1729);
  assign n2884 = n802 & n2465;
  assign n2885 = n802 & n2801 & (n18 | n2884);
  assign n2886 = n802 & n2472;
  assign n2887 = n802 & n2802 & (n18 | n2886);
  assign n2888 = (n2885 | n3915) & (n2887 | n3916);
  assign n2889 = n2624 & (n2805 | n3917);
  assign n2890 = n2801 & n2467;
  assign n2891 = n2888 & n2889 & (n2890 | n1729);
  assign n2892 = n802 & n2478;
  assign n2893 = n802 & n2803 & (n18 | n2892);
  assign n2894 = (n2891 | n3864) & (n2883 | n3867);
  assign n2895 = n4503 & n4501 & (n4400 | n3914);
  assign n2896 = n2894 & n2895 & (n2876 | n1322);
  assign n2897 = n802 & n2533;
  assign n2898 = n802 & n2821 & (n18 | n2897);
  assign n2899 = n802 & n2540;
  assign n2900 = n802 & n2822 & (n18 | n2899);
  assign n2901 = (n2898 | n3915) & (n2900 | n3916);
  assign n2902 = n2624 & (n4388 | n3917);
  assign n2903 = n2821 & n2535;
  assign n2904 = n2901 & n2902 & (n2903 | n1729);
  assign n2905 = n802 & n2520;
  assign n2906 = n802 & n2819 & (n18 | n2905);
  assign n2907 = n802 & n2525;
  assign n2908 = n802 & n2820 & (n18 | n2907);
  assign n2909 = (n2906 | n3915) & (n2908 | n3916);
  assign n2910 = n2624 & (n4389 | n3917);
  assign n2911 = n2909 & n2910 & (n2825 | n1729);
  assign n2912 = n802 & n2437;
  assign n2913 = n802 & n2795 & (n18 | n2912);
  assign n2914 = n802 & n2448;
  assign n2915 = n802 & n2796 & (n18 | n2914);
  assign n2916 = (n2913 | n3915) & (n2915 | n3916);
  assign n2917 = n2624 & (n2799 | n3917);
  assign n2918 = n2795 & n2440;
  assign n2919 = n2916 & n2917 & (n2918 | n1729);
  assign n2920 = n802 & n2455;
  assign n2921 = n802 & n2797 & (n18 | n2920);
  assign n2922 = (n2919 | n3864) & (n2911 | n3867);
  assign n2923 = n4500 & n4501 & (n4398 | n3914);
  assign n2924 = n2922 & n2923 & (n2904 | n1322);
  assign n2925 = n802 & n2609;
  assign n2926 = n802 & n2845 & (n18 | n2925);
  assign n2927 = n802 & n2614;
  assign n2928 = n802 & n2846 & (n18 | n2927);
  assign n2929 = (n2926 | n3915) & (n2928 | n3916);
  assign n2930 = n2624 & (n4394 | n3917);
  assign n2931 = n2845 & n2611;
  assign n2932 = n2929 & n2930 & (n2931 | n1729);
  assign n2933 = n802 & n2599;
  assign n2934 = n802 & n2843 & (n18 | n2933);
  assign n2935 = n802 & n2604;
  assign n2936 = n802 & n2844 & (n18 | n2935);
  assign n2937 = (n2934 | n3915) & (n2936 | n3916);
  assign n2938 = n2624 & (n4395 | n3917);
  assign n2939 = n2937 & n2938 & (n2849 | n1729);
  assign n2940 = n802 & n2503;
  assign n2941 = n802 & n2813 & (n18 | n2940);
  assign n2942 = n802 & n2508;
  assign n2943 = n802 & n2814 & (n18 | n2942);
  assign n2944 = (n2941 | n3915) & (n2943 | n3916);
  assign n2945 = n2624 & (n2817 | n3917);
  assign n2946 = n2813 & n2505;
  assign n2947 = n2944 & n2945 & (n2946 | n1729);
  assign n2948 = n802 & n2512;
  assign n2949 = n802 & n2815 & (n18 | n2948);
  assign n2950 = (n2947 | n3864) & (n2939 | n3867);
  assign n2951 = n4504 & n4501 & (n4401 | n3914);
  assign n2952 = n2950 & n2951 & (n2932 | n1322);
  assign n2953 = n802 & n2585;
  assign n2954 = n802 & n2837 & (n18 | n2953);
  assign n2955 = n802 & n2590;
  assign n2956 = n802 & n2838 & (n18 | n2955);
  assign n2957 = (n2954 | n3915) & (n2956 | n3916);
  assign n2958 = n2624 & (n4390 | n3917);
  assign n2959 = n2837 & n2587;
  assign n2960 = n2957 & n2958 & (n2959 | n1729);
  assign n2961 = n802 & n2575;
  assign n2962 = n802 & n2835 & (n18 | n2961);
  assign n2963 = n802 & n2580;
  assign n2964 = n802 & n2836 & (n18 | n2963);
  assign n2965 = (n2962 | n3915) & (n2964 | n3916);
  assign n2966 = n2624 & (n4391 | n3917);
  assign n2967 = n2965 & n2966 & (n2841 | n1729);
  assign n2968 = n802 & n2486;
  assign n2969 = n802 & n2807 & (n18 | n2968);
  assign n2970 = n802 & n2491;
  assign n2971 = n802 & n2808 & (n18 | n2970);
  assign n2972 = (n2969 | n3915) & (n2971 | n3916);
  assign n2973 = n2624 & (n2811 | n3917);
  assign n2974 = n2807 & n2488;
  assign n2975 = n2972 & n2973 & (n2974 | n1729);
  assign n2976 = n802 & n2495;
  assign n2977 = n802 & n2809 & (n18 | n2976);
  assign n2978 = (n2975 | n3864) & (n2967 | n3867);
  assign n2979 = n4502 & n4501 & (n4399 | n3914);
  assign n2980 = n2978 & n2979 & (n2960 | n1322);
  assign n2981 = ~n2272 & (~n4485 | ~n4486);
  assign n2982 = ~n2272 & (~n4466 | ~n4467);
  assign n2983 = n3696 | n4717 | n4719;
  assign n2984 = n2868 & (n2632 | (n4506 & n4505));
  assign n2985 = n2983 & n2984 & (n2867 | n1452);
  assign n2986 = (n2870 | n3901) & (n2872 | n3902);
  assign n2987 = n2634 & (n4392 | n3903);
  assign n2988 = n2986 & n2987 & (n2875 | n1868);
  assign n2989 = (n2878 | n3901) & (n2880 | n3902);
  assign n2990 = n2634 & (n4393 | n3903);
  assign n2991 = n2989 & n2990 & (n2833 | n1868);
  assign n2992 = (n2885 | n3901) & (n2887 | n3902);
  assign n2993 = n2634 & (n2805 | n3903);
  assign n2994 = n2992 & n2993 & (n2890 | n1868);
  assign n2995 = (n2994 | n3864) & (n2991 | n3867);
  assign n2996 = n4460 & n4458 & (n4400 | n3900);
  assign n2997 = n2995 & n2996 & (n2988 | n1322);
  assign n2998 = (n2898 | n3901) & (n2900 | n3902);
  assign n2999 = n2634 & (n4388 | n3903);
  assign n3000 = n2998 & n2999 & (n2903 | n1868);
  assign n3001 = (n2906 | n3901) & (n2908 | n3902);
  assign n3002 = n2634 & (n4389 | n3903);
  assign n3003 = n3001 & n3002 & (n2825 | n1868);
  assign n3004 = (n2913 | n3901) & (n2915 | n3902);
  assign n3005 = n2634 & (n2799 | n3903);
  assign n3006 = n3004 & n3005 & (n2918 | n1868);
  assign n3007 = (n3006 | n3864) & (n3003 | n3867);
  assign n3008 = n4457 & n4458 & (n4398 | n3900);
  assign n3009 = n3007 & n3008 & (n3000 | n1322);
  assign n3010 = (n2926 | n3901) & (n2928 | n3902);
  assign n3011 = n2634 & (n4394 | n3903);
  assign n3012 = n3010 & n3011 & (n2931 | n1868);
  assign n3013 = (n2934 | n3901) & (n2936 | n3902);
  assign n3014 = n2634 & (n4395 | n3903);
  assign n3015 = n3013 & n3014 & (n2849 | n1868);
  assign n3016 = (n2941 | n3901) & (n2943 | n3902);
  assign n3017 = n2634 & (n2817 | n3903);
  assign n3018 = n3016 & n3017 & (n2946 | n1868);
  assign n3019 = (n3018 | n3864) & (n3015 | n3867);
  assign n3020 = n4461 & n4458 & (n4401 | n3900);
  assign n3021 = n3019 & n3020 & (n3012 | n1322);
  assign n3022 = (n2954 | n3901) & (n2956 | n3902);
  assign n3023 = n2634 & (n4390 | n3903);
  assign n3024 = n3022 & n3023 & (n2959 | n1868);
  assign n3025 = (n2962 | n3901) & (n2964 | n3902);
  assign n3026 = n2634 & (n4391 | n3903);
  assign n3027 = n3025 & n3026 & (n2841 | n1868);
  assign n3028 = (n2969 | n3901) & (n2971 | n3902);
  assign n3029 = n2634 & (n2811 | n3903);
  assign n3030 = n3028 & n3029 & (n2974 | n1868);
  assign n3031 = (n3030 | n3864) & (n3027 | n3867);
  assign n3032 = n4459 & n4458 & (n4399 | n3900);
  assign n3033 = n3031 & n3032 & (n3024 | n1322);
  assign n3034 = (n2997 | n3884) & (n3021 | n3891);
  assign n3035 = (n3009 | n3870) & (n3033 | n3877);
  assign n3036 = n3034 & n3035;
  assign n3037 = n784 & n2424;
  assign n3038 = n2423 & (n3037 | n1919);
  assign n3039 = n3038 & (n1929 | (n4387 & n4385));
  assign n3040 = n2496 & (~Pi16 | n2513);
  assign n3041 = n3039 & (n3040 | n1923);
  assign n3042 = n3038 & (n1929 | (n4383 & n4381));
  assign n3043 = n2456 & (~Pi16 | n2479);
  assign n3044 = n3042 & (n3043 | n1923);
  assign n3045 = (n4414 | n3858) & (n2499 | n3860);
  assign n3046 = (Pi20 & n2492) | (n2487 & (~Pi20 | n2492));
  assign n3047 = n3045 & (n3046 | n1929);
  assign n3048 = ~n3740 & ((~n1929 & ~n2855) | ~n4416);
  assign n3049 = ~n2272 & (~n4417 | (~n1929 & ~n3094));
  assign n3050 = ~n3895 & ((~n1929 & ~n3091) | ~n4419);
  assign n3051 = ~n3743 & ((~n1929 & ~n2863) | ~n4420);
  assign n3052 = ~n3737 & ((~n1929 & ~n2864) | ~n4422);
  assign n3053 = (n4404 | n3858) & (n2459 | n3860);
  assign n3054 = n3053 & (n2851 | n1929);
  assign n3055 = ~n3740 & ((~n1929 & ~n2853) | ~n4406);
  assign n3056 = ~n2272 & (~n4407 | (~n1929 & ~n2857));
  assign n3057 = ~n3895 & ((~n1929 & ~n2858) | ~n4409);
  assign n3058 = ~n3743 & ((~n1929 & ~n2860) | ~n4410);
  assign n3059 = ~n3737 & ((~n1929 & ~n2861) | ~n4412);
  assign n3060 = (~Pi15 & n3044) | (n3041 & (Pi15 | n3044));
  assign n3061 = (n1448 | n3060) & (n1446 | ~n3997);
  assign n3062 = n2634 & (n2635 | n1919);
  assign n3063 = (n2869 | n3931) & (n2871 | n3932);
  assign n3064 = n3062 & n3063 & (n2861 | n1948);
  assign n3065 = (n2877 | n3931) & (n2879 | n3932);
  assign n3066 = n3062 & n3065 & (n2860 | n1948);
  assign n3067 = (n2884 | n3931) & (n2886 | n3932);
  assign n3068 = n3062 & n3067 & (n2853 | n1948);
  assign n3069 = (n3068 | n3864) & (n3066 | n3867);
  assign n3070 = n4453 & n4451 & (n2479 | n3930);
  assign n3071 = n3069 & n3070 & (n3064 | n1322);
  assign n3072 = (n2897 | n3931) & (n2899 | n3932);
  assign n3073 = n3062 & n3072 & (n2858 | n1948);
  assign n3074 = (n2905 | n3931) & (n2907 | n3932);
  assign n3075 = n3062 & n3074 & (n2857 | n1948);
  assign n3076 = (n2912 | n3931) & (n2914 | n3932);
  assign n3077 = n3062 & n3076 & (n2851 | n1948);
  assign n3078 = (n3077 | n3864) & (n3075 | n3867);
  assign n3079 = n4450 & n4451 & (n2456 | n3930);
  assign n3080 = n3078 & n3079 & (n3073 | n1322);
  assign n3081 = (n2925 | n3931) & (n2927 | n3932);
  assign n3082 = n3062 & n3081 & (n2864 | n1948);
  assign n3083 = (n2933 | n3931) & (n2935 | n3932);
  assign n3084 = n3062 & n3083 & (n2863 | n1948);
  assign n3085 = (n2940 | n3931) & (n2942 | n3932);
  assign n3086 = n3062 & n3085 & (n2855 | n1948);
  assign n3087 = (n3086 | n3864) & (n3084 | n3867);
  assign n3088 = n4454 & n4451 & (n2513 | n3930);
  assign n3089 = n3087 & n3088 & (n3082 | n1322);
  assign n3090 = (n2953 | n3931) & (n2955 | n3932);
  assign n3091 = (Pi20 & n2591) | (n2586 & (~Pi20 | n2591));
  assign n3092 = n3062 & n3090 & (n3091 | n1948);
  assign n3093 = (n2961 | n3931) & (n2963 | n3932);
  assign n3094 = (Pi20 & n2581) | (n2576 & (~Pi20 | n2581));
  assign n3095 = n3062 & n3093 & (n3094 | n1948);
  assign n3096 = (n2968 | n3931) & (n2970 | n3932);
  assign n3097 = n3062 & n3096 & (n3046 | n1948);
  assign n3098 = (n3097 | n3864) & (n3095 | n3867);
  assign n3099 = n4452 & n4451 & (n2496 | n3930);
  assign n3100 = n3098 & n3099 & (n3092 | n1322);
  assign n3101 = n2628 & (n2629 | n1919);
  assign n3102 = (n2861 | n3922) & (n2869 | n3923);
  assign n3103 = n3101 & n3102 & (n2871 | n1989);
  assign n3104 = (n2860 | n3922) & (n2877 | n3923);
  assign n3105 = n3101 & n3104 & (n2879 | n1989);
  assign n3106 = (n2853 | n3922) & (n2884 | n3923);
  assign n3107 = n3101 & n3106 & (n2886 | n1989);
  assign n3108 = (n3107 | n3864) & (n3105 | n3867);
  assign n3109 = n4446 & n4444 & (n2892 | n3921);
  assign n3110 = n3108 & n3109 & (n3103 | n1322);
  assign n3111 = (n2858 | n3922) & (n2897 | n3923);
  assign n3112 = n3101 & n3111 & (n2899 | n1989);
  assign n3113 = (n2857 | n3922) & (n2905 | n3923);
  assign n3114 = n3101 & n3113 & (n2907 | n1989);
  assign n3115 = (n2851 | n3922) & (n2912 | n3923);
  assign n3116 = n3101 & n3115 & (n2914 | n1989);
  assign n3117 = (n3116 | n3864) & (n3114 | n3867);
  assign n3118 = n4443 & n4444 & (n2920 | n3921);
  assign n3119 = n3117 & n3118 & (n3112 | n1322);
  assign n3120 = (n2864 | n3922) & (n2925 | n3923);
  assign n3121 = n3101 & n3120 & (n2927 | n1989);
  assign n3122 = (n2863 | n3922) & (n2933 | n3923);
  assign n3123 = n3101 & n3122 & (n2935 | n1989);
  assign n3124 = (n2855 | n3922) & (n2940 | n3923);
  assign n3125 = n3101 & n3124 & (n2942 | n1989);
  assign n3126 = (n3125 | n3864) & (n3123 | n3867);
  assign n3127 = n4447 & n4444 & (n2948 | n3921);
  assign n3128 = n3126 & n3127 & (n3121 | n1322);
  assign n3129 = (n3091 | n3922) & (n2953 | n3923);
  assign n3130 = n3101 & n3129 & (n2955 | n1989);
  assign n3131 = (n3094 | n3922) & (n2961 | n3923);
  assign n3132 = n3101 & n3131 & (n2963 | n1989);
  assign n3133 = (n3046 | n3922) & (n2968 | n3923);
  assign n3134 = n3101 & n3133 & (n2970 | n1989);
  assign n3135 = (n3134 | n3864) & (n3132 | n3867);
  assign n3136 = n4445 & n4444 & (n2976 | n3921);
  assign n3137 = n3135 & n3136 & (n3130 | n1322);
  assign n3138 = n2624 & (n2625 | n1919);
  assign n3139 = (n2869 | n3926) & (n2871 | n3927);
  assign n3140 = n3138 & n3139 & (n2861 | n2028);
  assign n3141 = (n2877 | n3926) & (n2879 | n3927);
  assign n3142 = n3138 & n3141 & (n2860 | n2028);
  assign n3143 = (n2884 | n3926) & (n2886 | n3927);
  assign n3144 = n3138 & n3143 & (n2853 | n2028);
  assign n3145 = (n3144 | n3864) & (n3142 | n3867);
  assign n3146 = n4439 & n4437 & (n2479 | n3925);
  assign n3147 = n3145 & n3146 & (n3140 | n1322);
  assign n3148 = (n2897 | n3926) & (n2899 | n3927);
  assign n3149 = n3138 & n3148 & (n2858 | n2028);
  assign n3150 = (n2905 | n3926) & (n2907 | n3927);
  assign n3151 = n3138 & n3150 & (n2857 | n2028);
  assign n3152 = (n2912 | n3926) & (n2914 | n3927);
  assign n3153 = n3138 & n3152 & (n2851 | n2028);
  assign n3154 = (n3153 | n3864) & (n3151 | n3867);
  assign n3155 = n4436 & n4437 & (n2456 | n3925);
  assign n3156 = n3154 & n3155 & (n3149 | n1322);
  assign n3157 = (n2925 | n3926) & (n2927 | n3927);
  assign n3158 = n3138 & n3157 & (n2864 | n2028);
  assign n3159 = (n2933 | n3926) & (n2935 | n3927);
  assign n3160 = n3138 & n3159 & (n2863 | n2028);
  assign n3161 = (n2940 | n3926) & (n2942 | n3927);
  assign n3162 = n3138 & n3161 & (n2855 | n2028);
  assign n3163 = (n3162 | n3864) & (n3160 | n3867);
  assign n3164 = n4440 & n4437 & (n2513 | n3925);
  assign n3165 = n3163 & n3164 & (n3158 | n1322);
  assign n3166 = (n2953 | n3926) & (n2955 | n3927);
  assign n3167 = n3138 & n3166 & (n3091 | n2028);
  assign n3168 = (n2961 | n3926) & (n2963 | n3927);
  assign n3169 = n3138 & n3168 & (n3094 | n2028);
  assign n3170 = (n2968 | n3926) & (n2970 | n3927);
  assign n3171 = n3138 & n3170 & (n3046 | n2028);
  assign n3172 = (n3171 | n3864) & (n3169 | n3867);
  assign n3173 = n4438 & n4437 & (n2496 | n3925);
  assign n3174 = n3172 & n3173 & (n3167 | n1322);
  assign n3175 = ~n3677 & (~n4455 | ~n4456);
  assign n3176 = ~n3805 & ~n4723 & (Ni10 | ~n4002);
  assign n3177 = ~n3937 & (n2751 | n2752 | ~n4532);
  assign n3178 = ~n3766 & (n2793 | n2794 | ~n4587);
  assign n3179 = ~n1671 & (~n4588 | (~Ni11 & ~n2633));
  assign n3180 = (Ni11 | n2622) & (~n1543 | n2621);
  assign n3181 = ~n3180 & (n2072 | (n2073 & n2074));
  assign n3182 = (~n3707 & ~n4010) | (~Ni32 & (n3707 | ~n4010));
  assign n3183 = Ni36 | ~Ni38;
  assign n3184 = Pi19 & Pi17;
  assign n3185 = ~Ni45 | n3186;
  assign n3186 = Ni45 & Ni46;
  assign n3187 = ~Ni40 | (Ni30 & n1353);
  assign n3188 = (~n2073 | ~n4014) & (~n2072 | n4013);
  assign n3189 = ~Ni41 | (Ni30 & n1353);
  assign n3190 = (~n2073 | ~n4018) & (~n2072 | n4017);
  assign n3191 = ~n3186 & (Ni45 | ~n3661);
  assign n3192 = ~Ni47 | ~Ni48;
  assign n3193 = ~n3186 & (Ni45 | n3192);
  assign n3194 = Ni38 | ~Ni39;
  assign n3195 = Ni39 | Ni38;
  assign n3196 = (n3191 | n3194) & (n3193 | n3195);
  assign n3197 = ~Ni37 | n3196;
  assign n3198 = n3193 & (n3203 | ~Ni42);
  assign n3199 = n3197 & (~n814 | n3198);
  assign n3200 = n3333 & (Ni42 | n3191);
  assign n3201 = n3197 & (~n814 | n3200);
  assign n3202 = ~n797 & (n1539 | n3193);
  assign n3203 = n3193 & (n3191 | n3331);
  assign n3204 = n3198 & (Ni41 | n3203);
  assign n3205 = n3203 & (n3191 | n923);
  assign n3206 = n3198 & (Ni41 | n3205);
  assign n3207 = n3200 | n3854;
  assign n3208 = n3211 | (n817 & n3968);
  assign n3209 = n3208 & n3207 & n3197;
  assign n3210 = Ni37 | n3976;
  assign n3211 = n3204 & (n3206 | ~Ni40);
  assign n3212 = n3210 & (~n783 | n3211);
  assign n3213 = n3209 & (~n2530 | n3212);
  assign n3214 = ~n2426 & ~n3191 & (n2441 | ~n3193);
  assign n3215 = Ni41 | ~Ni42;
  assign n3216 = ~n3214 & (n3203 | n3215);
  assign n3217 = n3200 | n3855;
  assign n3218 = n3220 | (n853 & n3968);
  assign n3219 = n3218 & n3217 & n3197;
  assign n3220 = n3247 & (n3206 | ~Ni40);
  assign n3221 = n3210 & (~n783 | n3220);
  assign n3222 = n3219 & (~n2530 | n3221);
  assign n3223 = Pi20 | Pi19;
  assign n3224 = ~Pi20 | Pi19;
  assign n3225 = (n3213 | n3223) & (n3222 | n3224);
  assign n3226 = n3197 & n3210 & (n3206 | ~Ni38);
  assign n3227 = Pi21 & Pi19;
  assign n3228 = Pi22 & ~n3550;
  assign n3229 = n3227 & (n810 | (~n3226 & n3228));
  assign n3230 = n3232 | (n817 & n3968);
  assign n3231 = n3230 & n3207 & n3197;
  assign n3232 = n3276 & (n3205 | ~Ni40);
  assign n3233 = n3210 & (~n783 | n3232);
  assign n3234 = n3231 & (~n2530 | n3233);
  assign n3235 = (~Ni41 | n3205) & n3216;
  assign n3236 = n3238 | (n853 & n3968);
  assign n3237 = n3236 & n3217 & n3197;
  assign n3238 = n3235 & (n3205 | ~Ni40);
  assign n3239 = n3210 & (~n783 | n3238);
  assign n3240 = n3237 & (~n2530 | n3239);
  assign n3241 = (n3234 | n3223) & (n3240 | n3224);
  assign n3242 = n3197 & n3210 & (n3205 | ~Ni38);
  assign n3243 = n3227 & (n810 | (n3228 & ~n3242));
  assign n3244 = n3247 | (n853 & n3968);
  assign n3245 = n3244 & n3217 & n3197;
  assign n3246 = n698 | n3976;
  assign n3247 = n3198 & n3216;
  assign n3248 = n3246 & n3245 & (n1216 | n3247);
  assign n3249 = n3247 & (Ni40 | n3206);
  assign n3250 = n3210 & (~n783 | n3249);
  assign n3251 = n3249 | (n853 & n3968);
  assign n3252 = n3251 & n3217 & n3197;
  assign n3253 = (~n2434 | n3250) & n3252;
  assign n3254 = n3235 | (n853 & n3968);
  assign n3255 = n3254 & n3217 & n3197;
  assign n3256 = n3246 & n3255 & (n1216 | n3235);
  assign n3257 = n3235 & (Ni40 | n3205);
  assign n3258 = n3210 & (~n783 | n3257);
  assign n3259 = n3257 | (n853 & n3968);
  assign n3260 = n3259 & n3217 & n3197;
  assign n3261 = (~n2434 | n3258) & n3260;
  assign n3262 = ~n799 & ~n3977;
  assign n3263 = (n3256 | n3743) & (n3261 | n3737);
  assign n3264 = (n3248 | n2272) & (n3253 | n3895);
  assign n3265 = n3262 & (~n3288 | (n3263 & n3264));
  assign n3266 = n3204 | (n817 & n3968);
  assign n3267 = n3266 & n3207 & n3197;
  assign n3268 = n3246 & n3267 & (n1216 | n3204);
  assign n3269 = n3204 & (Ni40 | n3206);
  assign n3270 = n3210 & (~n783 | n3269);
  assign n3271 = n3269 | (n817 & n3968);
  assign n3272 = n3271 & n3207 & n3197;
  assign n3273 = (~n2434 | n3270) & n3272;
  assign n3274 = n3276 | (n817 & n3968);
  assign n3275 = n3274 & n3207 & n3197;
  assign n3276 = n3203 & (~Ni41 | n3205);
  assign n3277 = n3246 & n3275 & (n1216 | n3276);
  assign n3278 = n3276 & (Ni40 | n3205);
  assign n3279 = n3210 & (~n783 | n3278);
  assign n3280 = n3278 | (n817 & n3968);
  assign n3281 = n3280 & n3207 & n3197;
  assign n3282 = (~n2434 | n3279) & n3281;
  assign n3283 = ~n4732 & (Pi22 | ~Pi21 | n3202);
  assign n3284 = ~n799 & n3283;
  assign n3285 = (n3277 | n3743) & (n3282 | n3737);
  assign n3286 = (n3268 | n2272) & (n3273 | n3895);
  assign n3287 = n3284 & (~n3288 | (n3285 & n3286));
  assign n3288 = ~n2254 & ~n3550;
  assign n3289 = ~n3978 & (n3229 | (~n3225 & n3288));
  assign n3290 = ~n3979 & (n3243 | (~n3241 & n3288));
  assign n3291 = (n3211 | n698) & (n3212 | n2434);
  assign n3292 = n3291 & n3209;
  assign n3293 = (n3220 | n698) & (n3221 | n2434);
  assign n3294 = n3293 & n3219;
  assign n3295 = (n3292 | n3223) & (n3294 | n3224);
  assign n3296 = n3197 & (n3206 | n690);
  assign n3297 = n3296 & (Ni36 | n3226);
  assign n3298 = ~n3297 & n3227 & n3228;
  assign n3299 = (n3232 | n698) & (n3233 | n2434);
  assign n3300 = n3299 & n3231;
  assign n3301 = (n3238 | n698) & (n3239 | n2434);
  assign n3302 = n3301 & n3237;
  assign n3303 = (n3300 | n3223) & (n3302 | n3224);
  assign n3304 = n3197 & (n3205 | n690);
  assign n3305 = n3304 & (Ni36 | n3242);
  assign n3306 = n3227 & (n810 | (n3228 & ~n3305));
  assign n3307 = n3245 & (n3247 | n698);
  assign n3308 = (n3249 | n698) & (n3250 | n2530);
  assign n3309 = n3308 & n3252;
  assign n3310 = n3255 & (n3235 | n698);
  assign n3311 = (n3257 | n698) & (n3258 | n2530);
  assign n3312 = n3311 & n3260;
  assign n3313 = (n3310 | n3743) & (n3312 | n3737);
  assign n3314 = (n3307 | n2272) & (n3309 | n3895);
  assign n3315 = n3262 & (~n3288 | (n3313 & n3314));
  assign n3316 = n3267 & (n3204 | n698);
  assign n3317 = (n3269 | n698) & (n3270 | n2530);
  assign n3318 = n3317 & n3272;
  assign n3319 = n3275 & (n3276 | n698);
  assign n3320 = (n3278 | n698) & (n3279 | n2530);
  assign n3321 = n3320 & n3281;
  assign n3322 = (n3319 | n3743) & (n3321 | n3737);
  assign n3323 = (n3316 | n2272) & (n3318 | n3895);
  assign n3324 = n3284 & (~n3288 | (n3322 & n3323));
  assign n3325 = ~n3978 & ((n3288 & ~n3295) | n3298);
  assign n3326 = ~n3979 & ((n3288 & ~n3303) | n3306);
  assign n3327 = Ni11 | n1446;
  assign n3328 = n3327 & (~n807 | (~n2254 & ~n3471));
  assign n3329 = ~n3944 & (n3325 | n3326 | ~n4030);
  assign n3330 = ~n2367 & (n3289 | n3290 | ~n4031);
  assign n3331 = ~Ni44 | Ni43;
  assign n3332 = ~n2426 & ~n3191 & (~n3193 | n3331);
  assign n3333 = n3193 & (n2441 | n3191);
  assign n3334 = ~n3332 & (n3215 | n3333);
  assign n3335 = n3193 & (n3191 | n3754);
  assign n3336 = n3335 & (n3333 | ~Ni42);
  assign n3337 = n3353 & (Ni40 | n3395);
  assign n3338 = n3337 | n817;
  assign n3339 = Ni37 | n3974;
  assign n3340 = n3337 | (~n783 & n3968);
  assign n3341 = n3340 & n3339 & n3197;
  assign n3342 = n3337 | n698;
  assign n3343 = n3341 & n3342 & (Ni35 | n3338);
  assign n3344 = ~n797 & n3480;
  assign n3345 = (~Ni33 | n3343) & n3344;
  assign n3346 = n3353 & (Ni40 | n3401);
  assign n3347 = n3346 | n853;
  assign n3348 = n3346 | (~n783 & n3968);
  assign n3349 = n3348 & n3339 & n3197;
  assign n3350 = n3346 | n698;
  assign n3351 = n3349 & n3350 & (Ni35 | n3347);
  assign n3352 = n3344 & (~Ni33 | n3351);
  assign n3353 = n3336 & n3836;
  assign n3354 = n3197 & n3339 & (n3353 | ~Ni38);
  assign n3355 = n3354 & (n3353 | n690);
  assign n3356 = n3344 & (~Ni33 | n3355);
  assign n3357 = (n3345 | n1408) & (n3352 | n914);
  assign n3358 = n807 & n3357 & (n3356 | n1702);
  assign n3359 = n3336 & (Ni40 | n3423);
  assign n3360 = n3359 | n817;
  assign n3361 = n3359 | (~n783 & n3968);
  assign n3362 = n3361 & n3339 & n3197;
  assign n3363 = n3359 | n698;
  assign n3364 = n3362 & n3363 & (Ni35 | n3360);
  assign n3365 = n3344 & (~Ni33 | n3364);
  assign n3366 = n3336 & (Ni40 | n3428);
  assign n3367 = n3366 | n853;
  assign n3368 = n3366 | (~n783 & n3968);
  assign n3369 = n3368 & n3339 & n3197;
  assign n3370 = n3366 | n698;
  assign n3371 = n3369 & n3370 & (Ni35 | n3367);
  assign n3372 = n3344 & (~Ni33 | n3371);
  assign n3373 = n3197 & n3339 & (n3336 | ~Ni38);
  assign n3374 = n3373 & (n3336 | n690);
  assign n3375 = n3344 & (~Ni33 | n3374);
  assign n3376 = (n3365 | n1408) & (n3372 | n914);
  assign n3377 = n807 & n3376 & (n3375 | n1702);
  assign n3378 = n3341 & (Ni35 | n3338);
  assign n3379 = n3344 & (~Ni33 | n3378);
  assign n3380 = n3349 & (Ni35 | n3347);
  assign n3381 = n3344 & (~Ni33 | n3380);
  assign n3382 = n3344 & (~Ni33 | n3354);
  assign n3383 = (n3379 | n1408) & (n3381 | n914);
  assign n3384 = n807 & n3383 & (n3382 | n1702);
  assign n3385 = n3362 & (Ni35 | n3360);
  assign n3386 = n3344 & (~Ni33 | n3385);
  assign n3387 = n3369 & (Ni35 | n3367);
  assign n3388 = n3344 & (~Ni33 | n3387);
  assign n3389 = n3344 & (~Ni33 | n3373);
  assign n3390 = (n3386 | n1408) & (n3388 | n914);
  assign n3391 = n807 & n3390 & (n3389 | n1702);
  assign n3392 = n3198 | n3854;
  assign n3393 = n3395 | (n817 & n3968);
  assign n3394 = n3393 & n3392 & n3197;
  assign n3395 = n3836 & n3334;
  assign n3396 = n3394 & (n3395 | n698);
  assign n3397 = n3344 & (~Ni33 | n3396);
  assign n3398 = n3198 | n3855;
  assign n3399 = n3401 | (n853 & n3968);
  assign n3400 = n3399 & n3398 & n3197;
  assign n3401 = n3333 & n3836;
  assign n3402 = n3400 & (n3401 | n698);
  assign n3403 = n3344 & (~Ni33 | n3402);
  assign n3404 = n3406 | (~n783 & n3968);
  assign n3405 = n3404 & n3339 & n3197;
  assign n3406 = n3353 & (n3395 | ~Ni40);
  assign n3407 = n3406 | n817;
  assign n3408 = n3406 | n698;
  assign n3409 = n3405 & n3408 & (~Ni35 | n3407);
  assign n3410 = n3344 & (~Ni33 | n3409);
  assign n3411 = n3413 | (~n783 & n3968);
  assign n3412 = n3411 & n3339 & n3197;
  assign n3413 = n3353 & (n3401 | ~Ni40);
  assign n3414 = n3413 | n853;
  assign n3415 = n3413 | n698;
  assign n3416 = n3412 & n3415 & (~Ni35 | n3414);
  assign n3417 = n3344 & (~Ni33 | n3416);
  assign n3418 = n807 & (n3410 | n3893);
  assign n3419 = (n3397 | n1408) & (n3403 | n914);
  assign n3420 = n3418 & n3419 & (n3417 | n2109);
  assign n3421 = n3423 | (n817 & n3968);
  assign n3422 = n3421 & n3392 & n3197;
  assign n3423 = n3336 & n3334;
  assign n3424 = n3422 & (n3423 | n698);
  assign n3425 = n3344 & (~Ni33 | n3424);
  assign n3426 = n3428 | (n853 & n3968);
  assign n3427 = n3426 & n3398 & n3197;
  assign n3428 = n3336 & (Ni41 | n3333);
  assign n3429 = n3427 & (n3428 | n698);
  assign n3430 = n3344 & (~Ni33 | n3429);
  assign n3431 = n3433 | (~n783 & n3968);
  assign n3432 = n3431 & n3339 & n3197;
  assign n3433 = n3336 & (n3423 | ~Ni40);
  assign n3434 = n3433 | n817;
  assign n3435 = n3433 | n698;
  assign n3436 = n3432 & n3435 & (~Ni35 | n3434);
  assign n3437 = n3344 & (~Ni33 | n3436);
  assign n3438 = n3440 | (~n783 & n3968);
  assign n3439 = n3438 & n3339 & n3197;
  assign n3440 = n3336 & (n3428 | ~Ni40);
  assign n3441 = n3440 | n853;
  assign n3442 = n3440 | n698;
  assign n3443 = n3439 & n3442 & (~Ni35 | n3441);
  assign n3444 = n3344 & (~Ni33 | n3443);
  assign n3445 = n807 & (n3437 | n3893);
  assign n3446 = (n3425 | n1408) & (n3430 | n914);
  assign n3447 = n3445 & n3446 & (n3444 | n2109);
  assign n3448 = n698 | n3974;
  assign n3449 = n3448 & n3394 & (n1216 | n3395);
  assign n3450 = n3344 & (~Ni33 | n3449);
  assign n3451 = n3448 & n3400 & (n1216 | n3401);
  assign n3452 = n3344 & (~Ni33 | n3451);
  assign n3453 = n3405 & (~Ni35 | n3407);
  assign n3454 = n3344 & (~Ni33 | n3453);
  assign n3455 = n3412 & (~Ni35 | n3414);
  assign n3456 = n3344 & (~Ni33 | n3455);
  assign n3457 = n807 & (n3454 | n3893);
  assign n3458 = (n3450 | n1408) & (n3452 | n914);
  assign n3459 = n3457 & n3458 & (n3456 | n2109);
  assign n3460 = n3448 & n3422 & (n1216 | n3423);
  assign n3461 = n3344 & (~Ni33 | n3460);
  assign n3462 = n3448 & n3427 & (n1216 | n3428);
  assign n3463 = n3344 & (~Ni33 | n3462);
  assign n3464 = n3432 & (~Ni35 | n3434);
  assign n3465 = n3344 & (~Ni33 | n3464);
  assign n3466 = n3439 & (~Ni35 | n3441);
  assign n3467 = n3344 & (~Ni33 | n3466);
  assign n3468 = n807 & (n3465 | n3893);
  assign n3469 = (n3461 | n1408) & (n3463 | n914);
  assign n3470 = n3468 & n3469 & (n3467 | n2109);
  assign n3471 = ~n809 & n3480;
  assign n3472 = n807 & (n3471 | n1919);
  assign n3473 = (~n2345 | n3389) & (n3382 | ~n3772);
  assign n3474 = ~n2272 & (~n3472 | ~n4604);
  assign n3475 = ~n3743 & (~n3472 | ~n4606);
  assign n3476 = (~n2345 | n3375) & (n3356 | ~n3772);
  assign n3477 = ~n3740 & (~n3472 | ~n4593);
  assign n3478 = ~n2272 & (~n3472 | ~n4594);
  assign n3479 = ~n3743 & (~n3472 | ~n4596);
  assign n3480 = n1539 | Ni33 | n3199;
  assign n3481 = ~Ni34 | n3201;
  assign n3482 = ~n797 & n3480 & (~Ni33 | n3481);
  assign n3483 = Ni34 | ~Ni33;
  assign n3484 = n3482 & (n3343 | n3483);
  assign n3485 = n3482 & (n3351 | n3483);
  assign n3486 = n3482 & (n3355 | n3483);
  assign n3487 = (n3484 | n1408) & (n3485 | n914);
  assign n3488 = n807 & n3487 & (n3486 | n1702);
  assign n3489 = n3482 & (n3364 | n3483);
  assign n3490 = n3482 & (n3371 | n3483);
  assign n3491 = n3482 & (n3374 | n3483);
  assign n3492 = (n3489 | n1408) & (n3490 | n914);
  assign n3493 = n807 & n3492 & (n3491 | n1702);
  assign n3494 = n3482 & (n3378 | n3483);
  assign n3495 = n3482 & (n3380 | n3483);
  assign n3496 = n3482 & (n3354 | n3483);
  assign n3497 = (n3494 | n1408) & (n3495 | n914);
  assign n3498 = n807 & n3497 & (n3496 | n1702);
  assign n3499 = n3482 & (n3385 | n3483);
  assign n3500 = n3482 & (n3387 | n3483);
  assign n3501 = n3482 & (n3373 | n3483);
  assign n3502 = (n3499 | n1408) & (n3500 | n914);
  assign n3503 = n807 & n3502 & (n3501 | n1702);
  assign n3504 = n3482 & (n3396 | n3483);
  assign n3505 = n3482 & (n3402 | n3483);
  assign n3506 = n3482 & (n3409 | n3483);
  assign n3507 = n3482 & (n3416 | n3483);
  assign n3508 = n807 & (n3506 | n3893);
  assign n3509 = (n3504 | n1408) & (n3505 | n914);
  assign n3510 = n3508 & n3509 & (n3507 | n2109);
  assign n3511 = n3482 & (n3424 | n3483);
  assign n3512 = n3482 & (n3429 | n3483);
  assign n3513 = n3482 & (n3436 | n3483);
  assign n3514 = n3482 & (n3443 | n3483);
  assign n3515 = n807 & (n3513 | n3893);
  assign n3516 = (n3511 | n1408) & (n3512 | n914);
  assign n3517 = n3515 & n3516 & (n3514 | n2109);
  assign n3518 = n3482 & (n3449 | n3483);
  assign n3519 = n3482 & (n3451 | n3483);
  assign n3520 = n3482 & (n3453 | n3483);
  assign n3521 = n3482 & (n3455 | n3483);
  assign n3522 = n807 & (n3520 | n3893);
  assign n3523 = (n3518 | n1408) & (n3519 | n914);
  assign n3524 = n3522 & n3523 & (n3521 | n2109);
  assign n3525 = n3482 & (n3460 | n3483);
  assign n3526 = n3482 & (n3462 | n3483);
  assign n3527 = n3482 & (n3464 | n3483);
  assign n3528 = n3482 & (n3466 | n3483);
  assign n3529 = n807 & (n3527 | n3893);
  assign n3530 = (n3525 | n1408) & (n3526 | n914);
  assign n3531 = n3529 & n3530 & (n3528 | n2109);
  assign n3532 = (~n2345 | n3501) & (n3496 | ~n3772);
  assign n3533 = ~n2272 & (~n3472 | ~n4625);
  assign n3534 = ~n3743 & (~n3472 | ~n4627);
  assign n3535 = (~n2345 | n3491) & (n3486 | ~n3772);
  assign n3536 = ~n3740 & (~n3472 | ~n4614);
  assign n3537 = ~n2272 & (~n3472 | ~n4615);
  assign n3538 = ~n3743 & (~n3472 | ~n4617);
  assign n3539 = n3975 | Ni34 | n3199;
  assign n3540 = ~n797 & n3539 & (~Ni33 | n3481);
  assign n3541 = n3292 | n3550;
  assign n3542 = n3541 & n3540 & (n3343 | n3483);
  assign n3543 = n3294 | n3550;
  assign n3544 = n3543 & n3540 & (n3351 | n3483);
  assign n3545 = (n3297 | n3550) & (n3355 | n3483);
  assign n3546 = n3545 & n3540;
  assign n3547 = (n3542 | n1408) & (n3544 | n914);
  assign n3548 = n807 & n3547 & (n3546 | n1702);
  assign n3549 = n3364 | n3483;
  assign n3550 = n1539 | n3953;
  assign n3551 = n3549 & n3540 & (n3300 | n3550);
  assign n3552 = n3371 | n3483;
  assign n3553 = n3552 & n3540 & (n3302 | n3550);
  assign n3554 = (n3305 | n3550) & (n3374 | n3483);
  assign n3555 = n3554 & n3540;
  assign n3556 = (n3551 | n1408) & (n3553 | n914);
  assign n3557 = n807 & n3556 & (n3555 | n1702);
  assign n3558 = n3213 | n3550;
  assign n3559 = n3558 & n3540 & (n3378 | n3483);
  assign n3560 = n3222 | n3550;
  assign n3561 = n3560 & n3540 & (n3380 | n3483);
  assign n3562 = (n3226 | n3550) & (n3354 | n3483);
  assign n3563 = n3562 & n3540;
  assign n3564 = (n3559 | n1408) & (n3561 | n914);
  assign n3565 = n807 & n3564 & (n3563 | n1702);
  assign n3566 = n3385 | n3483;
  assign n3567 = n3566 & n3540 & (n3234 | n3550);
  assign n3568 = n3387 | n3483;
  assign n3569 = n3568 & n3540 & (n3240 | n3550);
  assign n3570 = (n3242 | n3550) & (n3373 | n3483);
  assign n3571 = n3570 & n3540;
  assign n3572 = (n3567 | n1408) & (n3569 | n914);
  assign n3573 = n807 & n3572 & (n3571 | n1702);
  assign n3574 = n3316 | n3550;
  assign n3575 = n3574 & n3540 & (n3396 | n3483);
  assign n3576 = n3307 | n3550;
  assign n3577 = n3576 & n3540 & (n3402 | n3483);
  assign n3578 = n3318 | n3550;
  assign n3579 = n3578 & n3540 & (n3409 | n3483);
  assign n3580 = n3309 | n3550;
  assign n3581 = n3580 & n3540 & (n3416 | n3483);
  assign n3582 = n807 & (n3579 | n3893);
  assign n3583 = (n3575 | n1408) & (n3577 | n914);
  assign n3584 = n3582 & n3583 & (n3581 | n2109);
  assign n3585 = n3424 | n3483;
  assign n3586 = n3585 & n3540 & (n3319 | n3550);
  assign n3587 = n3429 | n3483;
  assign n3588 = n3587 & n3540 & (n3310 | n3550);
  assign n3589 = n3436 | n3483;
  assign n3590 = n3589 & n3540 & (n3321 | n3550);
  assign n3591 = n3443 | n3483;
  assign n3592 = n3591 & n3540 & (n3312 | n3550);
  assign n3593 = n807 & (n3590 | n3893);
  assign n3594 = (n3586 | n1408) & (n3588 | n914);
  assign n3595 = n3593 & n3594 & (n3592 | n2109);
  assign n3596 = n3268 | n3550;
  assign n3597 = n3596 & n3540 & (n3449 | n3483);
  assign n3598 = n3248 | n3550;
  assign n3599 = n3598 & n3540 & (n3451 | n3483);
  assign n3600 = n3273 | n3550;
  assign n3601 = n3600 & n3540 & (n3453 | n3483);
  assign n3602 = n3253 | n3550;
  assign n3603 = n3602 & n3540 & (n3455 | n3483);
  assign n3604 = n807 & (n3601 | n3893);
  assign n3605 = (n3597 | n1408) & (n3599 | n914);
  assign n3606 = n3604 & n3605 & (n3603 | n2109);
  assign n3607 = n3460 | n3483;
  assign n3608 = n3607 & n3540 & (n3277 | n3550);
  assign n3609 = n3462 | n3483;
  assign n3610 = n3609 & n3540 & (n3256 | n3550);
  assign n3611 = n3464 | n3483;
  assign n3612 = n3611 & n3540 & (n3282 | n3550);
  assign n3613 = n3466 | n3483;
  assign n3614 = n3613 & n3540 & (n3261 | n3550);
  assign n3615 = n807 & (n3612 | n3893);
  assign n3616 = (n3608 | n1408) & (n3610 | n914);
  assign n3617 = n3615 & n3616 & (n3614 | n2109);
  assign n3618 = n2254 | n3624;
  assign n3619 = n3561 & ~n3635 & (n3222 | n3618);
  assign n3620 = n3213 | n3618;
  assign n3621 = ~n798 & n3283;
  assign n3622 = n3620 & n3621 & (n3559 | n1929);
  assign n3623 = Pi25 | ~n809;
  assign n3624 = Pi25 | n3975;
  assign n3625 = n3623 & n3563 & (n3226 | n3624);
  assign n3626 = (n3622 | n3223) & (n3619 | n3224);
  assign n3627 = ~Pi22 | ~n3227;
  assign n3628 = n807 & n3626 & (n3625 | n3627);
  assign n3629 = n3623 & n3571 & (n3242 | n3624);
  assign n3630 = ~n3223 & (~n3621 | ~n4646);
  assign n3631 = ~n3630 & (n3224 | (~n3635 & n4647));
  assign n3632 = n807 & n3631 & (n3629 | n3627);
  assign n3633 = n3599 & ~n3635 & (n3248 | n3618);
  assign n3634 = n3603 & ~n3635 & (n3253 | n3618);
  assign n3635 = n798 | n3977;
  assign n3636 = ~n3743 & (n3635 | ~n4654);
  assign n3637 = ~n3737 & (n3635 | ~n4655);
  assign n3638 = ~n2272 & (~n3621 | ~n4648);
  assign n3639 = ~n3743 & (~n3621 | ~n4650);
  assign n3640 = n3544 & ~n3635 & (n3294 | n3618);
  assign n3641 = n3292 | n3618;
  assign n3642 = n3641 & n3621 & (n3542 | n1929);
  assign n3643 = n3623 & n3546 & (n3297 | n3624);
  assign n3644 = (n3642 | n3223) & (n3640 | n3224);
  assign n3645 = n807 & n3644 & (n3643 | n3627);
  assign n3646 = n3623 & n3555 & (n3305 | n3624);
  assign n3647 = ~n3223 & (~n3621 | ~n4634);
  assign n3648 = ~n3647 & (n3224 | (~n3635 & n4635));
  assign n3649 = n807 & n3648 & (n3646 | n3627);
  assign n3650 = n3577 & ~n3635 & (n3307 | n3618);
  assign n3651 = n3581 & ~n3635 & (n3309 | n3618);
  assign n3652 = ~n3743 & (n3635 | ~n4642);
  assign n3653 = ~n3737 & (n3635 | ~n4643);
  assign n3654 = ~n2272 & (~n3621 | ~n4636);
  assign n3655 = ~n3743 & (~n3621 | ~n4638);
  assign n3656 = ~n4739 & (~Pi17 | ~n4660 | ~n4661);
  assign n3657 = ~n3327 & ~n4740 & (~Ni10 | n3656);
  assign n3658 = (~n3707 & ~n4032) | (~Ni33 & (n3707 | ~n4032));
  assign n3659 = n3707 | n3805;
  assign n3660 = n4662 & (~n4029 | (~n1543 & ~Ni13));
  assign n3661 = ~Ni47 | ~n3192;
  assign n3662 = ~n900 & n3661 & (Pi20 | ~n3192);
  assign n3663 = Ni30 | n801;
  assign n3664 = Ni47 & (n801 | Ni30);
  assign n3665 = n1353 & Ni30;
  assign n3666 = n1463 & Ni30;
  assign n3667 = Ni12 | ~n3727;
  assign n3668 = n3665 & (n3666 | n3667);
  assign n3669 = n1354 & Ni30;
  assign n3670 = n1553 & n1542 & n1543;
  assign n3671 = n4750 & (Ni12 | n3679);
  assign n3672 = ~Pi26 & n3981;
  assign n3673 = n3670 & n3671 & (Ni14 | n3672);
  assign n3674 = (n3841 | n3696) & (n3838 | n2632);
  assign n3675 = ~n3842 & (n3670 | (Pi24 & n3666));
  assign n3676 = n3695 & (Pi26 | n3666);
  assign n3677 = n1446 | ~Ni11;
  assign n3678 = n3674 & n3675 & (n3676 | n3677);
  assign n3679 = Pi26 & n3981;
  assign n3680 = (n3672 | n2632) & (n3679 | n3677);
  assign n3681 = ~n3696 & ~n4775 & (n788 | ~n3841);
  assign n3682 = n3840 & (~Pi23 | (n3670 & n3680));
  assign n3683 = ~Pi24 & n3666;
  assign n3684 = ~n3681 & n3682 & (n3670 | n3683);
  assign n3685 = ~n3696 & ~n4775 & (n795 | ~n3841);
  assign n3686 = n3840 & (Pi23 | (n3670 & n3680));
  assign n3687 = ~n3685 & (n3670 | n3683) & n3686;
  assign n3688 = Ni7 | Ni8;
  assign n3689 = n3688 & n1670 & (Ni8 | Ni10);
  assign n3690 = (n3687 | n3766) & (n3673 | n3689);
  assign n3691 = (n3684 | n3937) & (n3678 | n2066);
  assign n3692 = n3690 & n3691;
  assign n3693 = ~n3692 & (~Ni6 | ~Ni5);
  assign n3694 = n2632 | Pi26 | n3841;
  assign n3695 = n3665 & (~Pi27 | n3666);
  assign n3696 = ~Ni12 | n2750;
  assign n3697 = n3694 & n3668 & (n3695 | n3696);
  assign n3698 = n3665 & (~Pi26 | n3677 | n3841);
  assign n3699 = n4663 & n4664 & (n3669 | n3982);
  assign n3700 = n3698 & n3699 & (Ni11 | n3697);
  assign n3701 = (Ni32 | n2399) & (n801 | ~Ni41);
  assign n3702 = ~Ni5 & (~Ni31 | ~Ni6 | ~n3980);
  assign n3703 = ~n3707 & (n780 | (~Ni6 & ~n3692));
  assign n3704 = Ni4 | n3711;
  assign n3705 = ~n3703 & ~Ni2 & (Ni31 | n3704);
  assign n3706 = n3701 & Ni30;
  assign n3707 = Ni2 | Ni3;
  assign n3708 = (n1353 | n3704) & (~n3700 | n3707);
  assign n3709 = n3702 | n3711 | ~Ni4 | ~n4752;
  assign n3710 = (~Ni5 | n3705) & (n3706 | n3983);
  assign n3711 = Ni2 | ~Ni3;
  assign n3712 = (~n3700 | n3707) & (n3711 | ~n4665);
  assign n3713 = (~n780 | n3707) & (n3980 | n3983);
  assign n3714 = ~Ni9 & ~Ni7;
  assign n3715 = ~n3707 & (~n3957 | (n3714 & ~n3767));
  assign n3716 = (~n795 | ~Ni7) & (n3688 | n3950);
  assign n3717 = n3716 & (Pi24 | ~Ni8);
  assign n3718 = ~Ni10 | n3707 | n3717 | ~n3957;
  assign n3719 = (~n788 | Ni10) & ~Ni9;
  assign n3720 = (n773 | n3688) & (~Ni8 | n3719);
  assign n3721 = (Ni10 | ~Ni7) & (n3720 | ~n3957);
  assign n3722 = (~n789 & ~Ni14) | (Pi27 & (~n789 | Ni14));
  assign n3723 = n3722 & ~Ni11 & ~Ni13;
  assign n3724 = (n785 | n1543) & (~Ni11 | ~n3761);
  assign n3725 = n3724 & (Pi27 | ~Ni12);
  assign n3726 = ~Ni14 | n3707 | n3725 | ~n3727;
  assign n3727 = ~Ni14 | ~Ni13;
  assign n3728 = n789 & ~Ni14 & Ni12;
  assign n3729 = ~n1543 & n785 & Ni14;
  assign n3730 = n3727 & (n3728 | n3729 | Ni13);
  assign n3731 = ~n3707 & ((Ni11 & ~Ni14) | n3730);
  assign n3732 = ~Ni42 | ~Ni43;
  assign n3733 = Ni44 | ~Ni43;
  assign n3734 = n3732 & (n2426 | n3733);
  assign n3735 = ~Ni41 | ~Ni43;
  assign n3736 = (n3740 | ~Ni43) & (n3844 | n3894);
  assign n3737 = ~Pi16 | n1322;
  assign n3738 = n3734 & n3736 & (n3735 | n3737);
  assign n3739 = (n3737 | ~Ni43) & (n3844 | n3895);
  assign n3740 = ~Pi16 | n3864;
  assign n3741 = n3734 & n3739 & (n3735 | n3740);
  assign n3742 = (n3738 & (n3741 | Ni40)) | (n3741 & ~Ni40);
  assign n3743 = ~Pi16 | n3867;
  assign n3744 = n3742 & (n3735 | n3743);
  assign n3745 = ~Ni44 | ~Ni43;
  assign n3746 = n3732 & (n2426 | n3745);
  assign n3747 = n3746 & n3736 & (n3735 | n3737);
  assign n3748 = n3746 & n3739 & (n3735 | n3740);
  assign n3749 = (n3747 & (n3748 | Ni40)) | (n3748 & ~Ni40);
  assign n3750 = n3749 & (n3735 | n3743);
  assign n3751 = Ni31 | n784;
  assign n3752 = (~n2345 | ~Ni43) & (~n3772 | n3844);
  assign n3753 = (~Pi20 & n3750) | (n3744 & (Pi20 | n3750));
  assign n3754 = Ni42 | ~Ni43;
  assign n3755 = n2426 | ~Ni40;
  assign n3756 = n3733 | n3755;
  assign n3757 = n3756 | (Ni30 & ~n3984);
  assign n3758 = (n801 | Ni41) & (~Ni31 | n887);
  assign n1090_1 = ~n3711;
  assign n3760 = Ni4 & ~n3711 & ~n2418 & ~n3701;
  assign n3761 = Pi27 | ~Pi26;
  assign n3762 = (~Ni12 | ~n3723) & (n3677 | n3761);
  assign n3763 = ~n3795 & (n3760 | (~n3758 & ~n3983));
  assign n3764 = Ni30 | n2418 | n3704 | ~n3973;
  assign n3765 = n887 & (~Ni32 | Ni41);
  assign n3766 = ~Ni10 | n2074 | ~Ni7;
  assign n3767 = (~Pi24 & (n788 | Ni10)) | (n788 & ~Ni10);
  assign n3768 = ~Ni8 | Ni9 | Ni7;
  assign n3769 = (n795 | n3766) & (n3767 | n3768);
  assign n3770 = n2418 | n3711 | n4764 | n4765;
  assign n3771 = n1353 | n3983 | Ni33 | n3765;
  assign n3772 = ~Pi16 & n3184;
  assign n3773 = ~n3472 & (n2345 | n3772);
  assign n986 = n2407 | n2408 | n2415 | ~n4379;
  assign n3775 = ~n2417 & (Pi21 | n801) & n3810;
  assign n946_1 = ~n3775;
  assign n3777 = n900 & n3837 & (~Ni47 | ~n3711);
  assign n936 = ~n3777;
  assign n3779 = n3845 & ((n655 & Ni30) | ~n4050);
  assign n3780 = ~n3754 & Ni41 & ~Pi16 & ~n806;
  assign n3781 = n3846 & ~n4758 & (Pi20 | ~n3757);
  assign n961_1 = n3781 | n3779 | n3780;
  assign n3783 = Pi20 & (~n905 | (~Pi21 & ~n1116));
  assign n3784 = ~Pi20 & (~n905 | (~Pi21 & ~n1091));
  assign n3785 = Pi20 & (~n905 | (~Pi21 & ~n1249));
  assign n3786 = ~Pi20 & (~n905 | (~Pi21 & ~n1239));
  assign n3787 = Pi20 & (~n905 | (~Pi21 & ~n1196));
  assign n3788 = ~Pi20 & (~n905 | (~Pi21 & ~n1172));
  assign n3789 = ~n901 | n1209 | n3787 | n3788;
  assign n3790 = Pi20 & (~n905 | (~Pi21 & ~n1281));
  assign n3791 = ~Pi20 & (~n905 | (~Pi21 & ~n1274));
  assign n3792 = ~n901 | n1288 | n3790 | n3791;
  assign n3793 = n1540 & n1354;
  assign n3794 = (~Pi27 | n1918) & n3793;
  assign n3795 = ~Ni30 | ~Ni33;
  assign n3796 = n1354 & (~n789 | ~Ni30);
  assign n3797 = n1353 & (~n789 | n1463);
  assign n3798 = ~Pi21 & ~n3796;
  assign n3799 = ~Pi22 & ~n3796;
  assign n3800 = ~Pi24 & (n3798 | n3799 | ~n4300);
  assign n3801 = n1354 & (Pi27 | ~Ni30);
  assign n3802 = n1353 & (Pi27 | n1463);
  assign n3803 = Ni14 & ~n3801 & (Pi24 | ~n3802);
  assign n3804 = ~n3803 & (n1540 | n2254);
  assign n3805 = Ni7 | n2074;
  assign n3806 = Ni34 & n3805 & (n3327 | ~n3995);
  assign n3807 = ~n665 | Ni33;
  assign n3808 = n2390 & (~Pi26 | ~n665) & n3807;
  assign n3809 = n2400 & (~Pi27 | ~n665) & n3807;
  assign n3810 = n903 & (~Ni45 | (~n2418 & ~n3704));
  assign n3811 = n2425 & (Ni42 | Ni47);
  assign n3812 = n784 & n811;
  assign n3813 = n802 & n2424;
  assign n3814 = (n3824 | n2254) & (Pi27 | n3822);
  assign n3815 = n801 & n811;
  assign n3816 = n2649 & n3814 & (n3815 | n2643);
  assign n3817 = (~Pi27 | n3037) & n3813;
  assign n3818 = n2623 & (~Pi26 | ~Ni32);
  assign n3819 = n802 & n811;
  assign n3820 = (~Pi27 | n3812) & n3819;
  assign n3821 = (~Pi26 | n3812) & n3820;
  assign n3822 = n2419 & n812;
  assign n3823 = (~Pi27 | n813) & n3815;
  assign n3824 = n801 & n2424;
  assign n3825 = n2424 & n812;
  assign n3826 = n3820 & (Pi26 | n3812);
  assign n3827 = n3969 & n3187;
  assign n3828 = n800 & n3827 & (~Pi26 | n3751);
  assign n3829 = n2406 & n3956;
  assign n3830 = ~n3828 & (Pi23 | ~n3827 | n3829);
  assign n3831 = n3972 & n3189;
  assign n3832 = n800 & n3831 & (~Pi27 | n3751);
  assign n3833 = ~n3832 & (Pi24 | n3829 | ~n3831);
  assign n3834 = ~Pi22 & (n797 | (~n1539 & ~n3191));
  assign n3835 = ~Pi21 & (n797 | (~n1539 & n3185));
  assign n3836 = n3200 | ~Ni41;
  assign n3837 = ~n3664 & (~Ni47 | (~n2418 & ~Ni4));
  assign n3838 = (~Pi26 | n3666) & n3695;
  assign n3839 = (n3838 | n2632) & (n3676 | n3677);
  assign n3840 = (~Pi24 | n3680) & n3839;
  assign n3841 = n3665 & (Pi27 | n3666);
  assign n3842 = ~Pi24 & (~n3680 | (~n3696 & ~n4775));
  assign n3843 = n3669 & (Ni11 | n3667);
  assign n3844 = Ni41 | ~Ni43;
  assign n3845 = ~n806 & (Ni30 | ~n986_1 | n3732);
  assign n3846 = Pi18 & ~Pi17;
  assign n3847 = n18 | n2254;
  assign n3848 = n2254 | ~n3184;
  assign n3849 = n677 & ~Ni47;
  assign n3850 = ~n18 | n2416;
  assign n3851 = Ni36 | n1241;
  assign n3852 = Ni37 | Ni36;
  assign n3853 = Ni38 | n3852;
  assign n3854 = n3853 | ~Ni39;
  assign n3855 = Ni39 | n3853;
  assign n3856 = Ni32 | n2434;
  assign n3857 = Pi20 | n2254;
  assign n3858 = Pi25 | n3857;
  assign n3859 = ~Pi20 | n2254;
  assign n3860 = Pi25 | n3859;
  assign n3861 = Pi20 & (~n905 | (~Pi21 & ~n868));
  assign n3862 = ~Pi20 & (~n905 | (~Pi21 & ~n835));
  assign n3863 = ~n901 | n909 | n3861 | n3862;
  assign n3864 = Pi19 | ~Pi17;
  assign n3865 = Pi20 & (~n905 | (~Pi21 & ~n1068));
  assign n3866 = ~Pi20 & (~n905 | (~Pi21 & ~n1053));
  assign n3867 = Pi17 | Pi19;
  assign n3868 = ~Ni32 | n2530;
  assign n3869 = Ni32 | n2530;
  assign n3870 = Pi16 | Pi15;
  assign n3871 = Pi20 & (~n905 | (~Pi21 & ~n1004));
  assign n3872 = ~Pi20 & (~n905 | (~Pi21 & ~n993));
  assign n3873 = ~n901 | n1015 | n3871 | n3872;
  assign n3874 = n677 & ~Ni45;
  assign n3875 = Pi20 & (~n905 | (~Pi21 & ~n1229));
  assign n3876 = ~Pi20 & (~n905 | (~Pi21 & ~n1220));
  assign n3877 = Pi16 | ~Pi15;
  assign n3878 = Pi20 & (~n905 | (~Pi21 & ~n954));
  assign n3879 = ~Pi20 & (~n905 | (~Pi21 & ~n930));
  assign n3880 = ~n901 | n978 | n3878 | n3879;
  assign n3881 = Pi20 & (~n905 | (~Pi21 & ~n1152));
  assign n3882 = ~Pi20 & (~n905 | (~Pi21 & ~n1138));
  assign n3883 = ~n901 | n1211 | n3881 | n3882;
  assign n3884 = ~Pi16 | Pi15;
  assign n3885 = Pi20 & (~n905 | (~Pi21 & ~n1029));
  assign n3886 = ~Pi20 & (~n905 | (~Pi21 & ~n1022));
  assign n3887 = ~n901 | n1040 | n3885 | n3886;
  assign n3888 = Pi20 & (~n905 | (~Pi21 & ~n1267));
  assign n3889 = ~Pi20 & (~n905 | (~Pi21 & ~n1260));
  assign n3890 = ~n901 | n1290 | n3888 | n3889;
  assign n3891 = ~Pi16 | ~Pi15;
  assign n3892 = Ni10 | ~n3327;
  assign n3893 = ~Pi19 | n3857;
  assign n3894 = Pi16 | n3864;
  assign n3895 = Pi16 | n1322;
  assign n3896 = Ni6 | Ni4 | Ni5;
  assign n3897 = Ni11 | Ni10;
  assign n3898 = n1446 & Ni11;
  assign n3899 = n3848 | n3761;
  assign n3900 = ~n3761 | n3848;
  assign n3901 = n3857 | n3761;
  assign n3902 = n3859 | n3761;
  assign n3903 = ~n3761 | n3859;
  assign n3904 = Pi27 | n1495;
  assign n3905 = Pi27 | n1497;
  assign n3906 = ~Pi27 | n1495;
  assign n3907 = ~Pi27 | n1497;
  assign n3908 = Pi27 | n3857;
  assign n3909 = Pi27 | n3859;
  assign n3910 = ~Pi27 | n3857;
  assign n3911 = ~Pi27 | n3859;
  assign n3912 = Ni13 | Ni14;
  assign n3913 = n3848 | n789;
  assign n3914 = ~n789 | n3848;
  assign n3915 = n3857 | n789;
  assign n3916 = n3859 | n789;
  assign n3917 = ~n789 | n3859;
  assign n3918 = n3799 | n3798;
  assign n3919 = Ni11 | ~Ni12;
  assign n3920 = Pi27 | n1923;
  assign n3921 = ~Pi27 | n1923;
  assign n3922 = Pi27 | n1929;
  assign n3923 = ~Pi27 | n2372;
  assign n3924 = n1923 | n789;
  assign n3925 = ~n789 | n1923;
  assign n3926 = n2372 | n789;
  assign n3927 = n1314 | n789;
  assign n3928 = Ni13 | n3919;
  assign n3929 = n1923 | n3761;
  assign n3930 = n1923 | ~n3761;
  assign n3931 = n2372 | n3761;
  assign n3932 = n1314 | n3761;
  assign n3933 = n3848 | n788;
  assign n3934 = ~n788 | n3848;
  assign n3935 = n3857 | n788;
  assign n3936 = ~n788 | n3857;
  assign n3937 = Ni10 | n3768;
  assign n3938 = ~Pi24 | n1495;
  assign n3939 = ~Pi24 | n1497;
  assign n3940 = Pi24 | n3857;
  assign n3941 = Pi24 | n3859;
  assign n3942 = ~Pi24 | n3857;
  assign n3943 = ~Pi24 | n3859;
  assign n3944 = Pi15 | n3327;
  assign n3945 = n3848 | n795;
  assign n3946 = ~n795 | n3848;
  assign n3947 = n3857 | n795;
  assign n3948 = ~n795 | n3857;
  assign n3949 = ~Pi25 | n2079;
  assign n3950 = ~n18 | Ni33;
  assign n3951 = ~Pi25 | Ni34 | n1539 | n3950;
  assign n3952 = n2254 | n2079;
  assign n3953 = ~Ni34 | Ni33;
  assign n3954 = n3952 | n3953;
  assign n3955 = n3954 & ~n792 & n2085;
  assign n3956 = Ni32 & Ni33;
  assign n3957 = ~Ni10 | ~Ni9;
  assign n3958 = Ni31 | n3795;
  assign n3959 = Ni39 | n3852;
  assign n3960 = n1241 | ~Ni38;
  assign n3961 = n3852 | ~Ni39;
  assign n3962 = n2389 | ~Ni38;
  assign n3963 = n2518 & n2430 & n2431;
  assign n3964 = n2523 & n2430 & n2444;
  assign n3965 = n2427 & n2430 & n2431;
  assign n3966 = n2442 & n2430 & n2444;
  assign n3967 = ~Pi26 | Pi24;
  assign n3968 = ~Ni37 | ~Ni38;
  assign n3969 = Ni32 | ~Ni40;
  assign n3970 = Ni33 | n3751;
  assign n3971 = ~Ni33 | n3751;
  assign n3972 = Ni32 | ~Ni41;
  assign n3973 = Ni31 & Ni33;
  assign n3974 = Ni38 | n3198;
  assign n3975 = Ni33 | n1539;
  assign n3976 = Ni38 | n3200;
  assign n3977 = n3834 | n3835;
  assign n3978 = ~Pi17 | Pi16;
  assign n3979 = ~Pi17 | ~Pi16;
  assign n3980 = ~Ni30 | n3701;
  assign n3981 = ~Pi27 & n3669;
  assign n3982 = n3688 | ~n3957;
  assign n3983 = n3704 | Ni6 | ~Ni5;
  assign n3984 = ~Ni32 & Ni30;
  assign n3985 = n3707 | n2393;
  assign n3986 = n2403 | Ni7 | n3707;
  assign n3987 = ~n4673 & (~n18 | ~n3707);
  assign n1026_1 = ~n3987;
  assign n3989 = (~Ni10 & ~n1944) | (~n1718 & (Ni10 | ~n1944));
  assign n3990 = (Pi15 & n4678) | (n4677 & (~Pi15 | n4678));
  assign n3991 = ~n4687 & (~Pi17 | ~n4171 | ~n4172);
  assign n3992 = ~n4686 & (Ni10 | ~n4195 | ~n4197);
  assign n3993 = n3797 & (n1540 | n2254) & ~n3800;
  assign n3994 = (~Ni10 | n2370) & n4700;
  assign n3995 = ~n4701 & (~Pi17 | (n4375 & n4376));
  assign n3996 = (~Ni10 & ~n3060) | (~n2867 & (Ni10 | ~n3060));
  assign n3997 = (Pi15 & n4715) | (n4714 & (~Pi15 | n4715));
  assign n3998 = ~n4725 & (~Pi17 | ~n4434 | ~n4435);
  assign n3999 = ~Pi22 & ~n3812 & (~Pi27 | ~n3819);
  assign n4000 = ~n4713 & (~Ni14 | ~n4448 | ~n4449);
  assign n4001 = (n4196 | n3060) & (Ni11 | n3061);
  assign n4002 = ~n3175 & n4001 & (n3928 | ~n4000);
  assign n4003 = (~Pi23 & n4724) | (~n2626 & (Pi23 | n4724));
  assign n4004 = (~n788 & ~n3816) | (~n2630 & (n788 | ~n3816));
  assign n4005 = (Pi24 & ~n3816) | (~n2630 & (~Pi24 | ~n3816));
  assign n4006 = (Pi24 & n4710) | (~n2626 & (~Pi24 | n4710));
  assign n4007 = (Pi24 & n4712) | (~n2636 & (~Pi24 | n4712));
  assign n4008 = (Pi23 & n4724) | (~n2626 & (~Pi23 | n4724));
  assign n4009 = (~n795 & ~n3816) | (~n2630 & (n795 | ~n3816));
  assign n4010 = n3896 & (n3178 | n3179 | ~n4589);
  assign n4011 = n3969 & (~Pi23 | n3970);
  assign n4012 = n3187 & n4011 & (~Ni40 | n3971);
  assign n4013 = n4728 & (n2393 | (n4590 & n3827));
  assign n4014 = (~n2403 & n4729) | (~n4013 & (n2403 | n4729));
  assign n4015 = (~Pi24 | n3970) & n3972;
  assign n4016 = n3189 & n4015 & (~Ni41 | n3971);
  assign n4017 = n4730 & (n2393 | (n4591 & n3831));
  assign n4018 = (~n2403 & n4731) | (~n4017 & (n2403 | n4731));
  assign n4019 = ~n3773 & (n3737 | (n3472 & n4607));
  assign n4020 = ~n3475 & (n3895 | (n3472 & n4605));
  assign n4021 = ~n3474 & (n3740 | (n3472 & n4603));
  assign n4022 = n4608 & (n3894 | (n4602 & n3472));
  assign n4023 = n4022 & n4021 & n4019 & n4020;
  assign n4024 = ~n3773 & (n3737 | (n3472 & n4628));
  assign n4025 = ~n3534 & (n3895 | (n3472 & n4626));
  assign n4026 = ~n3533 & (n3740 | (n3472 & n4624));
  assign n4027 = n4629 & (n3894 | (n4623 & n3472));
  assign n4028 = n4027 & n4026 & n4024 & n4025;
  assign n4029 = ~n4749 & (~Ni10 | (~n4747 & ~n4748));
  assign n4030 = (~Pi20 & n3324) | (n3315 & (Pi20 | n3324));
  assign n4031 = (~Pi20 & n3287) | (n3265 & (Pi20 | n3287));
  assign n4032 = n3805 & (n3328 | n3329 | n3330);
  assign n4033 = ~Ni4 | n780 | n3693;
  assign n4034 = n4033 & ~n4751 & (Ni5 | ~n3692);
  assign n4035 = ~n4755 & (~Ni4 | ~Ni2);
  assign n1081 = ~n4035;
  assign n4037 = n3957 | ~Ni8 | ~Ni7;
  assign n4038 = n3688 & (n795 | ~Ni10 | n2074);
  assign n4039 = n4037 & n4038 & (Ni7 | ~n3957);
  assign n4040 = (~n3707 & ~n4039) | (~Ni7 & (n3707 | ~n4039));
  assign n1066_1 = ~n4040;
  assign n4042 = (~Ni10 & (n3707 | n3721)) | (~n3707 & n3721);
  assign n1051 = ~n4042;
  assign n4044 = (Ni11 & (n1542 | n3727)) | (n1542 & ~n3727);
  assign n4045 = n1543 & n4044 & (n1446 | n3761);
  assign n4046 = (~n3707 & ~n4045) | (~Ni11 & (n3707 | ~n4045));
  assign n1046_1 = ~n4046;
  assign n4048 = ~n4757 & (Ni12 | n3707 | n3727);
  assign n1041_1 = ~n4048;
  assign n4050 = ~n4759 & (~n3733 | ~Ni42 | ~Ni39);
  assign n4051 = (~Pi26 | n4760) & n4761;
  assign n4052 = (~Pi23 | n4762) & n4763;
  assign n4053 = (n848 | n3857) & (n879 | n3859);
  assign n4054 = (n940 | n3857) & (n964 | n3859);
  assign n4055 = n1055 | (~Ni37 & n817);
  assign n4056 = n1051_1 | (~Ni37 & n817);
  assign n4057 = n1070 | (~Ni37 & n853);
  assign n4058 = n1067 | (~Ni37 & n853);
  assign n4059 = (n1060 | n3857) & (n1074 | n3859);
  assign n4060 = (n1101 | n3857) & (n1126 | n3859);
  assign n4061 = n1140 | (~Ni37 & n817);
  assign n4062 = n1137 | (~Ni37 & n817);
  assign n4063 = n1154 | (~Ni37 & n853);
  assign n4064 = n1151 | (~Ni37 & n853);
  assign n4065 = (n1144 | n3857) & (n1158 | n3859);
  assign n4066 = (n1182 | n3857) & (n1206 | n3859);
  assign n4067 = (n911 | ~n3772) & (n980 | ~n2345);
  assign n4068 = n975 | n1497;
  assign n4069 = n4068 & (n3894 | (~n3863 & n4053));
  assign n4070 = ~n1307 & (n3895 | (~n1295 & n4060));
  assign n4071 = n3850 | Ni32 | n884;
  assign n4072 = n3850 | Ni32 | n967;
  assign n4073 = (n999 | n3857) & (n1008 | n3859);
  assign n4074 = (n1026 | n3857) & (n1033 | n3859);
  assign n4075 = (n1226 | n3857) & (n1233 | n3859);
  assign n4076 = (n1245 | n3857) & (n1253 | n3859);
  assign n4077 = (n1264 | n3857) & (n1271 | n3859);
  assign n4078 = (n1278 | n3857) & (n1285 | n3859);
  assign n4079 = (n1017 | ~n3772) & (n1042 | ~n2345);
  assign n4080 = n1037 | n1497;
  assign n4081 = n4080 & (n3894 | (~n3873 & n4073));
  assign n4082 = ~n1300 & (n3895 | (~n1297 & n4076));
  assign n4083 = (n1102 | n3893) & (n1127 | n2109);
  assign n4084 = n4083 & (n1061_1 | n1408);
  assign n4085 = (n914 | n1075) & (Pi19 | ~n1306);
  assign n4086 = (n1246 | n3893) & (n1254 | n2109);
  assign n4087 = n4086 & (n1227 | n1408);
  assign n4088 = (n914 | n1234) & (Pi19 | ~n1299);
  assign n4089 = (n1215 | n3884) & (n1294 | n3891);
  assign n4090 = (n915 | n3870) & (n1020 | n3877);
  assign n4091 = (n983 | n3884) & (n1045 | n3891);
  assign n4092 = (n848 | n3858) & (n879 | n3860);
  assign n4093 = (n1060 | n3858) & (n1074 | n3860);
  assign n4094 = (n1101 | n3858) & (n1126 | n3860);
  assign n4095 = (n898 | n1923) & (n911 | ~n3184);
  assign n4096 = Pi25 | n3847;
  assign n4097 = (n999 | n3858) & (n1008 | n3860);
  assign n4098 = (n1226 | n3858) & (n1233 | n3860);
  assign n4099 = (n1245 | n3858) & (n1253 | n3860);
  assign n4100 = (n1013 | n1923) & (n1017 | ~n3184);
  assign n4101 = (n940 | n3858) & (n964 | n3860);
  assign n4102 = (n1144 | n3858) & (n1158 | n3860);
  assign n4103 = (n1182 | n3858) & (n1206 | n3860);
  assign n4104 = (n976 | n1923) & (n980 | ~n3184);
  assign n4105 = (n1026 | n3858) & (n1033 | n3860);
  assign n4106 = (n1264 | n3858) & (n1271 | n3860);
  assign n4107 = (n1278 | n3858) & (n1285 | n3860);
  assign n4108 = (n1038 | n1923) & (n1042 | ~n3184);
  assign n4109 = (n1332 | n3870) & (n1350 | n3877);
  assign n4110 = (n1323 | n3884) & (n1341 | n3891);
  assign n4111 = (n1937 | n3894) & (n1700 | n3740);
  assign n4112 = n4111 & (n1961 | n2272);
  assign n4113 = (n1958 | n3895) & (n1708 | n3743);
  assign n4114 = n4113 & (n1709 | n3737);
  assign n4115 = (n1704 | n3894) & (n1706 | n3740);
  assign n4116 = n4115 & (n1711 | n2272);
  assign n4117 = (n1712 | n3895) & (n1714 | n3743);
  assign n4118 = n4117 & (n1715 | n3737);
  assign n4119 = n1759 & n1404;
  assign n4120 = n1769 & n1400;
  assign n4121 = n1829 & n1429;
  assign n4122 = n1839 & n1425;
  assign n4123 = n1723 & n1417;
  assign n4124 = n1734 & n1413;
  assign n4125 = n1794 & n1441;
  assign n4126 = n1804 & n1437;
  assign n4127 = (n1687 | n3870) & (n1695 | n3877);
  assign n4128 = (n1691 | n3884) & (n1699 | n3891);
  assign n4129 = n1785 & n1361;
  assign n4130 = n1855 & n1380;
  assign n4131 = n1750 & n1371;
  assign n4132 = n1820 & n1389;
  assign n4133 = (n1674 | n3870) & (n1680 | n3877);
  assign n4134 = (n1677 | n3884) & (n1683 | n3891);
  assign n4135 = n1518 & n1357;
  assign n4136 = n1530 & n1367;
  assign n4137 = (n4136 | n3858) & (n1373 | n3860);
  assign n4138 = n1516 & n1400;
  assign n4139 = (n1407 | n3858) & (n4138 | n3860);
  assign n4140 = n1510 & n1402;
  assign n4141 = n1512 & n1404;
  assign n4142 = (n4140 | n3858) & (n4141 | n3860);
  assign n4143 = n1528 & n1413;
  assign n4144 = (n1420 | n3858) & (n4143 | n3860);
  assign n4145 = n1522 & n1415;
  assign n4146 = n1524 & n1417;
  assign n4147 = (n4145 | n3858) & (n4146 | n3860);
  assign n4148 = (n1926 | n1923) & (n1938 | n3894);
  assign n4149 = n1478 & n1376;
  assign n4150 = n1490 & n1385;
  assign n4151 = (n4150 | n3858) & (n1391 | n3860);
  assign n4152 = n1476 & n1425;
  assign n4153 = (n1432 | n3858) & (n4152 | n3860);
  assign n4154 = n1470 & n1427;
  assign n4155 = n1472 & n1429;
  assign n4156 = (n4154 | n3858) & (n4155 | n3860);
  assign n4157 = n1488 & n1437;
  assign n4158 = (n1444 | n3858) & (n4157 | n3860);
  assign n4159 = n1482 & n1439;
  assign n4160 = n1484 & n1441;
  assign n4161 = (n4159 | n3858) & (n4160 | n3860);
  assign n4162 = (n1922 | n1923) & (n1930 | n3894);
  assign n4163 = (n1961 | n1701) & (n1958 | n1702);
  assign n4164 = n4163 & (n1713 | n3877);
  assign n4165 = (n1710 | n3884) & (n1716 | n3891);
  assign n4166 = (n1937 | n1701) & (n1360 | n1702);
  assign n4167 = n4166 & (n1705 | n3877);
  assign n4168 = (n1703 | n3884) & (n1707 | n3891);
  assign n4169 = (n1409 | n3870) & (n1433 | n3877);
  assign n4170 = (n1421 | n3884) & (n1445 | n3891);
  assign n4171 = (n1365 | n3870) & (n1383 | n3877);
  assign n4172 = (n1374 | n3884) & (n1392 | n3891);
  assign n4173 = n1786 | n3924;
  assign n4174 = n2026 | ~n3184;
  assign n4175 = n1856 | n3924;
  assign n4176 = n1751 | n3924;
  assign n4177 = n1821 | n3924;
  assign n4178 = (n2045 | n3870) & (n2063 | n3877);
  assign n4179 = (n2036 | n3884) & (n2054 | n3891);
  assign n4180 = n1360 | n3920;
  assign n4181 = n1987 | ~n3184;
  assign n4182 = n1379 | n3920;
  assign n4183 = n1370 | n3920;
  assign n4184 = n1388 | n3920;
  assign n4185 = (n2006 | n3870) & (n2024 | n3877);
  assign n4186 = (n1997 | n3884) & (n2015 | n3891);
  assign n4187 = n1786 | n3929;
  assign n4188 = n1946 | ~n3184;
  assign n4189 = n1856 | n3929;
  assign n4190 = n1751 | n3929;
  assign n4191 = n1821 | n3929;
  assign n4192 = (n1967 | n3870) & (n1985 | n3877);
  assign n4193 = (n1956 | n3884) & (n1976 | n3891);
  assign n4194 = n3928 | n4675 | n4676;
  assign n4195 = n4194 & (n3677 | (n4193 & n4192));
  assign n4196 = n1452 & ~n3898;
  assign n4197 = (n4196 | n1944) & (Ni11 | n1945);
  assign n4198 = n1787 | n3899;
  assign n4199 = n1455 | ~n3184;
  assign n4200 = n1857 | n3899;
  assign n4201 = n1752 | n3899;
  assign n4202 = n1822 | n3899;
  assign n4203 = (n1783 | n3908) & (n1673 | n3909);
  assign n4204 = (n1777 | n3910) & (n1780 | n3911);
  assign n4205 = (n1748 | n3908) & (n1676 | n3909);
  assign n4206 = (n1742 | n3910) & (n1745 | n3911);
  assign n4207 = (n1686 | n3908) & (n4120 | n3909);
  assign n4208 = (n1768 | n3910) & (n1771 | n3911);
  assign n4209 = (n1764 | n3908) & (n4119 | n3909);
  assign n4210 = (n1758 | n3910) & (n1761 | n3911);
  assign n4211 = (n1690 | n3908) & (n4124 | n3909);
  assign n4212 = (n1733 | n3910) & (n1736 | n3911);
  assign n4213 = (n1728 | n3908) & (n4123 | n3909);
  assign n4214 = (n1722 | n3910) & (n1725 | n3911);
  assign n4215 = (n4129 | n3904) & (n4131 | n3905);
  assign n4216 = n1752 | n3907;
  assign n4217 = n4216 & (n3894 | (n4204 & n4203));
  assign n4218 = n4217 & (n3740 | (n4206 & n4205));
  assign n4219 = ~n1862 & (n3895 | (n4209 & n4210));
  assign n4220 = n4219 & (n3743 | (n4212 & n4211));
  assign n4221 = n1552 & (n3737 | (n4214 & n4213));
  assign n4222 = (n1853 | n3908) & (n1679 | n3909);
  assign n4223 = (n1847 | n3910) & (n1850 | n3911);
  assign n4224 = (n1818 | n3908) & (n1682 | n3909);
  assign n4225 = (n1812 | n3910) & (n1815 | n3911);
  assign n4226 = (n1694 | n3908) & (n4122 | n3909);
  assign n4227 = (n1838 | n3910) & (n1841 | n3911);
  assign n4228 = (n1834 | n3908) & (n4121 | n3909);
  assign n4229 = (n1828 | n3910) & (n1831 | n3911);
  assign n4230 = (n1698 | n3908) & (n4126 | n3909);
  assign n4231 = (n1803 | n3910) & (n1806 | n3911);
  assign n4232 = (n1799 | n3908) & (n4125 | n3909);
  assign n4233 = (n1793 | n3910) & (n1796 | n3911);
  assign n4234 = (n4130 | n3904) & (n4132 | n3905);
  assign n4235 = n1822 | n3907;
  assign n4236 = n4235 & (n3894 | (n4223 & n4222));
  assign n4237 = n4236 & (n3740 | (n4225 & n4224));
  assign n4238 = ~n1861 & (n3895 | (n4228 & n4229));
  assign n4239 = n4238 & (n3743 | (n4231 & n4230));
  assign n4240 = n1552 & (n3737 | (n4233 & n4232));
  assign n4241 = n1787 | n3913;
  assign n4242 = ~n3184 | ~n3918;
  assign n4243 = n1857 | n3913;
  assign n4244 = n1752 | n3913;
  assign n4245 = n1822 | n3913;
  assign n4246 = (n1790 | n3870) & (n1860 | n3877);
  assign n4247 = (n1755 | n3884) & (n1825 | n3891);
  assign n4248 = (n1917 | n3677) & (n1718 | ~n3898);
  assign n4249 = (~Ni14 & n4300) | (n1552 & (Ni14 | n4300));
  assign n4250 = n3804 & (~Pi23 | n4249);
  assign n4251 = n1507 | n3933;
  assign n4252 = ~n794 | ~n3184;
  assign n4253 = n1466 | n3933;
  assign n4254 = n1509 | n3933;
  assign n4255 = n1469 | n3933;
  assign n4256 = (n1578 | n3870) & (n1602 | n3877);
  assign n4257 = (n1566 | n3884) & (n1590 | n3891);
  assign n4258 = (n1540 | n2254) & (Pi24 | n3801);
  assign n4259 = (n4135 | n3940) & (n1364 | n3941);
  assign n4260 = (n1519 | n3942) & (n1521 | n3943);
  assign n4261 = (n4136 | n3940) & (n1373 | n3941);
  assign n4262 = (n1531 | n3942) & (n1533 | n3943);
  assign n4263 = (n1407 | n3940) & (n4138 | n3941);
  assign n4264 = (n1515 | n3942) & (n1517 | n3943);
  assign n4265 = (n4140 | n3940) & (n4141 | n3941);
  assign n4266 = (n1511 | n3942) & (n1513 | n3943);
  assign n4267 = (n1420 | n3940) & (n4143 | n3941);
  assign n4268 = (n1527 | n3942) & (n1529 | n3943);
  assign n4269 = (n4145 | n3940) & (n4146 | n3941);
  assign n4270 = (n1523 | n3942) & (n1525 | n3943);
  assign n4271 = (n1507 | n3938) & (n1509 | n3939);
  assign n4272 = ~n1537 & (n3740 | (n4261 & n4262));
  assign n4273 = n4271 & n4272 & (Pi24 | n1536);
  assign n4274 = ~n1538 & (n3895 | (n4265 & n4266));
  assign n4275 = n4274 & (n3743 | (n4268 & n4267));
  assign n4276 = n1460 & (n3737 | (n4270 & n4269));
  assign n4277 = (n4149 | n3940) & (n1382 | n3941);
  assign n4278 = (n1479 | n3942) & (n1481 | n3943);
  assign n4279 = (n4150 | n3940) & (n1391 | n3941);
  assign n4280 = (n1491 | n3942) & (n1493 | n3943);
  assign n4281 = (n1432 | n3940) & (n4152 | n3941);
  assign n4282 = (n1475 | n3942) & (n1477 | n3943);
  assign n4283 = (n4154 | n3940) & (n4155 | n3941);
  assign n4284 = (n1471 | n3942) & (n1473 | n3943);
  assign n4285 = (n1444 | n3940) & (n4157 | n3941);
  assign n4286 = (n1487 | n3942) & (n1489 | n3943);
  assign n4287 = (n4159 | n3940) & (n4160 | n3941);
  assign n4288 = (n1483 | n3942) & (n1485 | n3943);
  assign n4289 = (n1466 | n3938) & (n1469 | n3939);
  assign n4290 = ~n1500 & (n3895 | (n4283 & n4284));
  assign n4291 = (n1505 | n2367) & (n1462 | n1544);
  assign n4292 = n3804 & (Pi23 | n4249);
  assign n4293 = n1507 | n3945;
  assign n4294 = ~n796 | ~n3184;
  assign n4295 = n1466 | n3945;
  assign n4296 = n1509 | n3945;
  assign n4297 = n1469 | n3945;
  assign n4298 = (n1637 | n3870) & (n1661 | n3877);
  assign n4299 = (n1625 | n3884) & (n1649 | n3891);
  assign n4300 = n2025 | n2254;
  assign n4301 = ~n2386 & (n2382 | n3894);
  assign n4302 = (n2385 | n3740) & (n2381 | n2272);
  assign n4303 = (n2380 | n3895) & (n2384 | n3743);
  assign n4304 = (n2378 | n3740) & (n2374 | n2272);
  assign n4305 = ~n2379 & n4304 & (n2375 | n3894);
  assign n4306 = (n2373 | n3895) & (n2377 | n3743);
  assign n4307 = n2371 & n4306 & (n2376 | n3737);
  assign n4308 = (n2196 | n3949) & (~n1081_1 | n3951);
  assign n4309 = n2105 & (~Pi25 | n2313);
  assign n4310 = (n2228 | n3949) & (~n1235 | n3951);
  assign n4311 = n2120 & (~Pi25 | n2277);
  assign n4312 = (n2212 | n3949) & (~n1165 | n3951);
  assign n4313 = n2113 & (~Pi25 | n2320);
  assign n4314 = (n2244 | n3949) & (~n1273 | n3951);
  assign n4315 = n2127 & (~Pi25 | n2284);
  assign n4316 = (n2203 | n3870) & (n2235 | n3877);
  assign n4317 = (n2219 | n3884) & (n2251 | n3891);
  assign n4318 = (n2145 | n3870) & (n2173 | n3877);
  assign n4319 = (n2159 | n3884) & (n2187 | n3891);
  assign n4320 = (n2347 | n3847) & (n2140 | n3952);
  assign n4321 = (n2348 | n3847) & (n2154 | n3952);
  assign n4322 = (n2359 | n3847) & (n2132 | n3952);
  assign n4323 = (n2362 | n3847) & (n2146 | n3952);
  assign n4324 = (n2357 | n3847) & (n2188 | n3952);
  assign n4325 = (n2358 | n3847) & (n2196 | n3952);
  assign n4326 = (n2360 | n3847) & (n2204 | n3952);
  assign n4327 = (n2361 | n3847) & (n2212 | n3952);
  assign n4328 = ~n2363 & (n3740 | (n3955 & n4323));
  assign n4329 = n4328 & (n2272 | (n4324 & n3955));
  assign n4330 = ~n2364 & (n3895 | (n3955 & n4325));
  assign n4331 = n4330 & (n3737 | (n4327 & n3955));
  assign n4332 = (n2351 | n3847) & (n2136 | n3952);
  assign n4333 = (n2354 | n3847) & (n2150 | n3952);
  assign n4334 = (n2349 | n3847) & (n2192 | n3952);
  assign n4335 = (n2350 | n3847) & (n2197 | n3952);
  assign n4336 = (n2352 | n3847) & (n2208 | n3952);
  assign n4337 = (n2353 | n3847) & (n2213 | n3952);
  assign n4338 = ~n2355 & (n3740 | (n3955 & n4333));
  assign n4339 = n4338 & (n2272 | (n4334 & n3955));
  assign n4340 = ~n2356 & (n3895 | (n3955 & n4335));
  assign n4341 = n4340 & (n3737 | (n4337 & n3955));
  assign n4342 = ~n2365 & (~n3772 | (n3955 & n4320));
  assign n4343 = (n2327 | n3847) & (n2168 | n3952);
  assign n4344 = (n2328 | n3847) & (n2182 | n3952);
  assign n4345 = (n2339 | n3847) & (n2160 | n3952);
  assign n4346 = (n2342 | n3847) & (n2174 | n3952);
  assign n4347 = (n2337 | n3847) & (n2220 | n3952);
  assign n4348 = (n2338 | n3847) & (n2228 | n3952);
  assign n4349 = (n2340 | n3847) & (n2236 | n3952);
  assign n4350 = (n2341 | n3847) & (n2244 | n3952);
  assign n4351 = ~n2343 & (n3740 | (n3955 & n4346));
  assign n4352 = n4351 & (n2272 | (n4347 & n3955));
  assign n4353 = ~n2344 & (n3895 | (n3955 & n4348));
  assign n4354 = n4353 & (n3737 | (n4350 & n3955));
  assign n4355 = (n2331 | n3847) & (n2164 | n3952);
  assign n4356 = (n2334 | n3847) & (n2178 | n3952);
  assign n4357 = (n2329 | n3847) & (n2224 | n3952);
  assign n4358 = (n2330 | n3847) & (n2229 | n3952);
  assign n4359 = (n2332 | n3847) & (n2240 | n3952);
  assign n4360 = (n2333 | n3847) & (n2245 | n3952);
  assign n4361 = ~n2335 & (n3740 | (n3955 & n4356));
  assign n4362 = n4361 & (n2272 | (n4357 & n3955));
  assign n4363 = ~n2336 & (n3895 | (n3955 & n4358));
  assign n4364 = n4363 & (n3737 | (n4360 & n3955));
  assign n4365 = ~n2346 & (~n3772 | (n3955 & n4343));
  assign n4366 = (n2314 | n3895) & (n2318 | n3743);
  assign n4367 = (n2298 | n3895) & (n2302 | n3743);
  assign n4368 = (n2292 | ~n3772) & (n2294 | ~n2345);
  assign n4369 = (n2278 | n3895) & (n2282 | n3743);
  assign n4370 = (n2261 | n3895) & (n2265 | n3743);
  assign n4371 = ~n3327 | n4698 | n4699;
  assign n4372 = (~Pi20 & n2326) | (n2309 & (Pi20 | n2326));
  assign n4373 = (n2110 | n3870) & (n2124 | n3877);
  assign n4374 = (n2117 | n3884) & (n2131 | n3891);
  assign n4375 = (n2087 | n3870) & (n2097 | n3877);
  assign n4376 = (n2092 | n3884) & (n2102 | n3891);
  assign n4377 = (n1238 | n3958) & (~Pi23 | n3807);
  assign n4378 = (n886 | n3958) & (~Pi24 | n3807);
  assign n4379 = (Pi15 | n2414) & (n2413 | ~n3846);
  assign n4380 = (n2851 | n3894) & (n2853 | n3740);
  assign n4381 = n4380 & (n2857 | n2272);
  assign n4382 = (n2858 | n3895) & (n2860 | n3743);
  assign n4383 = n4382 & (n2861 | n3737);
  assign n4384 = (n3046 | n3894) & (n2855 | n3740);
  assign n4385 = n4384 & (n3094 | n2272);
  assign n4386 = (n3091 | n3895) & (n2863 | n3743);
  assign n4387 = n4386 & (n2864 | n3737);
  assign n4388 = n2822 & n2542;
  assign n4389 = n2820 & n2527;
  assign n4390 = n2838 & n2592;
  assign n4391 = n2836 & n2582;
  assign n4392 = n2830 & n2568;
  assign n4393 = n2828 & n2554;
  assign n4394 = n2846 & n2616;
  assign n4395 = n2844 & n2606;
  assign n4396 = (n2826 | n3870) & (n2842 | n3877);
  assign n4397 = (n2834 | n3884) & (n2850 | n3891);
  assign n4398 = n2797 & n2457;
  assign n4399 = n2809 & n2497;
  assign n4400 = n2803 & n2480;
  assign n4401 = n2815 & n2514;
  assign n4402 = (n2800 | n3870) & (n2812 | n3877);
  assign n4403 = (n2806 | n3884) & (n2818 | n3891);
  assign n4404 = n2436 & n2440;
  assign n4405 = n2464 & n2467;
  assign n4406 = (n4405 | n3858) & (n2482 | n3860);
  assign n4407 = (n2545 | n3858) & (n2721 | n3860);
  assign n4408 = n2532 & n2535;
  assign n4409 = (n4408 | n3858) & (n2718 | n3860);
  assign n4410 = (n2571 | n3858) & (n2710 | n3860);
  assign n4411 = n2558 & n2561;
  assign n4412 = (n4411 | n3858) & (n2706 | n3860);
  assign n4413 = (n3043 | n1923) & (n3054 | n3894);
  assign n4414 = n2485 & n2488;
  assign n4415 = n2502 & n2505;
  assign n4416 = (n4415 | n3858) & (n2516 | n3860);
  assign n4417 = (n2595 | n3858) & (n2743 | n3860);
  assign n4418 = n2584 & n2587;
  assign n4419 = (n4418 | n3858) & (n2740 | n3860);
  assign n4420 = (n2619 | n3858) & (n2732 | n3860);
  assign n4421 = n2608 & n2611;
  assign n4422 = (n4421 | n3858) & (n2729 | n3860);
  assign n4423 = (n3040 | n1923) & (n3047 | n3894);
  assign n4424 = (n3094 | n1701) & (n3091 | n1702);
  assign n4425 = n4424 & (n2859 | n3870);
  assign n4426 = (n2862 | n3884) & (n2865 | n3891);
  assign n4427 = (n3046 | n1701) & (n2496 | n1702);
  assign n4428 = n4427 & (n2852 | n3870);
  assign n4429 = (n2854 | n3884) & (n2856 | n3891);
  assign n4430 = (n3061 | n3897) & (~n1543 | ~n3996);
  assign n4431 = ~n2074 & (~n4430 | (~n2070 & ~n2868));
  assign n4432 = (n2546 | n3870) & (n2596 | n3877);
  assign n4433 = (n2572 | n3884) & (n2620 | n3891);
  assign n4434 = (n2460 | n3870) & (n2500 | n3877);
  assign n4435 = (n2483 | n3884) & (n2517 | n3891);
  assign n4436 = n2920 | n3924;
  assign n4437 = n3138 | ~n3184;
  assign n4438 = n2976 | n3924;
  assign n4439 = n2892 | n3924;
  assign n4440 = n2948 | n3924;
  assign n4441 = (n3156 | n3870) & (n3174 | n3877);
  assign n4442 = (n3147 | n3884) & (n3165 | n3891);
  assign n4443 = n2456 | n3920;
  assign n4444 = n3101 | ~n3184;
  assign n4445 = n2496 | n3920;
  assign n4446 = n2479 | n3920;
  assign n4447 = n2513 | n3920;
  assign n4448 = (n3119 | n3870) & (n3137 | n3877);
  assign n4449 = (n3110 | n3884) & (n3128 | n3891);
  assign n4450 = n2920 | n3929;
  assign n4451 = n3062 | ~n3184;
  assign n4452 = n2976 | n3929;
  assign n4453 = n2892 | n3929;
  assign n4454 = n2948 | n3929;
  assign n4455 = (n3080 | n3870) & (n3100 | n3877);
  assign n4456 = (n3071 | n3884) & (n3089 | n3891);
  assign n4457 = n2921 | n3899;
  assign n4458 = n2634 | ~n3184;
  assign n4459 = n2977 | n3899;
  assign n4460 = n2893 | n3899;
  assign n4461 = n2949 | n3899;
  assign n4462 = (n2918 | n3908) & (n2799 | n3909);
  assign n4463 = (n2913 | n3910) & (n2915 | n3911);
  assign n4464 = (n2890 | n3908) & (n2805 | n3909);
  assign n4465 = (n2885 | n3910) & (n2887 | n3911);
  assign n4466 = (n2825 | n3908) & (n4389 | n3909);
  assign n4467 = (n2906 | n3910) & (n2908 | n3911);
  assign n4468 = (n2903 | n3908) & (n4388 | n3909);
  assign n4469 = (n2898 | n3910) & (n2900 | n3911);
  assign n4470 = (n2833 | n3908) & (n4393 | n3909);
  assign n4471 = (n2878 | n3910) & (n2880 | n3911);
  assign n4472 = (n2875 | n3908) & (n4392 | n3909);
  assign n4473 = (n2870 | n3910) & (n2872 | n3911);
  assign n4474 = (n4398 | n3904) & (n4400 | n3905);
  assign n4475 = n2893 | n3907;
  assign n4476 = n4475 & (n3894 | (n4463 & n4462));
  assign n4477 = n4476 & (n3740 | (n4465 & n4464));
  assign n4478 = ~n2982 & (n3895 | (n4468 & n4469));
  assign n4479 = n4478 & (n3743 | (n4471 & n4470));
  assign n4480 = n2628 & (n3737 | (n4473 & n4472));
  assign n4481 = (n2974 | n3908) & (n2811 | n3909);
  assign n4482 = (n2969 | n3910) & (n2971 | n3911);
  assign n4483 = (n2946 | n3908) & (n2817 | n3909);
  assign n4484 = (n2941 | n3910) & (n2943 | n3911);
  assign n4485 = (n2841 | n3908) & (n4391 | n3909);
  assign n4486 = (n2962 | n3910) & (n2964 | n3911);
  assign n4487 = (n2959 | n3908) & (n4390 | n3909);
  assign n4488 = (n2954 | n3910) & (n2956 | n3911);
  assign n4489 = (n2849 | n3908) & (n4395 | n3909);
  assign n4490 = (n2934 | n3910) & (n2936 | n3911);
  assign n4491 = (n2931 | n3908) & (n4394 | n3909);
  assign n4492 = (n2926 | n3910) & (n2928 | n3911);
  assign n4493 = (n4399 | n3904) & (n4401 | n3905);
  assign n4494 = n2949 | n3907;
  assign n4495 = n4494 & (n3894 | (n4482 & n4481));
  assign n4496 = n4495 & (n3740 | (n4484 & n4483));
  assign n4497 = ~n2981 & (n3895 | (n4487 & n4488));
  assign n4498 = n4497 & (n3743 | (n4490 & n4489));
  assign n4499 = n2628 & (n3737 | (n4492 & n4491));
  assign n4500 = n2921 | n3913;
  assign n4501 = n2624 | ~n3184;
  assign n4502 = n2977 | n3913;
  assign n4503 = n2893 | n3913;
  assign n4504 = n2949 | n3913;
  assign n4505 = (n2924 | n3870) & (n2980 | n3877);
  assign n4506 = (n2896 | n3884) & (n2952 | n3891);
  assign n4507 = (n3036 | n3677) & (n2867 | ~n3898);
  assign n4508 = n3823 & (n813 | n3967);
  assign n4509 = n2647 & (n3825 | n3967);
  assign n4510 = n2646 & (n3822 | n3967);
  assign n4511 = (n2750 | ~n4004) & (n3912 | ~n4003);
  assign n4512 = (n2681 | n3935) & (n2682 | n1556);
  assign n4513 = (n2679 | n3935) & (n2680 | n1556);
  assign n4514 = (n2677 | n3935) & (n2678 | n1556);
  assign n4515 = n2699 | ~n3184;
  assign n4516 = n4515 & (n2675 | n3933);
  assign n4517 = (n2658 | n3935) & (n2659 | n1556);
  assign n4518 = (n2656 | n3935) & (n2657 | n1556);
  assign n4519 = (n2654 | n3935) & (n2655 | n1556);
  assign n4520 = n4515 & (n2652 | n3933);
  assign n4521 = (n2687 | n3935) & (n2688 | n1556);
  assign n4522 = (n2685 | n3935) & (n2686 | n1556);
  assign n4523 = (n2683 | n3935) & (n2684 | n1556);
  assign n4524 = n4515 & (n2676 | n3933);
  assign n4525 = (n2664 | n3935) & (n2665 | n1556);
  assign n4526 = (n2662 | n3935) & (n2663 | n1556);
  assign n4527 = (n2660 | n3935) & (n2661 | n1556);
  assign n4528 = n2653 | n3933;
  assign n4529 = (n2727 | n3870) & (n2749 | n3877);
  assign n4530 = (n2716 | n3884) & (n2738 | n3891);
  assign n4531 = n2700 | n2704;
  assign n4532 = n4531 & (n3327 | (n4530 & n4529));
  assign n4533 = (n4404 | n3940) & (n2459 | n3941);
  assign n4534 = (n2681 | n3942) & (n2682 | n3943);
  assign n4535 = (n4405 | n3940) & (n2482 | n3941);
  assign n4536 = (n2687 | n3942) & (n2688 | n3943);
  assign n4537 = (n2545 | n3940) & (n2721 | n3941);
  assign n4538 = (n2679 | n3942) & (n2680 | n3943);
  assign n4539 = (n4408 | n3940) & (n2718 | n3941);
  assign n4540 = (n2677 | n3942) & (n2678 | n3943);
  assign n4541 = (n2571 | n3940) & (n2710 | n3941);
  assign n4542 = (n2685 | n3942) & (n2686 | n3943);
  assign n4543 = (n4411 | n3940) & (n2706 | n3941);
  assign n4544 = (n2683 | n3942) & (n2684 | n3943);
  assign n4545 = (n2675 | n3938) & (n2676 | n3939);
  assign n4546 = ~n2692 & (n3894 | (n4533 & n4534));
  assign n4547 = n4545 & n4546 & (Pi24 | n2691);
  assign n4548 = ~n2693 & (n3895 | (n4539 & n4540));
  assign n4549 = n4548 & (n3743 | (n4542 & n4541));
  assign n4550 = n2639 & (n3737 | (n4544 & n4543));
  assign n4551 = (n4414 | n3940) & (n2499 | n3941);
  assign n4552 = (n2658 | n3942) & (n2659 | n3943);
  assign n4553 = (n4415 | n3940) & (n2516 | n3941);
  assign n4554 = (n2664 | n3942) & (n2665 | n3943);
  assign n4555 = (n2595 | n3940) & (n2743 | n3941);
  assign n4556 = (n2656 | n3942) & (n2657 | n3943);
  assign n4557 = (n4418 | n3940) & (n2740 | n3941);
  assign n4558 = (n2654 | n3942) & (n2655 | n3943);
  assign n4559 = (n2619 | n3940) & (n2732 | n3941);
  assign n4560 = (n2662 | n3942) & (n2663 | n3943);
  assign n4561 = (n4421 | n3940) & (n2729 | n3941);
  assign n4562 = (n2660 | n3942) & (n2661 | n3943);
  assign n4563 = (n2652 | n3938) & (n2653 | n3939);
  assign n4564 = ~n2669 & (n3894 | (n4551 & n4552));
  assign n4565 = ~n2670 & (n3895 | (n4557 & n4558));
  assign n4566 = (n2750 | ~n4009) & (n3912 | ~n4008);
  assign n4567 = (n2681 | n3947) & (n2682 | n1615);
  assign n4568 = (n2679 | n3947) & (n2680 | n1615);
  assign n4569 = (n2677 | n3947) & (n2678 | n1615);
  assign n4570 = n2754 | ~n3184;
  assign n4571 = n4570 & (n2675 | n3945);
  assign n4572 = (n2658 | n3947) & (n2659 | n1615);
  assign n4573 = (n2656 | n3947) & (n2657 | n1615);
  assign n4574 = (n2654 | n3947) & (n2655 | n1615);
  assign n4575 = n4570 & (n2652 | n3945);
  assign n4576 = (n2687 | n3947) & (n2688 | n1615);
  assign n4577 = (n2685 | n3947) & (n2686 | n1615);
  assign n4578 = (n2683 | n3947) & (n2684 | n1615);
  assign n4579 = n4570 & (n2676 | n3945);
  assign n4580 = (n2664 | n3947) & (n2665 | n1615);
  assign n4581 = (n2662 | n3947) & (n2663 | n1615);
  assign n4582 = (n2660 | n3947) & (n2661 | n1615);
  assign n4583 = n2653 | n3945;
  assign n4584 = (n2774 | n3870) & (n2792 | n3877);
  assign n4585 = (n2765 | n3884) & (n2783 | n3891);
  assign n4586 = n2704 | n2755;
  assign n4587 = n4586 & (n3327 | (n4585 & n4584));
  assign n4588 = (n2636 | n3677) & (n2621 | ~n3898);
  assign n4589 = ~n3176 & (n2066 | n2697) & ~n3177;
  assign n4590 = (~Pi26 | n3971) & (~Ni40 | n3970);
  assign n4591 = (~Pi27 | n3971) & (~Ni41 | n3970);
  assign n4592 = (n3345 | n2372) & (n3352 | n1314);
  assign n4593 = (n3365 | n2372) & (n3372 | n1314);
  assign n4594 = (n3397 | n2372) & (n3403 | n1314);
  assign n4595 = (n3410 | n2372) & (n3417 | n1314);
  assign n4596 = (n3425 | n2372) & (n3430 | n1314);
  assign n4597 = (n3437 | n2372) & (n3444 | n1314);
  assign n4598 = n3476 | n1929;
  assign n4599 = n4598 & (n3894 | (n4592 & n3472));
  assign n4600 = ~n3479 & (n3895 | (n3472 & n4595));
  assign n4601 = ~n3773 & (n3737 | (n3472 & n4597));
  assign n4602 = (n3379 | n2372) & (n3381 | n1314);
  assign n4603 = (n3386 | n2372) & (n3388 | n1314);
  assign n4604 = (n3450 | n2372) & (n3452 | n1314);
  assign n4605 = (n3454 | n2372) & (n3456 | n1314);
  assign n4606 = (n3461 | n2372) & (n3463 | n1314);
  assign n4607 = (n3465 | n2372) & (n3467 | n1314);
  assign n4608 = n3473 | n1929;
  assign n4609 = (n3420 | n3870) & (n3459 | n3877);
  assign n4610 = (n3447 | n3884) & (n3470 | n3891);
  assign n4611 = (n3358 | n3870) & (n3384 | n3877);
  assign n4612 = (n3377 | n3884) & (n3391 | n3891);
  assign n4613 = (n3484 | n2372) & (n3485 | n1314);
  assign n4614 = (n3489 | n2372) & (n3490 | n1314);
  assign n4615 = (n3504 | n2372) & (n3505 | n1314);
  assign n4616 = (n3506 | n2372) & (n3507 | n1314);
  assign n4617 = (n3511 | n2372) & (n3512 | n1314);
  assign n4618 = (n3513 | n2372) & (n3514 | n1314);
  assign n4619 = n3535 | n1929;
  assign n4620 = n4619 & (n3894 | (n4613 & n3472));
  assign n4621 = ~n3538 & (n3895 | (n3472 & n4616));
  assign n4622 = ~n3773 & (n3737 | (n3472 & n4618));
  assign n4623 = (n3494 | n2372) & (n3495 | n1314);
  assign n4624 = (n3499 | n2372) & (n3500 | n1314);
  assign n4625 = (n3518 | n2372) & (n3519 | n1314);
  assign n4626 = (n3520 | n2372) & (n3521 | n1314);
  assign n4627 = (n3525 | n2372) & (n3526 | n1314);
  assign n4628 = (n3527 | n2372) & (n3528 | n1314);
  assign n4629 = n3532 | n1929;
  assign n4630 = (n3510 | n3870) & (n3524 | n3877);
  assign n4631 = (n3517 | n3884) & (n3531 | n3891);
  assign n4632 = (n3488 | n3870) & (n3498 | n3877);
  assign n4633 = (n3493 | n3884) & (n3503 | n3891);
  assign n4634 = (n3300 | n3618) & (n3551 | n1929);
  assign n4635 = (n3302 | n3618) & (n3553 | n1929);
  assign n4636 = (n3316 | n3618) & (n3575 | n1929);
  assign n4637 = (n3318 | n3618) & (n3579 | n1929);
  assign n4638 = (n3319 | n3618) & (n3586 | n1929);
  assign n4639 = (n3321 | n3618) & (n3590 | n1929);
  assign n4640 = ~n3654 & (n3895 | (n3621 & n4637));
  assign n4641 = ~n3655 & (n3737 | (n3621 & n4639));
  assign n4642 = (n3310 | n3618) & (n3588 | n1929);
  assign n4643 = (n3312 | n3618) & (n3592 | n1929);
  assign n4644 = (n3650 | n2272) & (n3651 | n3895);
  assign n4645 = (n3645 | n3978) & (n3649 | n3979);
  assign n4646 = (n3234 | n3618) & (n3567 | n1929);
  assign n4647 = (n3240 | n3618) & (n3569 | n1929);
  assign n4648 = (n3268 | n3618) & (n3597 | n1929);
  assign n4649 = (n3273 | n3618) & (n3601 | n1929);
  assign n4650 = (n3277 | n3618) & (n3608 | n1929);
  assign n4651 = (n3282 | n3618) & (n3612 | n1929);
  assign n4652 = ~n3638 & (n3895 | (n3621 & n4649));
  assign n4653 = ~n3639 & (n3737 | (n3621 & n4651));
  assign n4654 = (n3256 | n3618) & (n3610 | n1929);
  assign n4655 = (n3261 | n3618) & (n3614 | n1929);
  assign n4656 = (n3633 | n2272) & (n3634 | n3895);
  assign n4657 = (n3628 | n3978) & (n3632 | n3979);
  assign n4658 = (n3584 | n3870) & (n3606 | n3877);
  assign n4659 = (n3595 | n3884) & (n3617 | n3891);
  assign n4660 = (n3548 | n3870) & (n3565 | n3877);
  assign n4661 = (n3557 | n3884) & (n3573 | n3891);
  assign n4662 = n3912 | n1543 | n4744 | n4745;
  assign n4663 = n2074 | n3669 | n795 | ~Ni10;
  assign n4664 = n3768 | n3669 | n3767;
  assign n4665 = Ni31 & (~Ni30 | ~Ni5 | Ni4);
  assign n4666 = (~Pi15 & n1312) | (n1305 & (Pi15 | n1312));
  assign n4667 = ~Pi17 & (n1296 | n1298 | ~n4089);
  assign n4668 = ~n4667 & (~Pi17 | (n4090 & n4091));
  assign n4669 = (~n3327 & n4668) | (n4666 & (n3327 | n4668));
  assign n4670 = n4110 & ~n3892 & n4109;
  assign n4671 = ~n2074 & (n4670 | (n3892 & n4668));
  assign n4672 = ~Ni7 & (n4671 | (n2074 & n4669));
  assign n4673 = ~n3707 & (n4672 | (Ni7 & n4669));
  assign n4674 = Ni14 & n4258 & n3802;
  assign n4675 = n4179 & ~Ni14 & n4178;
  assign n4676 = Ni14 & n4186 & n4185;
  assign n4677 = n1943 | ~n4148 | n1941 | n1942 | ~n1362 | ~n1536 | n1939 | n1940;
  assign n4678 = n1935 | ~n4162 | n1933 | n1934 | ~n1362 | ~n1498 | n1931 | n1932;
  assign n4679 = n1787 | n3906;
  assign n4680 = n4679 & n4221 & n4220 & n4218 & ~Pi15 & n4215;
  assign n4681 = n1857 | n3906;
  assign n4682 = Pi15 & n4239 & n4240 & n4237 & n4234 & n4681;
  assign n4683 = Pi17 & (~n4133 | ~n4134);
  assign n4684 = n4165 & n4164 & ~Pi17 & n1362;
  assign n4685 = Pi17 & n4167 & n4168 & n1362;
  assign n4686 = n4248 & Ni10 & (Ni11 | n1865);
  assign n4687 = n4170 & ~Pi17 & n4169;
  assign n4688 = n2383 | n3737;
  assign n4689 = n4688 & n4303 & n4302 & n4301 & ~Pi15 & n2371;
  assign n4690 = n18 | ~Ni34;
  assign n4691 = n1539 | Ni34 | n18;
  assign n4692 = n4317 & ~Pi17 & n4316;
  assign n4693 = Pi17 & n4319 & n4318;
  assign n4694 = Pi20 & (~n4339 | ~n4341);
  assign n4695 = ~n4694 & (Pi20 | (n4329 & n4331));
  assign n4696 = Pi20 & (~n4362 | ~n4364);
  assign n4697 = ~n4696 & (Pi20 | (n4352 & n4354));
  assign n4698 = n4695 & ~Pi15 & n4342;
  assign n4699 = Pi15 & n4365 & n4697;
  assign n4700 = n4692 | n4693 | n3327 | Ni10;
  assign n4701 = ~Pi17 & (~n4373 | ~n4374);
  assign n4702 = n2393 & n4377 & n2390;
  assign n4703 = ~n2393 & (n3808 | (~Pi23 & n2392));
  assign n4704 = n2393 & n4378 & n2400;
  assign n4705 = ~n2393 & (n3809 | (~Pi24 & n2401));
  assign n4706 = ~n2393 & (Ni33 | n886) & n2401;
  assign n4707 = ~Ni44 & ~Ni39 & (~n3733 | Ni42);
  assign n4708 = ~n4707 & (~Ni44 | ~n923 | ~Ni39);
  assign n4709 = Pi21 | n3818;
  assign n4710 = (~Pi26 & ~n2648) | (~n2644 & (Pi26 | ~n2648));
  assign n4711 = ~Pi21 & (~n2623 | (~Pi26 & Ni32));
  assign n4712 = (Pi26 & ~n2648) | (~n2644 & (~Pi26 | ~n2648));
  assign n4713 = n4442 & ~Ni14 & n4441;
  assign n4714 = n3059 | ~n4413 | n3057 | n3058 | ~n2423 | ~n2691 | n3055 | n3056;
  assign n4715 = n3052 | ~n4423 | n3050 | n3051 | ~n2423 | ~n2668 | n3048 | n3049;
  assign n4716 = n2921 | n3906;
  assign n4717 = n4716 & n4480 & n4479 & n4477 & ~Pi15 & n4474;
  assign n4718 = n2977 | n3906;
  assign n4719 = Pi15 & n4498 & n4499 & n4496 & n4493 & n4718;
  assign n4720 = Pi17 & (~n4402 | ~n4403);
  assign n4721 = n4426 & n4425 & ~Pi17 & n2423;
  assign n4722 = Pi17 & n4428 & n4429 & n2423;
  assign n4723 = n4507 & Ni10 & (Ni11 | n2985);
  assign n4724 = n2703 | n2701 | n2702;
  assign n4725 = n4433 & ~Pi17 & n4432;
  assign n4726 = ~Pi20 & n3968 & (n3183 | ~Ni39);
  assign n4727 = n3968 & Pi20 & (Ni39 | n3183);
  assign n4728 = ~n2393 | ~Ni40;
  assign n4729 = (n3830 & (~n2393 | ~n4012)) | (n2393 & ~n4012);
  assign n4730 = ~n2393 | ~Ni41;
  assign n4731 = (n3833 & (~n2393 | ~n4016)) | (n2393 & ~n4016);
  assign n4732 = ~Pi21 & (n797 | (~n1539 & n3186));
  assign n4733 = Pi20 & (n3652 | n3653 | ~n4644);
  assign n4734 = ~n4733 & (Pi20 | (n4640 & n4641));
  assign n4735 = Pi20 & (n3636 | n3637 | ~n4656);
  assign n4736 = ~n4735 & (Pi20 | (n4652 & n4653));
  assign n4737 = n4734 & ~Pi15 & n4645;
  assign n4738 = Pi15 & n4657 & n4736;
  assign n4739 = n4659 & ~Pi17 & n4658;
  assign n4740 = ~Ni10 & (n4737 | n4738);
  assign n4741 = n4601 & n4600 & n4599 & ~n3478 & ~Pi15 & ~n3477;
  assign n4742 = n4610 & ~Pi17 & n4609;
  assign n4743 = Pi17 & n4612 & n4611;
  assign n4744 = ~Ni10 & (n4741 | (Pi15 & n4023));
  assign n4745 = Ni10 & (n4742 | n4743);
  assign n4746 = n4622 & n4621 & n4620 & ~n3537 & ~Pi15 & ~n3536;
  assign n4747 = n4631 & ~Pi17 & n4630;
  assign n4748 = Pi17 & n4633 & n4632;
  assign n4749 = ~Ni10 & (n4746 | (Pi15 & n4028));
  assign n4750 = n4775 | ~Ni14 | ~Ni12;
  assign n4751 = ~Ni4 & (~Ni6 | ~Ni5 | ~n3700);
  assign n4752 = ~Ni5 | ~Ni31 | ~Ni6;
  assign n4753 = n4752 & Ni4 & (n2418 | n3980);
  assign n4754 = Ni3 & (n4753 | (~Ni4 & ~n4752));
  assign n4755 = ~Ni2 & (n4754 | (~Ni3 & n4034));
  assign n4756 = Ni6 & (Ni2 | (~Ni31 & Ni3));
  assign n4757 = Ni12 & (n3707 | (~n3723 & n3727));
  assign n4758 = Pi20 & (n806 | n3745 | n3755);
  assign n4759 = Ni42 & (~Ni44 | n3732) & ~Ni39;
  assign n4760 = Pi27 | n3985;
  assign n4761 = ~Pi27 | Pi26 | n3985;
  assign n4762 = Pi24 | n3986;
  assign n4763 = ~Pi24 | Pi23 | n3986;
  assign n4764 = ~Ni4 & (n2416 | n3973);
  assign n4765 = Ni4 & (Ni33 | n3980);
  assign n4766 = Ni33 & ~n1352;
  assign n4767 = ~Ni33 & ~n1352;
  assign n4768 = n698 | n2433;
  assign n4769 = ~n674 | Ni41;
  assign n4770 = ~n675 | Ni41;
  assign n4771 = ~Ni33 | n3201;
  assign n4772 = n1540 & n1463;
  assign n4773 = n1546 | n1547 | n1548 | ~n4291;
  assign n4774 = n3984 | n4726 | n4727;
  assign n4775 = n3669 & Pi27;
  assign n1085 = P__cmxcl_0;
  always @ (posedge clk) begin
    Ni48 <= n931_1;
    Ni47 <= n936;
    Ni46 <= n941_1;
    Ni45 <= n946_1;
    Ni44 <= n951_1;
    Ni43 <= n956_1;
    Ni42 <= n961_1;
    Ni41 <= n966_1;
    Ni40 <= n971;
    Ni39 <= n976_1;
    Ni38 <= n981_1;
    Ni37 <= n986;
    Ni36 <= n991_1;
    Ni35 <= n996_1;
    Ni34 <= n1001;
    Ni33 <= n1006_1;
    Ni32 <= n1011_1;
    Ni31 <= n1016_1;
    Ni30 <= n1021;
    n18 <= n1026_1;
    Ni14 <= n1031_1;
    Ni13 <= n1036;
    Ni12 <= n1041_1;
    Ni11 <= n1046_1;
    Ni10 <= n1051;
    Ni9 <= n1056_1;
    Ni8 <= n1061;
    Ni7 <= n1066_1;
    Ni6 <= n1071_1;
    Ni5 <= n1076;
    Ni4 <= n1081;
    Ni3 <= n1085;
    Ni2 <= n1090_1;
  end
endmodule


