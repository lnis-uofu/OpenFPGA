// Benchmark "TOP" written by ABC on Tue Mar  5 09:55:28 2019

module bigkey ( clock, 
    Pstart_0_, Pkey_255_, Pkey_254_, Pkey_253_, Pkey_252_, Pkey_251_,
    Pkey_250_, Pkey_249_, Pkey_248_, Pkey_247_, Pkey_246_, Pkey_245_,
    Pkey_244_, Pkey_243_, Pkey_242_, Pkey_241_, Pkey_240_, Pkey_239_,
    Pkey_238_, Pkey_237_, Pkey_236_, Pkey_235_, Pkey_234_, Pkey_233_,
    Pkey_232_, Pkey_231_, Pkey_230_, Pkey_229_, Pkey_228_, Pkey_227_,
    Pkey_226_, Pkey_225_, Pkey_224_, Pkey_223_, Pkey_222_, Pkey_221_,
    Pkey_220_, Pkey_219_, Pkey_218_, Pkey_217_, Pkey_216_, Pkey_215_,
    Pkey_214_, Pkey_213_, Pkey_212_, Pkey_211_, Pkey_210_, Pkey_209_,
    Pkey_208_, Pkey_207_, Pkey_206_, Pkey_205_, Pkey_204_, Pkey_203_,
    Pkey_202_, Pkey_201_, Pkey_200_, Pkey_199_, Pkey_198_, Pkey_197_,
    Pkey_196_, Pkey_195_, Pkey_194_, Pkey_193_, Pkey_192_, Pkey_191_,
    Pkey_190_, Pkey_189_, Pkey_188_, Pkey_187_, Pkey_186_, Pkey_185_,
    Pkey_184_, Pkey_183_, Pkey_182_, Pkey_181_, Pkey_180_, Pkey_179_,
    Pkey_178_, Pkey_177_, Pkey_176_, Pkey_175_, Pkey_174_, Pkey_173_,
    Pkey_172_, Pkey_171_, Pkey_170_, Pkey_169_, Pkey_168_, Pkey_167_,
    Pkey_166_, Pkey_165_, Pkey_164_, Pkey_163_, Pkey_162_, Pkey_161_,
    Pkey_160_, Pkey_159_, Pkey_158_, Pkey_157_, Pkey_156_, Pkey_155_,
    Pkey_154_, Pkey_153_, Pkey_152_, Pkey_151_, Pkey_150_, Pkey_149_,
    Pkey_148_, Pkey_147_, Pkey_146_, Pkey_145_, Pkey_144_, Pkey_143_,
    Pkey_142_, Pkey_141_, Pkey_140_, Pkey_139_, Pkey_138_, Pkey_137_,
    Pkey_136_, Pkey_135_, Pkey_134_, Pkey_133_, Pkey_132_, Pkey_131_,
    Pkey_130_, Pkey_129_, Pkey_128_, Pkey_127_, Pkey_126_, Pkey_125_,
    Pkey_124_, Pkey_123_, Pkey_122_, Pkey_121_, Pkey_120_, Pkey_119_,
    Pkey_118_, Pkey_117_, Pkey_116_, Pkey_115_, Pkey_114_, Pkey_113_,
    Pkey_112_, Pkey_111_, Pkey_110_, Pkey_109_, Pkey_108_, Pkey_107_,
    Pkey_106_, Pkey_105_, Pkey_104_, Pkey_103_, Pkey_102_, Pkey_101_,
    Pkey_100_, Pkey_99_, Pkey_98_, Pkey_97_, Pkey_96_, Pkey_95_, Pkey_94_,
    Pkey_93_, Pkey_92_, Pkey_91_, Pkey_90_, Pkey_89_, Pkey_88_, Pkey_87_,
    Pkey_86_, Pkey_85_, Pkey_84_, Pkey_83_, Pkey_82_, Pkey_81_, Pkey_80_,
    Pkey_79_, Pkey_78_, Pkey_77_, Pkey_76_, Pkey_75_, Pkey_74_, Pkey_73_,
    Pkey_72_, Pkey_71_, Pkey_70_, Pkey_69_, Pkey_68_, Pkey_67_, Pkey_66_,
    Pkey_65_, Pkey_64_, Pkey_63_, Pkey_62_, Pkey_61_, Pkey_60_, Pkey_59_,
    Pkey_58_, Pkey_57_, Pkey_56_, Pkey_55_, Pkey_54_, Pkey_53_, Pkey_52_,
    Pkey_51_, Pkey_50_, Pkey_49_, Pkey_48_, Pkey_47_, Pkey_46_, Pkey_45_,
    Pkey_44_, Pkey_43_, Pkey_42_, Pkey_41_, Pkey_40_, Pkey_39_, Pkey_38_,
    Pkey_37_, Pkey_36_, Pkey_35_, Pkey_34_, Pkey_33_, Pkey_32_, Pkey_31_,
    Pkey_30_, Pkey_29_, Pkey_28_, Pkey_27_, Pkey_26_, Pkey_25_, Pkey_24_,
    Pkey_23_, Pkey_22_, Pkey_21_, Pkey_20_, Pkey_19_, Pkey_18_, Pkey_17_,
    Pkey_16_, Pkey_15_, Pkey_14_, Pkey_13_, Pkey_12_, Pkey_11_, Pkey_10_,
    Pkey_9_, Pkey_8_, Pkey_7_, Pkey_6_, Pkey_5_, Pkey_4_, Pkey_3_, Pkey_2_,
    Pkey_1_, Pkey_0_, Pencrypt_0_, Pcount_3_, Pcount_2_, Pcount_1_,
    Pcount_0_, 
    Pnew_count_3_, Pnew_count_2_, Pnew_count_1_, Pnew_count_0_,
    Pdata_ready_0_, PKSi_191_, PKSi_190_, PKSi_189_, PKSi_188_, PKSi_187_,
    PKSi_186_, PKSi_185_, PKSi_184_, PKSi_183_, PKSi_182_, PKSi_181_,
    PKSi_180_, PKSi_179_, PKSi_178_, PKSi_177_, PKSi_176_, PKSi_175_,
    PKSi_174_, PKSi_173_, PKSi_172_, PKSi_171_, PKSi_170_, PKSi_169_,
    PKSi_168_, PKSi_167_, PKSi_166_, PKSi_165_, PKSi_164_, PKSi_163_,
    PKSi_162_, PKSi_161_, PKSi_160_, PKSi_159_, PKSi_158_, PKSi_157_,
    PKSi_156_, PKSi_155_, PKSi_154_, PKSi_153_, PKSi_152_, PKSi_151_,
    PKSi_150_, PKSi_149_, PKSi_148_, PKSi_147_, PKSi_146_, PKSi_145_,
    PKSi_144_, PKSi_143_, PKSi_142_, PKSi_141_, PKSi_140_, PKSi_139_,
    PKSi_138_, PKSi_137_, PKSi_136_, PKSi_135_, PKSi_134_, PKSi_133_,
    PKSi_132_, PKSi_131_, PKSi_130_, PKSi_129_, PKSi_128_, PKSi_127_,
    PKSi_126_, PKSi_125_, PKSi_124_, PKSi_123_, PKSi_122_, PKSi_121_,
    PKSi_120_, PKSi_119_, PKSi_118_, PKSi_117_, PKSi_116_, PKSi_115_,
    PKSi_114_, PKSi_113_, PKSi_112_, PKSi_111_, PKSi_110_, PKSi_109_,
    PKSi_108_, PKSi_107_, PKSi_106_, PKSi_105_, PKSi_104_, PKSi_103_,
    PKSi_102_, PKSi_101_, PKSi_100_, PKSi_99_, PKSi_98_, PKSi_97_,
    PKSi_96_, PKSi_95_, PKSi_94_, PKSi_93_, PKSi_92_, PKSi_91_, PKSi_90_,
    PKSi_89_, PKSi_88_, PKSi_87_, PKSi_86_, PKSi_85_, PKSi_84_, PKSi_83_,
    PKSi_82_, PKSi_81_, PKSi_80_, PKSi_79_, PKSi_78_, PKSi_77_, PKSi_76_,
    PKSi_75_, PKSi_74_, PKSi_73_, PKSi_72_, PKSi_71_, PKSi_70_, PKSi_69_,
    PKSi_68_, PKSi_67_, PKSi_66_, PKSi_65_, PKSi_64_, PKSi_63_, PKSi_62_,
    PKSi_61_, PKSi_60_, PKSi_59_, PKSi_58_, PKSi_57_, PKSi_56_, PKSi_55_,
    PKSi_54_, PKSi_53_, PKSi_52_, PKSi_51_, PKSi_50_, PKSi_49_, PKSi_48_,
    PKSi_47_, PKSi_46_, PKSi_45_, PKSi_44_, PKSi_43_, PKSi_42_, PKSi_41_,
    PKSi_40_, PKSi_39_, PKSi_38_, PKSi_37_, PKSi_36_, PKSi_35_, PKSi_34_,
    PKSi_33_, PKSi_32_, PKSi_31_, PKSi_30_, PKSi_29_, PKSi_28_, PKSi_27_,
    PKSi_26_, PKSi_25_, PKSi_24_, PKSi_23_, PKSi_22_, PKSi_21_, PKSi_20_,
    PKSi_19_, PKSi_18_, PKSi_17_, PKSi_16_, PKSi_15_, PKSi_14_, PKSi_13_,
    PKSi_12_, PKSi_11_, PKSi_10_, PKSi_9_, PKSi_8_, PKSi_7_, PKSi_6_,
    PKSi_5_, PKSi_4_, PKSi_3_, PKSi_2_, PKSi_1_, PKSi_0_  );
  input  Pstart_0_, Pkey_255_, Pkey_254_, Pkey_253_, Pkey_252_,
    Pkey_251_, Pkey_250_, Pkey_249_, Pkey_248_, Pkey_247_, Pkey_246_,
    Pkey_245_, Pkey_244_, Pkey_243_, Pkey_242_, Pkey_241_, Pkey_240_,
    Pkey_239_, Pkey_238_, Pkey_237_, Pkey_236_, Pkey_235_, Pkey_234_,
    Pkey_233_, Pkey_232_, Pkey_231_, Pkey_230_, Pkey_229_, Pkey_228_,
    Pkey_227_, Pkey_226_, Pkey_225_, Pkey_224_, Pkey_223_, Pkey_222_,
    Pkey_221_, Pkey_220_, Pkey_219_, Pkey_218_, Pkey_217_, Pkey_216_,
    Pkey_215_, Pkey_214_, Pkey_213_, Pkey_212_, Pkey_211_, Pkey_210_,
    Pkey_209_, Pkey_208_, Pkey_207_, Pkey_206_, Pkey_205_, Pkey_204_,
    Pkey_203_, Pkey_202_, Pkey_201_, Pkey_200_, Pkey_199_, Pkey_198_,
    Pkey_197_, Pkey_196_, Pkey_195_, Pkey_194_, Pkey_193_, Pkey_192_,
    Pkey_191_, Pkey_190_, Pkey_189_, Pkey_188_, Pkey_187_, Pkey_186_,
    Pkey_185_, Pkey_184_, Pkey_183_, Pkey_182_, Pkey_181_, Pkey_180_,
    Pkey_179_, Pkey_178_, Pkey_177_, Pkey_176_, Pkey_175_, Pkey_174_,
    Pkey_173_, Pkey_172_, Pkey_171_, Pkey_170_, Pkey_169_, Pkey_168_,
    Pkey_167_, Pkey_166_, Pkey_165_, Pkey_164_, Pkey_163_, Pkey_162_,
    Pkey_161_, Pkey_160_, Pkey_159_, Pkey_158_, Pkey_157_, Pkey_156_,
    Pkey_155_, Pkey_154_, Pkey_153_, Pkey_152_, Pkey_151_, Pkey_150_,
    Pkey_149_, Pkey_148_, Pkey_147_, Pkey_146_, Pkey_145_, Pkey_144_,
    Pkey_143_, Pkey_142_, Pkey_141_, Pkey_140_, Pkey_139_, Pkey_138_,
    Pkey_137_, Pkey_136_, Pkey_135_, Pkey_134_, Pkey_133_, Pkey_132_,
    Pkey_131_, Pkey_130_, Pkey_129_, Pkey_128_, Pkey_127_, Pkey_126_,
    Pkey_125_, Pkey_124_, Pkey_123_, Pkey_122_, Pkey_121_, Pkey_120_,
    Pkey_119_, Pkey_118_, Pkey_117_, Pkey_116_, Pkey_115_, Pkey_114_,
    Pkey_113_, Pkey_112_, Pkey_111_, Pkey_110_, Pkey_109_, Pkey_108_,
    Pkey_107_, Pkey_106_, Pkey_105_, Pkey_104_, Pkey_103_, Pkey_102_,
    Pkey_101_, Pkey_100_, Pkey_99_, Pkey_98_, Pkey_97_, Pkey_96_, Pkey_95_,
    Pkey_94_, Pkey_93_, Pkey_92_, Pkey_91_, Pkey_90_, Pkey_89_, Pkey_88_,
    Pkey_87_, Pkey_86_, Pkey_85_, Pkey_84_, Pkey_83_, Pkey_82_, Pkey_81_,
    Pkey_80_, Pkey_79_, Pkey_78_, Pkey_77_, Pkey_76_, Pkey_75_, Pkey_74_,
    Pkey_73_, Pkey_72_, Pkey_71_, Pkey_70_, Pkey_69_, Pkey_68_, Pkey_67_,
    Pkey_66_, Pkey_65_, Pkey_64_, Pkey_63_, Pkey_62_, Pkey_61_, Pkey_60_,
    Pkey_59_, Pkey_58_, Pkey_57_, Pkey_56_, Pkey_55_, Pkey_54_, Pkey_53_,
    Pkey_52_, Pkey_51_, Pkey_50_, Pkey_49_, Pkey_48_, Pkey_47_, Pkey_46_,
    Pkey_45_, Pkey_44_, Pkey_43_, Pkey_42_, Pkey_41_, Pkey_40_, Pkey_39_,
    Pkey_38_, Pkey_37_, Pkey_36_, Pkey_35_, Pkey_34_, Pkey_33_, Pkey_32_,
    Pkey_31_, Pkey_30_, Pkey_29_, Pkey_28_, Pkey_27_, Pkey_26_, Pkey_25_,
    Pkey_24_, Pkey_23_, Pkey_22_, Pkey_21_, Pkey_20_, Pkey_19_, Pkey_18_,
    Pkey_17_, Pkey_16_, Pkey_15_, Pkey_14_, Pkey_13_, Pkey_12_, Pkey_11_,
    Pkey_10_, Pkey_9_, Pkey_8_, Pkey_7_, Pkey_6_, Pkey_5_, Pkey_4_,
    Pkey_3_, Pkey_2_, Pkey_1_, Pkey_0_, Pencrypt_0_, Pcount_3_, Pcount_2_,
    Pcount_1_, Pcount_0_, clock;
  output Pnew_count_3_, Pnew_count_2_, Pnew_count_1_, Pnew_count_0_,
    Pdata_ready_0_, PKSi_191_, PKSi_190_, PKSi_189_, PKSi_188_, PKSi_187_,
    PKSi_186_, PKSi_185_, PKSi_184_, PKSi_183_, PKSi_182_, PKSi_181_,
    PKSi_180_, PKSi_179_, PKSi_178_, PKSi_177_, PKSi_176_, PKSi_175_,
    PKSi_174_, PKSi_173_, PKSi_172_, PKSi_171_, PKSi_170_, PKSi_169_,
    PKSi_168_, PKSi_167_, PKSi_166_, PKSi_165_, PKSi_164_, PKSi_163_,
    PKSi_162_, PKSi_161_, PKSi_160_, PKSi_159_, PKSi_158_, PKSi_157_,
    PKSi_156_, PKSi_155_, PKSi_154_, PKSi_153_, PKSi_152_, PKSi_151_,
    PKSi_150_, PKSi_149_, PKSi_148_, PKSi_147_, PKSi_146_, PKSi_145_,
    PKSi_144_, PKSi_143_, PKSi_142_, PKSi_141_, PKSi_140_, PKSi_139_,
    PKSi_138_, PKSi_137_, PKSi_136_, PKSi_135_, PKSi_134_, PKSi_133_,
    PKSi_132_, PKSi_131_, PKSi_130_, PKSi_129_, PKSi_128_, PKSi_127_,
    PKSi_126_, PKSi_125_, PKSi_124_, PKSi_123_, PKSi_122_, PKSi_121_,
    PKSi_120_, PKSi_119_, PKSi_118_, PKSi_117_, PKSi_116_, PKSi_115_,
    PKSi_114_, PKSi_113_, PKSi_112_, PKSi_111_, PKSi_110_, PKSi_109_,
    PKSi_108_, PKSi_107_, PKSi_106_, PKSi_105_, PKSi_104_, PKSi_103_,
    PKSi_102_, PKSi_101_, PKSi_100_, PKSi_99_, PKSi_98_, PKSi_97_,
    PKSi_96_, PKSi_95_, PKSi_94_, PKSi_93_, PKSi_92_, PKSi_91_, PKSi_90_,
    PKSi_89_, PKSi_88_, PKSi_87_, PKSi_86_, PKSi_85_, PKSi_84_, PKSi_83_,
    PKSi_82_, PKSi_81_, PKSi_80_, PKSi_79_, PKSi_78_, PKSi_77_, PKSi_76_,
    PKSi_75_, PKSi_74_, PKSi_73_, PKSi_72_, PKSi_71_, PKSi_70_, PKSi_69_,
    PKSi_68_, PKSi_67_, PKSi_66_, PKSi_65_, PKSi_64_, PKSi_63_, PKSi_62_,
    PKSi_61_, PKSi_60_, PKSi_59_, PKSi_58_, PKSi_57_, PKSi_56_, PKSi_55_,
    PKSi_54_, PKSi_53_, PKSi_52_, PKSi_51_, PKSi_50_, PKSi_49_, PKSi_48_,
    PKSi_47_, PKSi_46_, PKSi_45_, PKSi_44_, PKSi_43_, PKSi_42_, PKSi_41_,
    PKSi_40_, PKSi_39_, PKSi_38_, PKSi_37_, PKSi_36_, PKSi_35_, PKSi_34_,
    PKSi_33_, PKSi_32_, PKSi_31_, PKSi_30_, PKSi_29_, PKSi_28_, PKSi_27_,
    PKSi_26_, PKSi_25_, PKSi_24_, PKSi_23_, PKSi_22_, PKSi_21_, PKSi_20_,
    PKSi_19_, PKSi_18_, PKSi_17_, PKSi_16_, PKSi_15_, PKSi_14_, PKSi_13_,
    PKSi_12_, PKSi_11_, PKSi_10_, PKSi_9_, PKSi_8_, PKSi_7_, PKSi_6_,
    PKSi_5_, PKSi_4_, PKSi_3_, PKSi_2_, PKSi_1_, PKSi_0_;
  reg PKSi_79_, PKSi_92_, \[333] , N_N2737, PKSi_75_, PKSi_84_, N_N2741,
    PKSi_82_, PKSi_93_, PKSi_85_, N_N2746, PKSi_73_, N_N2749, PKSi_80_,
    PKSi_72_, PKSi_94_, PKSi_86_, PKSi_74_, PKSi_83_, N_N2757, PKSi_89_,
    PKSi_91_, PKSi_81_, PKSi_77_, PKSi_87_, PKSi_78_, PKSi_95_, PKSi_76_,
    PKSi_55_, PKSi_68_, PKSi_64_, N_N2770, PKSi_51_, PKSi_60_, N_N2774,
    PKSi_58_, PKSi_69_, PKSi_61_, N_N2779, PKSi_49_, PKSi_66_, PKSi_56_,
    PKSi_48_, PKSi_70_, PKSi_62_, PKSi_50_, PKSi_59_, N_N2789, PKSi_65_,
    PKSi_67_, PKSi_57_, PKSi_53_, PKSi_63_, PKSi_54_, PKSi_71_, PKSi_52_,
    PKSi_31_, PKSi_44_, PKSi_40_, N_N2802, PKSi_27_, PKSi_36_, N_N2806,
    PKSi_34_, PKSi_45_, PKSi_37_, N_N2811, PKSi_25_, PKSi_42_, PKSi_32_,
    PKSi_24_, PKSi_46_, PKSi_38_, PKSi_26_, PKSi_35_, N_N2821, PKSi_41_,
    PKSi_43_, PKSi_33_, PKSi_29_, PKSi_39_, PKSi_30_, PKSi_47_, PKSi_28_,
    PKSi_7_, PKSi_20_, PKSi_16_, N_N2834, PKSi_3_, PKSi_12_, N_N2838,
    PKSi_10_, PKSi_21_, PKSi_13_, N_N2843, PKSi_1_, PKSi_18_, PKSi_8_,
    PKSi_0_, PKSi_22_, PKSi_14_, PKSi_2_, PKSi_11_, N_N2853, PKSi_17_,
    PKSi_19_, PKSi_9_, PKSi_5_, PKSi_15_, PKSi_6_, PKSi_23_, PKSi_4_,
    PKSi_183_, PKSi_173_, N_N2865, PKSi_185_, PKSi_169_, PKSi_176_,
    PKSi_188_, \[253] , PKSi_179_, PKSi_172_, PKSi_186_, PKSi_177_,
    PKSi_180_, N_N2877, N_N2879, N_N2881, PKSi_175_, PKSi_182_, N_N2885,
    PKSi_171_, PKSi_189_, N_N2889, PKSi_184_, PKSi_178_, \[234] ,
    PKSi_170_, PKSi_174_, PKSi_190_, PKSi_159_, PKSi_149_, N_N2899,
    PKSi_161_, PKSi_145_, PKSi_152_, PKSi_164_, PKSi_157_, PKSi_155_,
    PKSi_148_, PKSi_162_, N_N2909, PKSi_156_, PKSi_153_, PKSi_163_,
    PKSi_144_, PKSi_151_, PKSi_158_, N_N2917, PKSi_147_, PKSi_165_,
    N_N2921, PKSi_160_, PKSi_154_, PKSi_167_, PKSi_146_, PKSi_150_,
    PKSi_166_, PKSi_135_, PKSi_125_, N_N2931, PKSi_137_, PKSi_121_,
    PKSi_128_, PKSi_140_, PKSi_133_, PKSi_131_, PKSi_124_, PKSi_138_,
    PKSi_129_, PKSi_132_, N_N2943, N_N2945, PKSi_120_, PKSi_127_,
    PKSi_134_, N_N2950, PKSi_123_, PKSi_141_, N_N2954, PKSi_136_,
    PKSi_130_, \[282] , PKSi_122_, PKSi_126_, PKSi_142_, PKSi_111_,
    PKSi_101_, N_N2964, PKSi_113_, PKSi_97_, PKSi_104_, PKSi_116_,
    PKSi_109_, PKSi_107_, PKSi_100_, PKSi_114_, PKSi_105_, PKSi_108_,
    N_N2976, PKSi_115_, PKSi_96_, PKSi_103_, PKSi_110_, N_N2982, PKSi_99_,
    PKSi_117_, N_N2986, PKSi_112_, PKSi_106_, PKSi_119_, PKSi_98_,
    PKSi_102_, PKSi_118_;
  wire n1137, n1138, n1139_1, n1140, n1141, n1142, n1143_1, n1144, n1145,
    n1146, n1148, n1150, n1152, n1154, n1156, n1158, n1160, n1162, n1164,
    n1166, n1168, n1170, n1172_1, n1174, n1176_1, n1178, n1180_1, n1182,
    n1184, n1186, n1188, n1190, n1192, n1194, n1196, n1198, n1200, n1202_1,
    n1204, n1206_1, n1208, n1210_1, n1212, n1214_1, n1216, n1218_1, n1220,
    n1222_1, n1224, n1226_1, n1228, n1230_1, n1232, n1234_1, n1236, n1238,
    n1240, n1242, n1244, n1246, n1248, n1250, n1252, n1254, n1256, n1258,
    n1260, n1262, n1264, n1266, n1268, n1270, n1272, n1274, n1276, n1278,
    n1280, n1282, n1284, n1286, n1288_1, n1290, n1292, n1294, n1296, n1298,
    n1300, n1302, n1304, n1306, n1308, n1310, n1312, n1314, n1316, n1318,
    n1320, n1322, n1324, n1326, n1328, n1330, n1332, n1334, n1336, n1338,
    n1340, n1342, n1344, n1346, n1348, n1350, n1352, n1354, n1356, n1358,
    n1360, n1362, n1364, n1366, n1368, n1370, n1372, n1374, n1376, n1378,
    n1380, n1382, n1384, n1386, n1388, n1390, n1392, n1394, n1396, n1398,
    n1400, n1402, n1404, n1406, n1408, n1410, n1412, n1414, n1416, n1418,
    n1420, n1422, n1424, n1426, n1428, n1430, n1432, n1434, n1436, n1438,
    n1440, n1442, n1444, n1446, n1448, n1450, n1452, n1454, n1456, n1458,
    n1460, n1462, n1464, n1466, n1468, n1470, n1472, n1474, n1476, n1478,
    n1480, n1482, n1484, n1486, n1488, n1490, n1492, n1494, n1496, n1498,
    n1500, n1502, n1504, n1506, n1508, n1510, n1512, n1514, n1516, n1518,
    n1520, n1522, n1524, n1526, n1528, n1530, n1532, n1534, n1536, n1538,
    n1540, n1542, n1544, n1546, n1548, n1550, n1552, n1554, n1556, n1558,
    n1560, n1562, n1564, n1566, n1568, n1570, n1572, n1574, n1576, n1578,
    n1580, n1582, n1584, n1586, n1588, n1590, n1592, n1594, n1595, n1596,
    n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
    n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
    n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
    n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
    n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
    n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
    n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
    n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
    n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
    n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
    n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
    n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
    n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
    n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
    n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745_1, n1746,
    n1747, n1748, n1749_1, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
    n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
    n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
    n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
    n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
    n1797, n1798, n1799_1, n1800, n1801, n1802, n1803_1, n1804, n1805,
    n1806, n1807_1, n1808, n1809, n1810, n1811_1, n1812, n1813, n1814,
    n1815_1, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
    n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833_1, n1834,
    n1835, n1836, n1837_1, n1838, n1839, n1840, n1841_1, n1842, n1843,
    n1844, n1845_1, n1846, n1847, n1848, n1849_1, n1850, n1851, n1852,
    n1853_1, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
    n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
    n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
    n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
    n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
    n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
    n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
    n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
    n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
    n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
    n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
    n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
    n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
    n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
    n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
    n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
    n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
    n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
    n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
    n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
    n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
    n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
    n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
    n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
    n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
    n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
    n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
    n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
    n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
    n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
    n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
    n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
    n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
    n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
    n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
    n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
    n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
    n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
    n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
    n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
    n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
    n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
    n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
    n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
    n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
    n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
    n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
    n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
    n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
    n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
    n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
    n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
    n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
    n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
    n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
    n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
    n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
    n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
    n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
    n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
    n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
    n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
    n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
    n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
    n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
    n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
    n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
    n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
    n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
    n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
    n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
    n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
    n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
    n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
    n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
    n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
    n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
    n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
    n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
    n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
    n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
    n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
    n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
    n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
    n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
    n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
    n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
    n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
    n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n921,
    n925_1, n929_1, n934_1, n939_1, n943, n947, n952_1, n956_1, n960_1,
    n964_1, n969, n973, n978_1, n982_1, n986_1, n990_1, n994_1, n998_1,
    n1002_1, n1007, n1011, n1015, n1019, n1023, n1027, n1031, n1035, n1039,
    n1043, n1047, n1051, n1056_1, n1060_1, n1064_1, n1069, n1073, n1077,
    n1081, n1086_1, n1090_1, n1094_1, n1098_1, n1102_1, n1106_1, n1110_1,
    n1114_1, n1118_1, n1123, n1127, n1131, n1135, n1139, n1143, n1147,
    n1151, n1155, n1159, n1163, n1167_1, n1172, n1176, n1180, n1185, n1189,
    n1193, n1197, n1202, n1206, n1210, n1214, n1218, n1222, n1226, n1230,
    n1234, n1239, n1243, n1247, n1251, n1255, n1259, n1263, n1267, n1271,
    n1275, n1279, n1283, n1288, n1292_1, n1296_1, n1301_1, n1305_1,
    n1309_1, n1313_1, n1318_1, n1322_1, n1326_1, n1330_1, n1334_1, n1338_1,
    n1342_1, n1346_1, n1350_1, n1355_1, n1359_1, n1363_1, n1367_1, n1371_1,
    n1375_1, n1379_1, n1383_1, n1387_1, n1391_1, n1395_1, n1400_1, n1404_1,
    n1408_1, n1412_1, n1416_1, n1421_1, n1425_1, n1429_1, n1433_1, n1437_1,
    n1441_1, n1446_1, n1451_1, n1456_1, n1460_1, n1464_1, n1469_1, n1473_1,
    n1477_1, n1482_1, n1486_1, n1490_1, n1495_1, n1499_1, n1503_1, n1507_1,
    n1511_1, n1515, n1520_1, n1524_1, n1528_1, n1532_1, n1536_1, n1540_1,
    n1544_1, n1548_1, n1552_1, n1557_1, n1561_1, n1565_1, n1569_1, n1573_1,
    n1577_1, n1581_1, n1586_1, n1590_1, n1594_1, n1599_1, n1603_1, n1607_1,
    n1611_1, n1615_1, n1619_1, n1623_1, n1627_1, n1631_1, n1636_1, n1640_1,
    n1644_1, n1648_1, n1652_1, n1656_1, n1660_1, n1664_1, n1668_1, n1672_1,
    n1676_1, n1681_1, n1686_1, n1690_1, n1694_1, n1698_1, n1703_1, n1707_1,
    n1711_1, n1716_1, n1720_1, n1724_1, n1729_1, n1733_1, n1737_1, n1741_1,
    n1745, n1749, n1754_1, n1758_1, n1762_1, n1766_1, n1770_1, n1774_1,
    n1778_1, n1782_1, n1786_1, n1790_1, n1794_1, n1799, n1803, n1807,
    n1811, n1815, n1820_1, n1824_1, n1828_1, n1833, n1837, n1841, n1845,
    n1849, n1853;
  assign Pnew_count_3_ = ~n1142;
  assign Pnew_count_2_ = ~n1143_1;
  assign Pnew_count_1_ = ~n1144;
  assign Pnew_count_0_ = ~n1145;
  assign Pdata_ready_0_ = ~n1141;
  assign n1137 = ~Pstart_0_ | Pencrypt_0_;
  assign n1138 = ~Pstart_0_ | ~Pencrypt_0_;
  assign n1139_1 = n1597 | Pstart_0_ | Pencrypt_0_;
  assign n1140 = n1597 & ~Pstart_0_ & ~Pencrypt_0_;
  assign n1141 = n2049 & (Pstart_0_ | n2050);
  assign n1142 = n1137 & (Pstart_0_ | n2058);
  assign n1143_1 = ~n2053 & (Pencrypt_0_ | n1595) & n2054;
  assign n1144 = n1137 & n2051 & (~Pcount_0_ | n2052);
  assign n1145 = n1137 & (Pstart_0_ | Pcount_0_);
  assign n1146 = n1823 & (~Pkey_62_ | n1138) & n1824;
  assign n1387_1 = ~n1146;
  assign n1148 = n1821 & (~Pkey_195_ | n1138) & n1822;
  assign n1391_1 = ~n1148;
  assign n1150 = n1819 & (~Pkey_203_ | n1138) & n1820;
  assign n1395_1 = ~n1150;
  assign n1152 = n1817 & (~Pkey_211_ | n1138) & n1818;
  assign n1400_1 = ~n1152;
  assign n1154 = n1815_1 & (~Pkey_219_ | n1138) & n1816;
  assign n1404_1 = ~n1154;
  assign n1156 = n1813 & (~Pkey_196_ | n1138) & n1814;
  assign n1408_1 = ~n1156;
  assign n1158 = n1811_1 & (~Pkey_204_ | n1138) & n1812;
  assign n1412_1 = ~n1158;
  assign n1160 = n1809 & (~Pkey_212_ | n1138) & n1810;
  assign n1416_1 = ~n1160;
  assign n1162 = n1807_1 & (~Pkey_220_ | n1138) & n1808;
  assign n1421_1 = ~n1162;
  assign n1164 = n1805 & (~Pkey_228_ | n1138) & n1806;
  assign n1425_1 = ~n1164;
  assign n1166 = n1803_1 & (~Pkey_172_ | n1138) & n1804;
  assign n1429_1 = ~n1166;
  assign n1168 = n1801 & (~Pkey_244_ | n1138) & n1802;
  assign n1433_1 = ~n1168;
  assign n1170 = n1799_1 & (~Pkey_252_ | n1138) & n1800;
  assign n1437_1 = ~n1170;
  assign n1172_1 = n1797 & (~Pkey_197_ | n1138) & n1798;
  assign n1441_1 = ~n1172_1;
  assign n1174 = n1795 & (~Pkey_205_ | n1138) & n1796;
  assign n1446_1 = ~n1174;
  assign n1176_1 = n1793 & (~Pkey_213_ | n1138) & n1794;
  assign n1451_1 = ~n1176_1;
  assign n1178 = n1791 & (~Pkey_221_ | n1138) & n1792;
  assign n1456_1 = ~n1178;
  assign n1180_1 = n1789 & (~Pkey_229_ | n1138) & n1790;
  assign n1460_1 = ~n1180_1;
  assign n1182 = n1787 & (~Pkey_237_ | n1138) & n1788;
  assign n1464_1 = ~n1182;
  assign n1184 = n1785 & (~Pkey_245_ | n1138) & n1786;
  assign n1469_1 = ~n1184;
  assign n1186 = n1783 & (~Pkey_253_ | n1138) & n1784;
  assign n1473_1 = ~n1186;
  assign n1188 = n1781 & (~Pkey_198_ | n1138) & n1782;
  assign n1477_1 = ~n1188;
  assign n1190 = n1779 & (~Pkey_206_ | n1138) & n1780;
  assign n1482_1 = ~n1190;
  assign n1192 = n1777 & (~Pkey_214_ | n1138) & n1778;
  assign n1486_1 = ~n1192;
  assign n1194 = n1775 & (~Pkey_222_ | n1138) & n1776;
  assign n1490_1 = ~n1194;
  assign n1196 = n1773 & (~Pkey_230_ | n1138) & n1774;
  assign n1495_1 = ~n1196;
  assign n1198 = n1771 & (~Pkey_238_ | n1138) & n1772;
  assign n1499_1 = ~n1198;
  assign n1200 = n1769 & (~Pkey_246_ | n1138) & n1770;
  assign n1503_1 = ~n1200;
  assign n1202_1 = n1767 & (~Pkey_254_ | n1138) & n1768;
  assign n1507_1 = ~n1202_1;
  assign n1204 = n1765 & (~Pkey_131_ | n1138) & n1766;
  assign n1511_1 = ~n1204;
  assign n1206_1 = n1763 & (~Pkey_139_ | n1138) & n1764;
  assign n1515 = ~n1206_1;
  assign n1208 = n1761 & (~Pkey_147_ | n1138) & n1762;
  assign n1520_1 = ~n1208;
  assign n1210_1 = n1759 & (~Pkey_155_ | n1138) & n1760;
  assign n1524_1 = ~n1210_1;
  assign n1212 = n1757 & (~Pkey_132_ | n1138) & n1758;
  assign n1528_1 = ~n1212;
  assign n1214_1 = n1755 & (~Pkey_140_ | n1138) & n1756;
  assign n1532_1 = ~n1214_1;
  assign n1216 = n1753 & (~Pkey_148_ | n1138) & n1754;
  assign n1536_1 = ~n1216;
  assign n1218_1 = n1751 & (~Pkey_156_ | n1138) & n1752;
  assign n1540_1 = ~n1218_1;
  assign n1220 = n1749_1 & (~Pkey_164_ | n1138) & n1750;
  assign n1544_1 = ~n1220;
  assign n1222_1 = n1747 & (~Pkey_172_ | n1138) & n1748;
  assign n1548_1 = ~n1222_1;
  assign n1224 = n1745_1 & (~Pkey_180_ | n1138) & n1746;
  assign n1552_1 = ~n1224;
  assign n1226_1 = n1743 & (~Pkey_188_ | n1138) & n1744;
  assign n1557_1 = ~n1226_1;
  assign n1228 = n1741 & (~Pkey_133_ | n1138) & n1742;
  assign n1561_1 = ~n1228;
  assign n1230_1 = n1739 & (~Pkey_141_ | n1138) & n1740;
  assign n1565_1 = ~n1230_1;
  assign n1232 = n1737 & (~Pkey_149_ | n1138) & n1738;
  assign n1569_1 = ~n1232;
  assign n1234_1 = n1735 & (~Pkey_157_ | n1138) & n1736;
  assign n1573_1 = ~n1234_1;
  assign n1236 = n1733 & (~Pkey_165_ | n1138) & n1734;
  assign n1577_1 = ~n1236;
  assign n1238 = n1731 & (~Pkey_173_ | n1138) & n1732;
  assign n1581_1 = ~n1238;
  assign n1240 = n1729 & (~Pkey_181_ | n1138) & n1730;
  assign n1586_1 = ~n1240;
  assign n1242 = n1727 & (~Pkey_189_ | n1138) & n1728;
  assign n1590_1 = ~n1242;
  assign n1244 = n1725 & (~Pkey_134_ | n1138) & n1726;
  assign n1594_1 = ~n1244;
  assign n1246 = n1723 & (~Pkey_142_ | n1138) & n1724;
  assign n1599_1 = ~n1246;
  assign n1248 = n1721 & (~Pkey_150_ | n1138) & n1722;
  assign n1603_1 = ~n1248;
  assign n1250 = n1719 & (~Pkey_158_ | n1138) & n1720;
  assign n1607_1 = ~n1250;
  assign n1252 = n1717 & (~Pkey_166_ | n1138) & n1718;
  assign n1611_1 = ~n1252;
  assign n1254 = n1715 & (~Pkey_174_ | n1138) & n1716;
  assign n1615_1 = ~n1254;
  assign n1256 = n1713 & (~Pkey_182_ | n1138) & n1714;
  assign n1619_1 = ~n1256;
  assign n1258 = n1711 & (~Pkey_190_ | n1138) & n1712;
  assign n1623_1 = ~n1258;
  assign n1260 = n1709 & (~Pkey_67_ | n1138) & n1710;
  assign n1627_1 = ~n1260;
  assign n1262 = n1707 & (~Pkey_75_ | n1138) & n1708;
  assign n1631_1 = ~n1262;
  assign n1264 = n1705 & (~Pkey_83_ | n1138) & n1706;
  assign n1636_1 = ~n1264;
  assign n1266 = n1703 & (~Pkey_91_ | n1138) & n1704;
  assign n1640_1 = ~n1266;
  assign n1268 = n1701 & (~Pkey_68_ | n1138) & n1702;
  assign n1644_1 = ~n1268;
  assign n1270 = n1699 & (~Pkey_76_ | n1138) & n1700;
  assign n1648_1 = ~n1270;
  assign n1272 = n1697 & (~Pkey_84_ | n1138) & n1698;
  assign n1652_1 = ~n1272;
  assign n1274 = n1695 & (~Pkey_92_ | n1138) & n1696;
  assign n1656_1 = ~n1274;
  assign n1276 = n1693 & (~Pkey_100_ | n1138) & n1694;
  assign n1660_1 = ~n1276;
  assign n1278 = n1691 & (~Pkey_44_ | n1138) & n1692;
  assign n1664_1 = ~n1278;
  assign n1280 = n1689 & (~Pkey_116_ | n1138) & n1690;
  assign n1668_1 = ~n1280;
  assign n1282 = n1687 & (~Pkey_124_ | n1138) & n1688;
  assign n1672_1 = ~n1282;
  assign n1284 = n1685 & (~Pkey_69_ | n1138) & n1686;
  assign n1676_1 = ~n1284;
  assign n1286 = n1683 & (~Pkey_77_ | n1138) & n1684;
  assign n1681_1 = ~n1286;
  assign n1288_1 = n1681 & (~Pkey_85_ | n1138) & n1682;
  assign n1686_1 = ~n1288_1;
  assign n1290 = n1679 & (~Pkey_93_ | n1138) & n1680;
  assign n1690_1 = ~n1290;
  assign n1292 = n1677 & (~Pkey_101_ | n1138) & n1678;
  assign n1694_1 = ~n1292;
  assign n1294 = n1675 & (~Pkey_109_ | n1138) & n1676;
  assign n1698_1 = ~n1294;
  assign n1296 = n1673 & (~Pkey_117_ | n1138) & n1674;
  assign n1703_1 = ~n1296;
  assign n1298 = n1671 & (~Pkey_125_ | n1138) & n1672;
  assign n1707_1 = ~n1298;
  assign n1300 = n1669 & (~Pkey_70_ | n1138) & n1670;
  assign n1711_1 = ~n1300;
  assign n1302 = n1667 & (~Pkey_78_ | n1138) & n1668;
  assign n1716_1 = ~n1302;
  assign n1304 = n1665 & (~Pkey_86_ | n1138) & n1666;
  assign n1720_1 = ~n1304;
  assign n1306 = n1663 & (~Pkey_94_ | n1138) & n1664;
  assign n1724_1 = ~n1306;
  assign n1308 = n1661 & (~Pkey_102_ | n1138) & n1662;
  assign n1729_1 = ~n1308;
  assign n1310 = n1659 & (~Pkey_110_ | n1138) & n1660;
  assign n1733_1 = ~n1310;
  assign n1312 = n1657 & (~Pkey_118_ | n1138) & n1658;
  assign n1737_1 = ~n1312;
  assign n1314 = n1655 & (~Pkey_126_ | n1138) & n1656;
  assign n1741_1 = ~n1314;
  assign n1316 = n1653 & (~Pkey_3_ | n1138) & n1654;
  assign n1745 = ~n1316;
  assign n1318 = n1651 & (~Pkey_11_ | n1138) & n1652;
  assign n1749 = ~n1318;
  assign n1320 = n1649 & (~Pkey_19_ | n1138) & n1650;
  assign n1754_1 = ~n1320;
  assign n1322 = n1647 & (~Pkey_27_ | n1138) & n1648;
  assign n1758_1 = ~n1322;
  assign n1324 = n1645 & (~Pkey_4_ | n1138) & n1646;
  assign n1762_1 = ~n1324;
  assign n1326 = n1643 & (~Pkey_12_ | n1138) & n1644;
  assign n1766_1 = ~n1326;
  assign n1328 = n1641 & (~Pkey_20_ | n1138) & n1642;
  assign n1770_1 = ~n1328;
  assign n1330 = n1639 & (~Pkey_28_ | n1138) & n1640;
  assign n1774_1 = ~n1330;
  assign n1332 = n1637 & (~Pkey_36_ | n1138) & n1638;
  assign n1778_1 = ~n1332;
  assign n1334 = n1635 & (~Pkey_44_ | n1138) & n1636;
  assign n1782_1 = ~n1334;
  assign n1336 = n1633 & (~Pkey_52_ | n1138) & n1634;
  assign n1786_1 = ~n1336;
  assign n1338 = n1631 & (~Pkey_60_ | n1138) & n1632;
  assign n1790_1 = ~n1338;
  assign n1340 = n1629 & (~Pkey_5_ | n1138) & n1630;
  assign n1794_1 = ~n1340;
  assign n1342 = n1627 & (~Pkey_13_ | n1138) & n1628;
  assign n1799 = ~n1342;
  assign n1344 = n1625 & (~Pkey_21_ | n1138) & n1626;
  assign n1803 = ~n1344;
  assign n1346 = n1623 & (~Pkey_29_ | n1138) & n1624;
  assign n1807 = ~n1346;
  assign n1348 = n1621 & (~Pkey_37_ | n1138) & n1622;
  assign n1811 = ~n1348;
  assign n1350 = n1619 & (~Pkey_45_ | n1138) & n1620;
  assign n1815 = ~n1350;
  assign n1352 = n1617 & (~Pkey_53_ | n1138) & n1618;
  assign n1820_1 = ~n1352;
  assign n1354 = n1615 & (~Pkey_61_ | n1138) & n1616;
  assign n1824_1 = ~n1354;
  assign n1356 = n1613 & (~Pkey_6_ | n1138) & n1614;
  assign n1828_1 = ~n1356;
  assign n1358 = n1611 & (~Pkey_14_ | n1138) & n1612;
  assign n1833 = ~n1358;
  assign n1360 = n1609 & (~Pkey_22_ | n1138) & n1610;
  assign n1837 = ~n1360;
  assign n1362 = n1607 & (~Pkey_30_ | n1138) & n1608;
  assign n1841 = ~n1362;
  assign n1364 = n1605 & (~Pkey_38_ | n1138) & n1606;
  assign n1845 = ~n1364;
  assign n1366 = n1603 & (~Pkey_46_ | n1138) & n1604;
  assign n1849 = ~n1366;
  assign n1368 = n1601 & (~Pkey_54_ | n1138) & n1602;
  assign n1853 = ~n1368;
  assign n1370 = n2047 & (~Pkey_56_ | n1138) & n2048;
  assign n921 = ~n1370;
  assign n1372 = n2045 & (~Pkey_227_ | n1138) & n2046;
  assign n925_1 = ~n1372;
  assign n1374 = n2043 & (~Pkey_235_ | n1138) & n2044;
  assign n929_1 = ~n1374;
  assign n1376 = n2041 & (~Pkey_243_ | n1138) & n2042;
  assign n934_1 = ~n1376;
  assign n1378 = n2039 & (~Pkey_251_ | n1138) & n2040;
  assign n939_1 = ~n1378;
  assign n1380 = n2037 & (~Pkey_194_ | n1138) & n2038;
  assign n943 = ~n1380;
  assign n1382 = n2035 & (~Pkey_202_ | n1138) & n2036;
  assign n947 = ~n1382;
  assign n1384 = n2033 & (~Pkey_210_ | n1138) & n2034;
  assign n952_1 = ~n1384;
  assign n1386 = n2031 & (~Pkey_218_ | n1138) & n2032;
  assign n956_1 = ~n1386;
  assign n1388 = n2029 & (~Pkey_226_ | n1138) & n2030;
  assign n960_1 = ~n1388;
  assign n1390 = n2027 & (~Pkey_234_ | n1138) & n2028;
  assign n964_1 = ~n1390;
  assign n1392 = n2025 & (~Pkey_242_ | n1138) & n2026;
  assign n969 = ~n1392;
  assign n1394 = n2023 & (~Pkey_250_ | n1138) & n2024;
  assign n973 = ~n1394;
  assign n1396 = n2021 & (~Pkey_193_ | n1138) & n2022;
  assign n978_1 = ~n1396;
  assign n1398 = n2019 & (~Pkey_201_ | n1138) & n2020;
  assign n982_1 = ~n1398;
  assign n1400 = n2017 & (~Pkey_209_ | n1138) & n2018;
  assign n986_1 = ~n1400;
  assign n1402 = n2015 & (~Pkey_217_ | n1138) & n2016;
  assign n990_1 = ~n1402;
  assign n1404 = n2013 & (~Pkey_225_ | n1138) & n2014;
  assign n994_1 = ~n1404;
  assign n1406 = n2011 & (~Pkey_233_ | n1138) & n2012;
  assign n998_1 = ~n1406;
  assign n1408 = n2009 & (~Pkey_241_ | n1138) & n2010;
  assign n1002_1 = ~n1408;
  assign n1410 = n2007 & (~Pkey_249_ | n1138) & n2008;
  assign n1007 = ~n1410;
  assign n1412 = n2005 & (~Pkey_192_ | n1138) & n2006;
  assign n1011 = ~n1412;
  assign n1414 = n2003 & (~Pkey_200_ | n1138) & n2004;
  assign n1015 = ~n1414;
  assign n1416 = n2001 & (~Pkey_208_ | n1138) & n2002;
  assign n1019 = ~n1416;
  assign n1418 = n1999 & (~Pkey_216_ | n1138) & n2000;
  assign n1023 = ~n1418;
  assign n1420 = n1997 & (~Pkey_224_ | n1138) & n1998;
  assign n1027 = ~n1420;
  assign n1422 = n1995 & (~Pkey_232_ | n1138) & n1996;
  assign n1031 = ~n1422;
  assign n1424 = n1993 & (~Pkey_240_ | n1138) & n1994;
  assign n1035 = ~n1424;
  assign n1426 = n1991 & (~Pkey_248_ | n1138) & n1992;
  assign n1039 = ~n1426;
  assign n1428 = n1989 & (~Pkey_163_ | n1138) & n1990;
  assign n1043 = ~n1428;
  assign n1430 = n1987 & (~Pkey_171_ | n1138) & n1988;
  assign n1047 = ~n1430;
  assign n1432 = n1985 & (~Pkey_179_ | n1138) & n1986;
  assign n1051 = ~n1432;
  assign n1434 = n1983 & (~Pkey_187_ | n1138) & n1984;
  assign n1056_1 = ~n1434;
  assign n1436 = n1981 & (~Pkey_130_ | n1138) & n1982;
  assign n1060_1 = ~n1436;
  assign n1438 = n1979 & (~Pkey_138_ | n1138) & n1980;
  assign n1064_1 = ~n1438;
  assign n1440 = n1977 & (~Pkey_146_ | n1138) & n1978;
  assign n1069 = ~n1440;
  assign n1442 = n1975 & (~Pkey_154_ | n1138) & n1976;
  assign n1073 = ~n1442;
  assign n1444 = n1973 & (~Pkey_162_ | n1138) & n1974;
  assign n1077 = ~n1444;
  assign n1446 = n1971 & (~Pkey_170_ | n1138) & n1972;
  assign n1081 = ~n1446;
  assign n1448 = n1969 & (~Pkey_178_ | n1138) & n1970;
  assign n1086_1 = ~n1448;
  assign n1450 = n1967 & (~Pkey_186_ | n1138) & n1968;
  assign n1090_1 = ~n1450;
  assign n1452 = n1965 & (~Pkey_129_ | n1138) & n1966;
  assign n1094_1 = ~n1452;
  assign n1454 = n1963 & (~Pkey_137_ | n1138) & n1964;
  assign n1098_1 = ~n1454;
  assign n1456 = n1961 & (~Pkey_145_ | n1138) & n1962;
  assign n1102_1 = ~n1456;
  assign n1458 = n1959 & (~Pkey_153_ | n1138) & n1960;
  assign n1106_1 = ~n1458;
  assign n1460 = n1957 & (~Pkey_161_ | n1138) & n1958;
  assign n1110_1 = ~n1460;
  assign n1462 = n1955 & (~Pkey_169_ | n1138) & n1956;
  assign n1114_1 = ~n1462;
  assign n1464 = n1953 & (~Pkey_177_ | n1138) & n1954;
  assign n1118_1 = ~n1464;
  assign n1466 = n1951 & (~Pkey_185_ | n1138) & n1952;
  assign n1123 = ~n1466;
  assign n1468 = n1949 & (~Pkey_128_ | n1138) & n1950;
  assign n1127 = ~n1468;
  assign n1470 = n1947 & (~Pkey_136_ | n1138) & n1948;
  assign n1131 = ~n1470;
  assign n1472 = n1945 & (~Pkey_144_ | n1138) & n1946;
  assign n1135 = ~n1472;
  assign n1474 = n1943 & (~Pkey_152_ | n1138) & n1944;
  assign n1139 = ~n1474;
  assign n1476 = n1941 & (~Pkey_160_ | n1138) & n1942;
  assign n1143 = ~n1476;
  assign n1478 = n1939 & (~Pkey_168_ | n1138) & n1940;
  assign n1147 = ~n1478;
  assign n1480 = n1937 & (~Pkey_176_ | n1138) & n1938;
  assign n1151 = ~n1480;
  assign n1482 = n1935 & (~Pkey_184_ | n1138) & n1936;
  assign n1155 = ~n1482;
  assign n1484 = n1933 & (~Pkey_99_ | n1138) & n1934;
  assign n1159 = ~n1484;
  assign n1486 = n1931 & (~Pkey_107_ | n1138) & n1932;
  assign n1163 = ~n1486;
  assign n1488 = n1929 & (~Pkey_115_ | n1138) & n1930;
  assign n1167_1 = ~n1488;
  assign n1490 = n1927 & (~Pkey_123_ | n1138) & n1928;
  assign n1172 = ~n1490;
  assign n1492 = n1925 & (~Pkey_66_ | n1138) & n1926;
  assign n1176 = ~n1492;
  assign n1494 = n1923 & (~Pkey_74_ | n1138) & n1924;
  assign n1180 = ~n1494;
  assign n1496 = n1921 & (~Pkey_82_ | n1138) & n1922;
  assign n1185 = ~n1496;
  assign n1498 = n1919 & (~Pkey_90_ | n1138) & n1920;
  assign n1189 = ~n1498;
  assign n1500 = n1917 & (~Pkey_98_ | n1138) & n1918;
  assign n1193 = ~n1500;
  assign n1502 = n1915 & (~Pkey_106_ | n1138) & n1916;
  assign n1197 = ~n1502;
  assign n1504 = n1913 & (~Pkey_114_ | n1138) & n1914;
  assign n1202 = ~n1504;
  assign n1506 = n1911 & (~Pkey_122_ | n1138) & n1912;
  assign n1206 = ~n1506;
  assign n1508 = n1909 & (~Pkey_65_ | n1138) & n1910;
  assign n1210 = ~n1508;
  assign n1510 = n1907 & (~Pkey_73_ | n1138) & n1908;
  assign n1214 = ~n1510;
  assign n1512 = n1905 & (~Pkey_81_ | n1138) & n1906;
  assign n1218 = ~n1512;
  assign n1514 = n1903 & (~Pkey_89_ | n1138) & n1904;
  assign n1222 = ~n1514;
  assign n1516 = n1901 & (~Pkey_97_ | n1138) & n1902;
  assign n1226 = ~n1516;
  assign n1518 = n1899 & (~Pkey_105_ | n1138) & n1900;
  assign n1230 = ~n1518;
  assign n1520 = n1897 & (~Pkey_113_ | n1138) & n1898;
  assign n1234 = ~n1520;
  assign n1522 = n1895 & (~Pkey_121_ | n1138) & n1896;
  assign n1239 = ~n1522;
  assign n1524 = n1893 & (~Pkey_64_ | n1138) & n1894;
  assign n1243 = ~n1524;
  assign n1526 = n1891 & (~Pkey_72_ | n1138) & n1892;
  assign n1247 = ~n1526;
  assign n1528 = n1889 & (~Pkey_80_ | n1138) & n1890;
  assign n1251 = ~n1528;
  assign n1530 = n1887 & (~Pkey_88_ | n1138) & n1888;
  assign n1255 = ~n1530;
  assign n1532 = n1885 & (~Pkey_96_ | n1138) & n1886;
  assign n1259 = ~n1532;
  assign n1534 = n1883 & (~Pkey_104_ | n1138) & n1884;
  assign n1263 = ~n1534;
  assign n1536 = n1881 & (~Pkey_112_ | n1138) & n1882;
  assign n1267 = ~n1536;
  assign n1538 = n1879 & (~Pkey_120_ | n1138) & n1880;
  assign n1271 = ~n1538;
  assign n1540 = n1877 & (~Pkey_35_ | n1138) & n1878;
  assign n1275 = ~n1540;
  assign n1542 = n1875 & (~Pkey_43_ | n1138) & n1876;
  assign n1279 = ~n1542;
  assign n1544 = n1873 & (~Pkey_51_ | n1138) & n1874;
  assign n1283 = ~n1544;
  assign n1546 = n1871 & (~Pkey_59_ | n1138) & n1872;
  assign n1288 = ~n1546;
  assign n1548 = n1869 & (~Pkey_2_ | n1138) & n1870;
  assign n1292_1 = ~n1548;
  assign n1550 = n1867 & (~Pkey_10_ | n1138) & n1868;
  assign n1296_1 = ~n1550;
  assign n1552 = n1865 & (~Pkey_18_ | n1138) & n1866;
  assign n1301_1 = ~n1552;
  assign n1554 = n1863 & (~Pkey_26_ | n1138) & n1864;
  assign n1305_1 = ~n1554;
  assign n1556 = n1861 & (~Pkey_34_ | n1138) & n1862;
  assign n1309_1 = ~n1556;
  assign n1558 = n1859 & (~Pkey_42_ | n1138) & n1860;
  assign n1313_1 = ~n1558;
  assign n1560 = n1857 & (~Pkey_50_ | n1138) & n1858;
  assign n1318_1 = ~n1560;
  assign n1562 = n1855 & (~Pkey_58_ | n1138) & n1856;
  assign n1322_1 = ~n1562;
  assign n1564 = n1853_1 & (~Pkey_1_ | n1138) & n1854;
  assign n1326_1 = ~n1564;
  assign n1566 = n1851 & (~Pkey_9_ | n1138) & n1852;
  assign n1330_1 = ~n1566;
  assign n1568 = n1849_1 & (~Pkey_17_ | n1138) & n1850;
  assign n1334_1 = ~n1568;
  assign n1570 = n1847 & (~Pkey_25_ | n1138) & n1848;
  assign n1338_1 = ~n1570;
  assign n1572 = n1845_1 & (~Pkey_33_ | n1138) & n1846;
  assign n1342_1 = ~n1572;
  assign n1574 = n1843 & (~Pkey_41_ | n1138) & n1844;
  assign n1346_1 = ~n1574;
  assign n1576 = n1841_1 & (~Pkey_49_ | n1138) & n1842;
  assign n1350_1 = ~n1576;
  assign n1578 = n1839 & (~Pkey_57_ | n1138) & n1840;
  assign n1355_1 = ~n1578;
  assign n1580 = n1837_1 & (~Pkey_0_ | n1138) & n1838;
  assign n1359_1 = ~n1580;
  assign n1582 = n1835 & (~Pkey_8_ | n1138) & n1836;
  assign n1363_1 = ~n1582;
  assign n1584 = n1833_1 & (~Pkey_16_ | n1138) & n1834;
  assign n1367_1 = ~n1584;
  assign n1586 = n1831 & (~Pkey_24_ | n1138) & n1832;
  assign n1371_1 = ~n1586;
  assign n1588 = n1829 & (~Pkey_32_ | n1138) & n1830;
  assign n1375_1 = ~n1588;
  assign n1590 = n1827 & (~Pkey_40_ | n1138) & n1828;
  assign n1379_1 = ~n1590;
  assign n1592 = n1825 & (~Pkey_48_ | n1138) & n1826;
  assign n1383_1 = ~n1592;
  assign n1594 = Pcount_3_ | Pcount_1_ | Pcount_2_;
  assign n1595 = Pcount_0_ | Pcount_1_ | Pcount_2_;
  assign n1596 = ~Pcount_2_ | ~Pcount_1_ | ~Pcount_0_;
  assign n1597 = n1594 & n1595 & (~Pcount_3_ | n1596);
  assign n1598 = ~Pcount_3_ | ~Pcount_2_ | ~Pcount_1_ | Pcount_0_;
  assign n1599 = Pcount_3_ | n1596;
  assign n1600 = n1598 & n1599 & (Pcount_3_ | n1595);
  assign n1601 = n2179 & (~PKSi_118_ | ~PKSi_4_ | n2172);
  assign n1602 = (~Pkey_62_ | n1137) & n2180;
  assign n1603 = n2181 & (~PKSi_102_ | ~PKSi_23_ | n2172);
  assign n1604 = (~Pkey_54_ | n1137) & n2182;
  assign n1605 = n2183 & (~PKSi_98_ | ~PKSi_6_ | n2172);
  assign n1606 = (~Pkey_46_ | n1137) & n2184;
  assign n1607 = n2185 & (~PKSi_119_ | ~PKSi_15_ | n2172);
  assign n1608 = (~Pkey_38_ | n1137) & n2186;
  assign n1609 = n2187 & (~PKSi_106_ | ~PKSi_5_ | n2172);
  assign n1610 = (~Pkey_30_ | n1137) & n2188;
  assign n1611 = n2189 & (~PKSi_112_ | ~PKSi_9_ | n2172);
  assign n1612 = (~Pkey_22_ | n1137) & n2190;
  assign n1613 = n2191 & (~PKSi_19_ | ~N_N2986 | n2172);
  assign n1614 = (~Pkey_14_ | n1137) & n2192;
  assign n1615 = n2193 & (~PKSi_117_ | ~PKSi_17_ | n2172);
  assign n1616 = (~Pkey_6_ | n1137) & n2194;
  assign n1617 = n2195 & (~PKSi_99_ | n2172 | ~N_N2853);
  assign n1618 = (~Pkey_61_ | n1137) & n2196;
  assign n1619 = n2197 & (~PKSi_11_ | ~N_N2982 | n2172);
  assign n1620 = (~Pkey_53_ | n1137) & n2198;
  assign n1621 = n2199 & (~PKSi_110_ | ~PKSi_2_ | n2172);
  assign n1622 = (~Pkey_45_ | n1137) & n2200;
  assign n1623 = n2201 & (~PKSi_103_ | ~PKSi_14_ | n2172);
  assign n1624 = (~Pkey_37_ | n1137) & n2202;
  assign n1625 = n2203 & (~PKSi_96_ | ~PKSi_22_ | n2172);
  assign n1626 = (~Pkey_29_ | n1137) & n2204;
  assign n1627 = n2205 & (~PKSi_115_ | ~PKSi_0_ | n2172);
  assign n1628 = (~Pkey_21_ | n1137) & n2206;
  assign n1629 = n2207 & (~PKSi_8_ | ~N_N2976 | n2172);
  assign n1630 = (~Pkey_13_ | n1137) & n2208;
  assign n1631 = n2209 & (~PKSi_108_ | ~PKSi_18_ | n2172);
  assign n1632 = (~Pkey_5_ | n1137) & n2210;
  assign n1633 = n2211 & (~PKSi_105_ | ~PKSi_1_ | n2172);
  assign n1634 = (~Pkey_60_ | n1137) & n2212;
  assign n1635 = n2213 & (~PKSi_114_ | n2172 | ~N_N2843);
  assign n1636 = (~Pkey_52_ | n1137) & n2214;
  assign n1637 = n2215 & (~PKSi_100_ | ~PKSi_13_ | n2172);
  assign n1638 = (~Pkey_44_ | n1137) & n2216;
  assign n1639 = n2217 & (~PKSi_107_ | ~PKSi_21_ | n2172);
  assign n1640 = (~Pkey_36_ | n1137) & n2218;
  assign n1641 = n2219 & (~PKSi_109_ | ~PKSi_10_ | n2172);
  assign n1642 = (~Pkey_28_ | n1137) & n2220;
  assign n1643 = n2221 & (~PKSi_116_ | n2172 | ~N_N2838);
  assign n1644 = (~Pkey_20_ | n1137) & n2222;
  assign n1645 = n2223 & (~PKSi_104_ | ~PKSi_12_ | n2172);
  assign n1646 = (~Pkey_12_ | n1137) & n2224;
  assign n1647 = n2225 & (~PKSi_97_ | ~PKSi_3_ | n2172);
  assign n1648 = (~Pkey_4_ | n1137) & n2226;
  assign n1649 = n2227 & (~PKSi_113_ | n2172 | ~N_N2834);
  assign n1650 = (~Pkey_27_ | n1137) & n2228;
  assign n1651 = n2229 & (~PKSi_16_ | ~N_N2964 | n2172);
  assign n1652 = (~Pkey_19_ | n1137) & n2230;
  assign n1653 = n2231 & (~PKSi_101_ | ~PKSi_20_ | n2172);
  assign n1654 = (~Pkey_11_ | n1137) & n2232;
  assign n1655 = n2233 & (~PKSi_111_ | ~PKSi_7_ | n2172);
  assign n1656 = (~Pkey_3_ | n1137) & n2234;
  assign n1657 = n2235 & (~PKSi_142_ | ~PKSi_28_ | n2172);
  assign n1658 = (~Pkey_126_ | n1137) & n2236;
  assign n1659 = n2237 & (~PKSi_126_ | ~PKSi_47_ | n2172);
  assign n1660 = (~Pkey_118_ | n1137) & n2238;
  assign n1661 = n2239 & (~PKSi_122_ | ~PKSi_30_ | n2172);
  assign n1662 = (~Pkey_110_ | n1137) & n2240;
  assign n1663 = n2241 & (~\[282]  | ~PKSi_39_ | n2172);
  assign n1664 = (~Pkey_102_ | n1137) & n2242;
  assign n1665 = n2243 & (~PKSi_130_ | ~PKSi_29_ | n2172);
  assign n1666 = (~Pkey_94_ | n1137) & n2244;
  assign n1667 = n2245 & (~PKSi_136_ | ~PKSi_33_ | n2172);
  assign n1668 = (~Pkey_86_ | n1137) & n2246;
  assign n1669 = n2247 & (~PKSi_43_ | ~N_N2954 | n2172);
  assign n1670 = (~Pkey_78_ | n1137) & n2248;
  assign n1671 = n2249 & (~PKSi_141_ | ~PKSi_41_ | n2172);
  assign n1672 = (~Pkey_70_ | n1137) & n2250;
  assign n1673 = n2251 & (~PKSi_123_ | n2172 | ~N_N2821);
  assign n1674 = (~Pkey_125_ | n1137) & n2252;
  assign n1675 = n2253 & (~PKSi_35_ | ~N_N2950 | n2172);
  assign n1676 = (~Pkey_117_ | n1137) & n2254;
  assign n1677 = n2255 & (~PKSi_134_ | ~PKSi_26_ | n2172);
  assign n1678 = (~Pkey_109_ | n1137) & n2256;
  assign n1679 = n2257 & (~PKSi_127_ | ~PKSi_38_ | n2172);
  assign n1680 = (~Pkey_101_ | n1137) & n2258;
  assign n1681 = n2259 & (~PKSi_120_ | ~PKSi_46_ | n2172);
  assign n1682 = (~Pkey_93_ | n1137) & n2260;
  assign n1683 = n2261 & (~PKSi_24_ | ~N_N2945 | n2172);
  assign n1684 = (~Pkey_85_ | n1137) & n2262;
  assign n1685 = n2263 & (~PKSi_32_ | ~N_N2943 | n2172);
  assign n1686 = (~Pkey_77_ | n1137) & n2264;
  assign n1687 = n2265 & (~PKSi_132_ | ~PKSi_42_ | n2172);
  assign n1688 = (~Pkey_69_ | n1137) & n2266;
  assign n1689 = n2267 & (~PKSi_129_ | ~PKSi_25_ | n2172);
  assign n1690 = (~Pkey_124_ | n1137) & n2268;
  assign n1691 = n2269 & (~PKSi_138_ | n2172 | ~N_N2811);
  assign n1692 = (~Pkey_116_ | n1137) & n2270;
  assign n1693 = n2271 & (~PKSi_124_ | ~PKSi_37_ | n2172);
  assign n1694 = (~Pkey_44_ | n1137) & n2272;
  assign n1695 = n2273 & (~PKSi_131_ | ~PKSi_45_ | n2172);
  assign n1696 = (~Pkey_100_ | n1137) & n2274;
  assign n1697 = n2275 & (~PKSi_133_ | ~PKSi_34_ | n2172);
  assign n1698 = (~Pkey_92_ | n1137) & n2276;
  assign n1699 = n2277 & (~PKSi_140_ | n2172 | ~N_N2806);
  assign n1700 = (~Pkey_84_ | n1137) & n2278;
  assign n1701 = n2279 & (~PKSi_128_ | ~PKSi_36_ | n2172);
  assign n1702 = (~Pkey_76_ | n1137) & n2280;
  assign n1703 = n2281 & (~PKSi_121_ | ~PKSi_27_ | n2172);
  assign n1704 = (~Pkey_68_ | n1137) & n2282;
  assign n1705 = n2283 & (~PKSi_137_ | n2172 | ~N_N2802);
  assign n1706 = (~Pkey_91_ | n1137) & n2284;
  assign n1707 = n2285 & (~PKSi_40_ | ~N_N2931 | n2172);
  assign n1708 = (~Pkey_83_ | n1137) & n2286;
  assign n1709 = n2287 & (~PKSi_125_ | ~PKSi_44_ | n2172);
  assign n1710 = (~Pkey_75_ | n1137) & n2288;
  assign n1711 = n2289 & (~PKSi_135_ | ~PKSi_31_ | n2172);
  assign n1712 = (~Pkey_67_ | n1137) & n2290;
  assign n1713 = n2291 & (~PKSi_166_ | ~PKSi_52_ | n2172);
  assign n1714 = (~Pkey_190_ | n1137) & n2292;
  assign n1715 = n2293 & (~PKSi_150_ | ~PKSi_71_ | n2172);
  assign n1716 = (~Pkey_182_ | n1137) & n2294;
  assign n1717 = n2295 & (~PKSi_146_ | ~PKSi_54_ | n2172);
  assign n1718 = (~Pkey_174_ | n1137) & n2296;
  assign n1719 = n2297 & (~PKSi_167_ | ~PKSi_63_ | n2172);
  assign n1720 = (~Pkey_166_ | n1137) & n2298;
  assign n1721 = n2299 & (~PKSi_154_ | ~PKSi_53_ | n2172);
  assign n1722 = (~Pkey_158_ | n1137) & n2300;
  assign n1723 = n2301 & (~PKSi_160_ | ~PKSi_57_ | n2172);
  assign n1724 = (~Pkey_150_ | n1137) & n2302;
  assign n1725 = n2303 & (~PKSi_67_ | ~N_N2921 | n2172);
  assign n1726 = (~Pkey_142_ | n1137) & n2304;
  assign n1727 = n2305 & (~PKSi_165_ | ~PKSi_65_ | n2172);
  assign n1728 = (~Pkey_134_ | n1137) & n2306;
  assign n1729 = n2307 & (~PKSi_147_ | n2172 | ~N_N2789);
  assign n1730 = (~Pkey_189_ | n1137) & n2308;
  assign n1731 = n2309 & (~PKSi_59_ | ~N_N2917 | n2172);
  assign n1732 = (~Pkey_181_ | n1137) & n2310;
  assign n1733 = n2311 & (~PKSi_158_ | ~PKSi_50_ | n2172);
  assign n1734 = (~Pkey_173_ | n1137) & n2312;
  assign n1735 = n2313 & (~PKSi_151_ | ~PKSi_62_ | n2172);
  assign n1736 = (~Pkey_165_ | n1137) & n2314;
  assign n1737 = n2315 & (~PKSi_144_ | ~PKSi_70_ | n2172);
  assign n1738 = (~Pkey_157_ | n1137) & n2316;
  assign n1739 = n2317 & (~PKSi_163_ | ~PKSi_48_ | n2172);
  assign n1740 = (~Pkey_149_ | n1137) & n2318;
  assign n1741 = n2319 & (~PKSi_153_ | ~PKSi_56_ | n2172);
  assign n1742 = (~Pkey_141_ | n1137) & n2320;
  assign n1743 = n2321 & (~PKSi_156_ | ~PKSi_66_ | n2172);
  assign n1744 = (~Pkey_133_ | n1137) & n2322;
  assign n1745_1 = n2323 & (~PKSi_49_ | ~N_N2909 | n2172);
  assign n1746 = (~Pkey_188_ | n1137) & n2324;
  assign n1747 = n2325 & (~PKSi_162_ | n2172 | ~N_N2779);
  assign n1748 = (~Pkey_180_ | n1137) & n2326;
  assign n1749_1 = n2327 & (~PKSi_148_ | ~PKSi_61_ | n2172);
  assign n1750 = (~Pkey_172_ | n1137) & n2328;
  assign n1751 = n2329 & (~PKSi_155_ | ~PKSi_69_ | n2172);
  assign n1752 = (~Pkey_164_ | n1137) & n2330;
  assign n1753 = n2331 & (~PKSi_157_ | ~PKSi_58_ | n2172);
  assign n1754 = (~Pkey_156_ | n1137) & n2332;
  assign n1755 = n2333 & (~PKSi_164_ | n2172 | ~N_N2774);
  assign n1756 = (~Pkey_148_ | n1137) & n2334;
  assign n1757 = n2335 & (~PKSi_152_ | ~PKSi_60_ | n2172);
  assign n1758 = (~Pkey_140_ | n1137) & n2336;
  assign n1759 = n2337 & (~PKSi_145_ | ~PKSi_51_ | n2172);
  assign n1760 = (~Pkey_132_ | n1137) & n2338;
  assign n1761 = n2339 & (~PKSi_161_ | n2172 | ~N_N2770);
  assign n1762 = (~Pkey_155_ | n1137) & n2340;
  assign n1763 = n2341 & (~PKSi_64_ | ~N_N2899 | n2172);
  assign n1764 = (~Pkey_147_ | n1137) & n2342;
  assign n1765 = n2343 & (~PKSi_149_ | ~PKSi_68_ | n2172);
  assign n1766 = (~Pkey_139_ | n1137) & n2344;
  assign n1767 = n2345 & (~PKSi_159_ | ~PKSi_55_ | n2172);
  assign n1768 = (~Pkey_131_ | n1137) & n2346;
  assign n1769 = n2347 & (~PKSi_190_ | ~PKSi_76_ | n2172);
  assign n1770 = (~Pkey_254_ | n1137) & n2348;
  assign n1771 = n2349 & (~PKSi_174_ | ~PKSi_95_ | n2172);
  assign n1772 = (~Pkey_246_ | n1137) & n2350;
  assign n1773 = n2351 & (~PKSi_170_ | ~PKSi_78_ | n2172);
  assign n1774 = (~Pkey_238_ | n1137) & n2352;
  assign n1775 = n2353 & (~\[234]  | ~PKSi_87_ | n2172);
  assign n1776 = (~Pkey_230_ | n1137) & n2354;
  assign n1777 = n2355 & (~PKSi_178_ | ~PKSi_77_ | n2172);
  assign n1778 = (~Pkey_222_ | n1137) & n2356;
  assign n1779 = n2357 & (~PKSi_184_ | ~PKSi_81_ | n2172);
  assign n1780 = (~Pkey_214_ | n1137) & n2358;
  assign n1781 = n2359 & (~PKSi_91_ | ~N_N2889 | n2172);
  assign n1782 = (~Pkey_206_ | n1137) & n2360;
  assign n1783 = n2361 & (~PKSi_189_ | ~PKSi_89_ | n2172);
  assign n1784 = (~Pkey_198_ | n1137) & n2362;
  assign n1785 = n2363 & (~PKSi_171_ | n2172 | ~N_N2757);
  assign n1786 = (~Pkey_253_ | n1137) & n2364;
  assign n1787 = n2365 & (~PKSi_83_ | ~N_N2885 | n2172);
  assign n1788 = (~Pkey_245_ | n1137) & n2366;
  assign n1789 = n2367 & (~PKSi_182_ | ~PKSi_74_ | n2172);
  assign n1790 = (~Pkey_237_ | n1137) & n2368;
  assign n1791 = n2369 & (~PKSi_175_ | ~PKSi_86_ | n2172);
  assign n1792 = (~Pkey_229_ | n1137) & n2370;
  assign n1793 = n2371 & (~PKSi_94_ | ~N_N2881 | n2172);
  assign n1794 = (~Pkey_221_ | n1137) & n2372;
  assign n1795 = n2373 & (~PKSi_72_ | ~N_N2879 | n2172);
  assign n1796 = (~Pkey_213_ | n1137) & n2374;
  assign n1797 = n2375 & (~PKSi_80_ | ~N_N2877 | n2172);
  assign n1798 = (~Pkey_205_ | n1137) & n2376;
  assign n1799_1 = n2377 & (~PKSi_180_ | n2172 | ~N_N2749);
  assign n1800 = (~Pkey_197_ | n1137) & n2378;
  assign n1801 = n2379 & (~PKSi_177_ | ~PKSi_73_ | n2172);
  assign n1802 = (~Pkey_252_ | n1137) & n2380;
  assign n1803_1 = n2381 & (~PKSi_186_ | n2172 | ~N_N2746);
  assign n1804 = (~Pkey_244_ | n1137) & n2382;
  assign n1805 = n2383 & (~PKSi_172_ | ~PKSi_85_ | n2172);
  assign n1806 = (~Pkey_172_ | n1137) & n2384;
  assign n1807_1 = n2385 & (~PKSi_179_ | ~PKSi_93_ | n2172);
  assign n1808 = (~Pkey_228_ | n1137) & n2386;
  assign n1809 = n2387 & (~\[253]  | ~PKSi_82_ | n2172);
  assign n1810 = (~Pkey_220_ | n1137) & n2388;
  assign n1811_1 = n2389 & (~PKSi_188_ | n2172 | ~N_N2741);
  assign n1812 = (~Pkey_212_ | n1137) & n2390;
  assign n1813 = n2391 & (~PKSi_176_ | ~PKSi_84_ | n2172);
  assign n1814 = (~Pkey_204_ | n1137) & n2392;
  assign n1815_1 = n2393 & (~PKSi_169_ | ~PKSi_75_ | n2172);
  assign n1816 = (~Pkey_196_ | n1137) & n2394;
  assign n1817 = n2395 & (~PKSi_185_ | n2172 | ~N_N2737);
  assign n1818 = (~Pkey_219_ | n1137) & n2396;
  assign n1819 = n2397 & (~\[333]  | ~N_N2865 | n2172);
  assign n1820 = (~Pkey_211_ | n1137) & n2398;
  assign n1821 = n2399 & (~PKSi_173_ | ~PKSi_92_ | n2172);
  assign n1822 = (~Pkey_203_ | n1137) & n2400;
  assign n1823 = n2401 & (~PKSi_183_ | ~PKSi_79_ | n2172);
  assign n1824 = (~Pkey_195_ | n1137) & n2402;
  assign n1825 = (n2059 | n2176) & (~n2175 | n2403);
  assign n1826 = (~Pkey_56_ | n1137) & n2404;
  assign n1827 = (n2060 | n2176) & (~n2175 | n2405);
  assign n1828 = (~Pkey_48_ | n1137) & n2406;
  assign n1829 = (n2061 | n2176) & (~n2175 | n2407);
  assign n1830 = (~Pkey_40_ | n1137) & n2408;
  assign n1831 = (n2062 | n2176) & (~n2175 | n2409);
  assign n1832 = (~Pkey_32_ | n1137) & n2410;
  assign n1833_1 = (n2063 | n2176) & (~n2175 | n2411);
  assign n1834 = (~Pkey_24_ | n1137) & n2412;
  assign n1835 = (n2064 | n2176) & (~n2175 | n2413);
  assign n1836 = (~Pkey_16_ | n1137) & n2414;
  assign n1837_1 = (n2065 | n2176) & (~n2175 | n2415);
  assign n1838 = (~Pkey_8_ | n1137) & n2416;
  assign n1839 = (n2066 | n2176) & (~n2175 | n2417);
  assign n1840 = (~Pkey_0_ | n1137) & n2418;
  assign n1841_1 = (n2067 | n2176) & (~n2175 | n2419);
  assign n1842 = (~Pkey_57_ | n1137) & n2420;
  assign n1843 = (n2068 | n2176) & (~n2175 | n2421);
  assign n1844 = (~Pkey_49_ | n1137) & n2422;
  assign n1845_1 = (n2069 | n2176) & (~n2175 | n2423);
  assign n1846 = (~Pkey_41_ | n1137) & n2424;
  assign n1847 = (n2070 | n2176) & (~n2175 | n2425);
  assign n1848 = (~Pkey_33_ | n1137) & n2426;
  assign n1849_1 = (n2071 | n2176) & (~n2175 | n2427);
  assign n1850 = (~Pkey_25_ | n1137) & n2428;
  assign n1851 = (n2072 | n2176) & (~n2175 | n2429);
  assign n1852 = (~Pkey_17_ | n1137) & n2430;
  assign n1853_1 = (n2073 | n2176) & (~n2175 | n2431);
  assign n1854 = (~Pkey_9_ | n1137) & n2432;
  assign n1855 = (n2074 | n2176) & (~n2175 | n2433);
  assign n1856 = (~Pkey_1_ | n1137) & n2434;
  assign n1857 = (n2075 | n2176) & (~n2175 | n2435);
  assign n1858 = (~Pkey_58_ | n1137) & n2436;
  assign n1859 = (n2076 | n2176) & (~n2175 | n2437);
  assign n1860 = (~Pkey_50_ | n1137) & n2438;
  assign n1861 = (n2077 | n2176) & (~n2175 | n2439);
  assign n1862 = (~Pkey_42_ | n1137) & n2440;
  assign n1863 = (n2078 | n2176) & (~n2175 | n2441);
  assign n1864 = (~Pkey_34_ | n1137) & n2442;
  assign n1865 = (n2079 | n2176) & (~n2175 | n2443);
  assign n1866 = (~Pkey_26_ | n1137) & n2444;
  assign n1867 = (n2080 | n2176) & (~n2175 | n2445);
  assign n1868 = (~Pkey_18_ | n1137) & n2446;
  assign n1869 = (n2081 | n2176) & (~n2175 | n2447);
  assign n1870 = (~Pkey_10_ | n1137) & n2448;
  assign n1871 = (n2082 | n2176) & (~n2175 | n2449);
  assign n1872 = (~Pkey_2_ | n1137) & n2450;
  assign n1873 = (n2083 | n2176) & (~n2175 | n2451);
  assign n1874 = (~Pkey_59_ | n1137) & n2452;
  assign n1875 = (n2084 | n2176) & (~n2175 | n2453);
  assign n1876 = (~Pkey_51_ | n1137) & n2454;
  assign n1877 = (n2085 | n2176) & (~n2175 | n2455);
  assign n1878 = (~Pkey_43_ | n1137) & n2456;
  assign n1879 = (n2086 | n2176) & (~n2175 | n2457);
  assign n1880 = (~Pkey_35_ | n1137) & n2458;
  assign n1881 = (n2087 | n2176) & (~n2175 | n2459);
  assign n1882 = (~Pkey_120_ | n1137) & n2460;
  assign n1883 = (n2088 | n2176) & (~n2175 | n2461);
  assign n1884 = (~Pkey_112_ | n1137) & n2462;
  assign n1885 = (n2089 | n2176) & (~n2175 | n2463);
  assign n1886 = (~Pkey_104_ | n1137) & n2464;
  assign n1887 = (n2090 | n2176) & (~n2175 | n2465);
  assign n1888 = (~Pkey_96_ | n1137) & n2466;
  assign n1889 = (n2091 | n2176) & (~n2175 | n2467);
  assign n1890 = (~Pkey_88_ | n1137) & n2468;
  assign n1891 = (n2092 | n2176) & (~n2175 | n2469);
  assign n1892 = (~Pkey_80_ | n1137) & n2470;
  assign n1893 = (n2093 | n2176) & (~n2175 | n2471);
  assign n1894 = (~Pkey_72_ | n1137) & n2472;
  assign n1895 = (n2094 | n2176) & (~n2175 | n2473);
  assign n1896 = (~Pkey_64_ | n1137) & n2474;
  assign n1897 = (n2095 | n2176) & (~n2175 | n2475);
  assign n1898 = (~Pkey_121_ | n1137) & n2476;
  assign n1899 = (n2096 | n2176) & (~n2175 | n2477);
  assign n1900 = (~Pkey_113_ | n1137) & n2478;
  assign n1901 = (n2097 | n2176) & (~n2175 | n2479);
  assign n1902 = (~Pkey_105_ | n1137) & n2480;
  assign n1903 = (n2098 | n2176) & (~n2175 | n2481);
  assign n1904 = (~Pkey_97_ | n1137) & n2482;
  assign n1905 = (n2099 | n2176) & (~n2175 | n2483);
  assign n1906 = (~Pkey_89_ | n1137) & n2484;
  assign n1907 = (n2100 | n2176) & (~n2175 | n2485);
  assign n1908 = (~Pkey_81_ | n1137) & n2486;
  assign n1909 = (n2101 | n2176) & (~n2175 | n2487);
  assign n1910 = (~Pkey_73_ | n1137) & n2488;
  assign n1911 = (n2102 | n2176) & (~n2175 | n2489);
  assign n1912 = (~Pkey_65_ | n1137) & n2490;
  assign n1913 = (n2103 | n2176) & (~n2175 | n2491);
  assign n1914 = (~Pkey_122_ | n1137) & n2492;
  assign n1915 = (n2104 | n2176) & (~n2175 | n2493);
  assign n1916 = (~Pkey_114_ | n1137) & n2494;
  assign n1917 = (n2105 | n2176) & (~n2175 | n2495);
  assign n1918 = (~Pkey_106_ | n1137) & n2496;
  assign n1919 = (n2106 | n2176) & (~n2175 | n2497);
  assign n1920 = (~Pkey_98_ | n1137) & n2498;
  assign n1921 = (n2107 | n2176) & (~n2175 | n2499);
  assign n1922 = (~Pkey_90_ | n1137) & n2500;
  assign n1923 = (n2108 | n2176) & (~n2175 | n2501);
  assign n1924 = (~Pkey_82_ | n1137) & n2502;
  assign n1925 = (n2109 | n2176) & (~n2175 | n2503);
  assign n1926 = (~Pkey_74_ | n1137) & n2504;
  assign n1927 = (n2110 | n2176) & (~n2175 | n2505);
  assign n1928 = (~Pkey_66_ | n1137) & n2506;
  assign n1929 = (n2111 | n2176) & (~n2175 | n2507);
  assign n1930 = (~Pkey_123_ | n1137) & n2508;
  assign n1931 = (n2112 | n2176) & (~n2175 | n2509);
  assign n1932 = (~Pkey_115_ | n1137) & n2510;
  assign n1933 = (n2113 | n2176) & (~n2175 | n2511);
  assign n1934 = (~Pkey_107_ | n1137) & n2512;
  assign n1935 = (n2114 | n2176) & (~n2175 | n2513);
  assign n1936 = (~Pkey_99_ | n1137) & n2514;
  assign n1937 = (n2115 | n2176) & (~n2175 | n2515);
  assign n1938 = (~Pkey_184_ | n1137) & n2516;
  assign n1939 = (n2116 | n2176) & (~n2175 | n2517);
  assign n1940 = (~Pkey_176_ | n1137) & n2518;
  assign n1941 = (n2117 | n2176) & (~n2175 | n2519);
  assign n1942 = (~Pkey_168_ | n1137) & n2520;
  assign n1943 = (n2118 | n2176) & (~n2175 | n2521);
  assign n1944 = (~Pkey_160_ | n1137) & n2522;
  assign n1945 = (n2119 | n2176) & (~n2175 | n2523);
  assign n1946 = (~Pkey_152_ | n1137) & n2524;
  assign n1947 = (n2120 | n2176) & (~n2175 | n2525);
  assign n1948 = (~Pkey_144_ | n1137) & n2526;
  assign n1949 = (n2121 | n2176) & (~n2175 | n2527);
  assign n1950 = (~Pkey_136_ | n1137) & n2528;
  assign n1951 = (n2122 | n2176) & (~n2175 | n2529);
  assign n1952 = (~Pkey_128_ | n1137) & n2530;
  assign n1953 = (n2123 | n2176) & (~n2175 | n2531);
  assign n1954 = (~Pkey_185_ | n1137) & n2532;
  assign n1955 = (n2124 | n2176) & (~n2175 | n2533);
  assign n1956 = (~Pkey_177_ | n1137) & n2534;
  assign n1957 = (n2125 | n2176) & (~n2175 | n2535);
  assign n1958 = (~Pkey_169_ | n1137) & n2536;
  assign n1959 = (n2126 | n2176) & (~n2175 | n2537);
  assign n1960 = (~Pkey_161_ | n1137) & n2538;
  assign n1961 = (n2127 | n2176) & (~n2175 | n2539);
  assign n1962 = (~Pkey_153_ | n1137) & n2540;
  assign n1963 = (n2128 | n2176) & (~n2175 | n2541);
  assign n1964 = (~Pkey_145_ | n1137) & n2542;
  assign n1965 = (n2129 | n2176) & (~n2175 | n2543);
  assign n1966 = (~Pkey_137_ | n1137) & n2544;
  assign n1967 = (n2130 | n2176) & (~n2175 | n2545);
  assign n1968 = (~Pkey_129_ | n1137) & n2546;
  assign n1969 = (n2131 | n2176) & (~n2175 | n2547);
  assign n1970 = (~Pkey_186_ | n1137) & n2548;
  assign n1971 = (n2132 | n2176) & (~n2175 | n2549);
  assign n1972 = (~Pkey_178_ | n1137) & n2550;
  assign n1973 = (n2133 | n2176) & (~n2175 | n2551);
  assign n1974 = (~Pkey_170_ | n1137) & n2552;
  assign n1975 = (n2134 | n2176) & (~n2175 | n2553);
  assign n1976 = (~Pkey_162_ | n1137) & n2554;
  assign n1977 = (n2135 | n2176) & (~n2175 | n2555);
  assign n1978 = (~Pkey_154_ | n1137) & n2556;
  assign n1979 = (n2136 | n2176) & (~n2175 | n2557);
  assign n1980 = (~Pkey_146_ | n1137) & n2558;
  assign n1981 = (n2137 | n2176) & (~n2175 | n2559);
  assign n1982 = (~Pkey_138_ | n1137) & n2560;
  assign n1983 = (n2138 | n2176) & (~n2175 | n2561);
  assign n1984 = (~Pkey_130_ | n1137) & n2562;
  assign n1985 = (n2139 | n2176) & (~n2175 | n2563);
  assign n1986 = (~Pkey_187_ | n1137) & n2564;
  assign n1987 = (n2140 | n2176) & (~n2175 | n2565);
  assign n1988 = (~Pkey_179_ | n1137) & n2566;
  assign n1989 = (n2141 | n2176) & (~n2175 | n2567);
  assign n1990 = (~Pkey_171_ | n1137) & n2568;
  assign n1991 = (n2142 | n2176) & (~n2175 | n2569);
  assign n1992 = (~Pkey_163_ | n1137) & n2570;
  assign n1993 = (n2143 | n2176) & (~n2175 | n2571);
  assign n1994 = (~Pkey_248_ | n1137) & n2572;
  assign n1995 = (n2144 | n2176) & (~n2175 | n2573);
  assign n1996 = (~Pkey_240_ | n1137) & n2574;
  assign n1997 = (n2145 | n2176) & (~n2175 | n2575);
  assign n1998 = (~Pkey_232_ | n1137) & n2576;
  assign n1999 = (n2146 | n2176) & (~n2175 | n2577);
  assign n2000 = (~Pkey_224_ | n1137) & n2578;
  assign n2001 = (n2147 | n2176) & (~n2175 | n2579);
  assign n2002 = (~Pkey_216_ | n1137) & n2580;
  assign n2003 = (n2148 | n2176) & (~n2175 | n2581);
  assign n2004 = (~Pkey_208_ | n1137) & n2582;
  assign n2005 = (n2149 | n2176) & (~n2175 | n2583);
  assign n2006 = (~Pkey_200_ | n1137) & n2584;
  assign n2007 = (n2150 | n2176) & (~n2175 | n2585);
  assign n2008 = (~Pkey_192_ | n1137) & n2586;
  assign n2009 = (n2151 | n2176) & (~n2175 | n2587);
  assign n2010 = (~Pkey_249_ | n1137) & n2588;
  assign n2011 = (n2152 | n2176) & (~n2175 | n2589);
  assign n2012 = (~Pkey_241_ | n1137) & n2590;
  assign n2013 = (n2153 | n2176) & (~n2175 | n2591);
  assign n2014 = (~Pkey_233_ | n1137) & n2592;
  assign n2015 = (n2154 | n2176) & (~n2175 | n2593);
  assign n2016 = (~Pkey_225_ | n1137) & n2594;
  assign n2017 = (n2155 | n2176) & (~n2175 | n2595);
  assign n2018 = (~Pkey_217_ | n1137) & n2596;
  assign n2019 = (n2156 | n2176) & (~n2175 | n2597);
  assign n2020 = (~Pkey_209_ | n1137) & n2598;
  assign n2021 = (n2157 | n2176) & (~n2175 | n2599);
  assign n2022 = (~Pkey_201_ | n1137) & n2600;
  assign n2023 = (n2158 | n2176) & (~n2175 | n2601);
  assign n2024 = (~Pkey_193_ | n1137) & n2602;
  assign n2025 = (n2159 | n2176) & (~n2175 | n2603);
  assign n2026 = (~Pkey_250_ | n1137) & n2604;
  assign n2027 = (n2160 | n2176) & (~n2175 | n2605);
  assign n2028 = (~Pkey_242_ | n1137) & n2606;
  assign n2029 = (n2161 | n2176) & (~n2175 | n2607);
  assign n2030 = (~Pkey_234_ | n1137) & n2608;
  assign n2031 = (n2162 | n2176) & (~n2175 | n2609);
  assign n2032 = (~Pkey_226_ | n1137) & n2610;
  assign n2033 = (n2163 | n2176) & (~n2175 | n2611);
  assign n2034 = (~Pkey_218_ | n1137) & n2612;
  assign n2035 = (n2164 | n2176) & (~n2175 | n2613);
  assign n2036 = (~Pkey_210_ | n1137) & n2614;
  assign n2037 = (n2165 | n2176) & (~n2175 | n2615);
  assign n2038 = (~Pkey_202_ | n1137) & n2616;
  assign n2039 = (n2166 | n2176) & (~n2175 | n2617);
  assign n2040 = (~Pkey_194_ | n1137) & n2618;
  assign n2041 = (n2167 | n2176) & (~n2175 | n2619);
  assign n2042 = (~Pkey_251_ | n1137) & n2620;
  assign n2043 = (n2168 | n2176) & (~n2175 | n2621);
  assign n2044 = (~Pkey_243_ | n1137) & n2622;
  assign n2045 = (n2169 | n2176) & (~n2175 | n2623);
  assign n2046 = (~Pkey_235_ | n1137) & n2624;
  assign n2047 = (n2170 | n2176) & (~n2175 | n2625);
  assign n2048 = (~Pkey_227_ | n1137) & n2626;
  assign n2049 = ~Pcount_3_ | n1596 | n2177;
  assign n2050 = n1595 | Pcount_3_ | Pencrypt_0_;
  assign n2051 = (n2739 & (~Pcount_1_ | n2740)) | (Pcount_1_ & n2740);
  assign n2052 = Pencrypt_0_ | ~Pcount_1_;
  assign n2053 = Pcount_2_ & (~n2052 | ~n2740);
  assign n2054 = n1137 & (Pstart_0_ | ~Pcount_0_ | ~n2178);
  assign n2055 = ~Pcount_2_ & ~Pcount_0_;
  assign n2056 = (~Pencrypt_0_ | n1599) & n2050;
  assign n2057 = (~n1596 & (Pencrypt_0_ | n2055)) | (~Pencrypt_0_ & n2055);
  assign n2058 = n2056 & (~Pcount_3_ | (n2052 & n2057));
  assign n2059 = ~PKSi_118_ ^ PKSi_4_;
  assign n2060 = ~PKSi_102_ ^ PKSi_23_;
  assign n2061 = ~PKSi_98_ ^ PKSi_6_;
  assign n2062 = ~PKSi_119_ ^ PKSi_15_;
  assign n2063 = ~PKSi_106_ ^ PKSi_5_;
  assign n2064 = ~PKSi_112_ ^ PKSi_9_;
  assign n2065 = ~PKSi_19_ ^ N_N2986;
  assign n2066 = ~PKSi_117_ ^ PKSi_17_;
  assign n2067 = ~PKSi_99_ ^ N_N2853;
  assign n2068 = ~PKSi_11_ ^ N_N2982;
  assign n2069 = ~PKSi_110_ ^ PKSi_2_;
  assign n2070 = ~PKSi_103_ ^ PKSi_14_;
  assign n2071 = ~PKSi_96_ ^ PKSi_22_;
  assign n2072 = ~PKSi_115_ ^ PKSi_0_;
  assign n2073 = ~PKSi_8_ ^ N_N2976;
  assign n2074 = ~PKSi_108_ ^ PKSi_18_;
  assign n2075 = ~PKSi_105_ ^ PKSi_1_;
  assign n2076 = ~PKSi_114_ ^ N_N2843;
  assign n2077 = ~PKSi_100_ ^ PKSi_13_;
  assign n2078 = ~PKSi_107_ ^ PKSi_21_;
  assign n2079 = ~PKSi_109_ ^ PKSi_10_;
  assign n2080 = ~PKSi_116_ ^ N_N2838;
  assign n2081 = ~PKSi_104_ ^ PKSi_12_;
  assign n2082 = ~PKSi_97_ ^ PKSi_3_;
  assign n2083 = ~PKSi_113_ ^ N_N2834;
  assign n2084 = ~PKSi_16_ ^ N_N2964;
  assign n2085 = ~PKSi_101_ ^ PKSi_20_;
  assign n2086 = ~PKSi_111_ ^ PKSi_7_;
  assign n2087 = ~PKSi_142_ ^ PKSi_28_;
  assign n2088 = ~PKSi_126_ ^ PKSi_47_;
  assign n2089 = ~PKSi_122_ ^ PKSi_30_;
  assign n2090 = ~\[282]  ^ PKSi_39_;
  assign n2091 = ~PKSi_130_ ^ PKSi_29_;
  assign n2092 = ~PKSi_136_ ^ PKSi_33_;
  assign n2093 = ~PKSi_43_ ^ N_N2954;
  assign n2094 = ~PKSi_141_ ^ PKSi_41_;
  assign n2095 = ~PKSi_123_ ^ N_N2821;
  assign n2096 = ~PKSi_35_ ^ N_N2950;
  assign n2097 = ~PKSi_134_ ^ PKSi_26_;
  assign n2098 = ~PKSi_127_ ^ PKSi_38_;
  assign n2099 = ~PKSi_120_ ^ PKSi_46_;
  assign n2100 = ~PKSi_24_ ^ N_N2945;
  assign n2101 = ~PKSi_32_ ^ N_N2943;
  assign n2102 = ~PKSi_132_ ^ PKSi_42_;
  assign n2103 = ~PKSi_129_ ^ PKSi_25_;
  assign n2104 = ~PKSi_138_ ^ N_N2811;
  assign n2105 = ~PKSi_124_ ^ PKSi_37_;
  assign n2106 = ~PKSi_131_ ^ PKSi_45_;
  assign n2107 = ~PKSi_133_ ^ PKSi_34_;
  assign n2108 = ~PKSi_140_ ^ N_N2806;
  assign n2109 = ~PKSi_128_ ^ PKSi_36_;
  assign n2110 = ~PKSi_121_ ^ PKSi_27_;
  assign n2111 = ~PKSi_137_ ^ N_N2802;
  assign n2112 = ~PKSi_40_ ^ N_N2931;
  assign n2113 = ~PKSi_125_ ^ PKSi_44_;
  assign n2114 = ~PKSi_135_ ^ PKSi_31_;
  assign n2115 = ~PKSi_166_ ^ PKSi_52_;
  assign n2116 = ~PKSi_150_ ^ PKSi_71_;
  assign n2117 = ~PKSi_146_ ^ PKSi_54_;
  assign n2118 = ~PKSi_167_ ^ PKSi_63_;
  assign n2119 = ~PKSi_154_ ^ PKSi_53_;
  assign n2120 = ~PKSi_160_ ^ PKSi_57_;
  assign n2121 = ~PKSi_67_ ^ N_N2921;
  assign n2122 = ~PKSi_165_ ^ PKSi_65_;
  assign n2123 = ~PKSi_147_ ^ N_N2789;
  assign n2124 = ~PKSi_59_ ^ N_N2917;
  assign n2125 = ~PKSi_158_ ^ PKSi_50_;
  assign n2126 = ~PKSi_151_ ^ PKSi_62_;
  assign n2127 = ~PKSi_144_ ^ PKSi_70_;
  assign n2128 = ~PKSi_163_ ^ PKSi_48_;
  assign n2129 = ~PKSi_153_ ^ PKSi_56_;
  assign n2130 = ~PKSi_156_ ^ PKSi_66_;
  assign n2131 = ~PKSi_49_ ^ N_N2909;
  assign n2132 = ~PKSi_162_ ^ N_N2779;
  assign n2133 = ~PKSi_148_ ^ PKSi_61_;
  assign n2134 = ~PKSi_155_ ^ PKSi_69_;
  assign n2135 = ~PKSi_157_ ^ PKSi_58_;
  assign n2136 = ~PKSi_164_ ^ N_N2774;
  assign n2137 = ~PKSi_152_ ^ PKSi_60_;
  assign n2138 = ~PKSi_145_ ^ PKSi_51_;
  assign n2139 = ~PKSi_161_ ^ N_N2770;
  assign n2140 = ~PKSi_64_ ^ N_N2899;
  assign n2141 = ~PKSi_149_ ^ PKSi_68_;
  assign n2142 = ~PKSi_159_ ^ PKSi_55_;
  assign n2143 = ~PKSi_190_ ^ PKSi_76_;
  assign n2144 = ~PKSi_174_ ^ PKSi_95_;
  assign n2145 = ~PKSi_170_ ^ PKSi_78_;
  assign n2146 = ~\[234]  ^ PKSi_87_;
  assign n2147 = ~PKSi_178_ ^ PKSi_77_;
  assign n2148 = ~PKSi_184_ ^ PKSi_81_;
  assign n2149 = ~PKSi_91_ ^ N_N2889;
  assign n2150 = ~PKSi_189_ ^ PKSi_89_;
  assign n2151 = ~PKSi_171_ ^ N_N2757;
  assign n2152 = ~PKSi_83_ ^ N_N2885;
  assign n2153 = ~PKSi_182_ ^ PKSi_74_;
  assign n2154 = ~PKSi_175_ ^ PKSi_86_;
  assign n2155 = ~PKSi_94_ ^ N_N2881;
  assign n2156 = ~PKSi_72_ ^ N_N2879;
  assign n2157 = ~PKSi_80_ ^ N_N2877;
  assign n2158 = ~PKSi_180_ ^ N_N2749;
  assign n2159 = ~PKSi_177_ ^ PKSi_73_;
  assign n2160 = ~PKSi_186_ ^ N_N2746;
  assign n2161 = ~PKSi_172_ ^ PKSi_85_;
  assign n2162 = ~PKSi_179_ ^ PKSi_93_;
  assign n2163 = ~\[253]  ^ PKSi_82_;
  assign n2164 = ~PKSi_188_ ^ N_N2741;
  assign n2165 = ~PKSi_176_ ^ PKSi_84_;
  assign n2166 = ~PKSi_169_ ^ PKSi_75_;
  assign n2167 = ~PKSi_185_ ^ N_N2737;
  assign n2168 = ~\[333]  ^ N_N2865;
  assign n2169 = ~PKSi_173_ ^ PKSi_92_;
  assign n2170 = ~PKSi_183_ ^ PKSi_79_;
  assign n2171 = Pencrypt_0_ & ~n1600;
  assign n2172 = Pstart_0_ | n2171;
  assign n2173 = Pstart_0_ | ~n2171;
  assign n2174 = ~Pencrypt_0_ | ~n1600;
  assign n2175 = ~Pstart_0_ & n2174;
  assign n2176 = Pstart_0_ | n2174;
  assign n2177 = Pstart_0_ | ~Pencrypt_0_;
  assign n2178 = n2741 & ((Pencrypt_0_ & ~Pcount_2_) | ~Pcount_1_);
  assign n2179 = n2059 | n2173;
  assign n2180 = (~n1140 & ~n2627) | (n1139_1 & (~n1140 | n2627));
  assign n2181 = n2060 | n2173;
  assign n2182 = (~n1140 & ~n2628) | (n1139_1 & (~n1140 | n2628));
  assign n2183 = n2061 | n2173;
  assign n2184 = (~n1140 & ~n2629) | (n1139_1 & (~n1140 | n2629));
  assign n2185 = n2062 | n2173;
  assign n2186 = (~n1140 & ~n2630) | (n1139_1 & (~n1140 | n2630));
  assign n2187 = n2063 | n2173;
  assign n2188 = (~n1140 & ~n2631) | (n1139_1 & (~n1140 | n2631));
  assign n2189 = n2064 | n2173;
  assign n2190 = (~n1140 & ~n2632) | (n1139_1 & (~n1140 | n2632));
  assign n2191 = n2065 | n2173;
  assign n2192 = (~n1140 & ~n2633) | (n1139_1 & (~n1140 | n2633));
  assign n2193 = n2066 | n2173;
  assign n2194 = (~n1140 & ~n2634) | (n1139_1 & (~n1140 | n2634));
  assign n2195 = n2067 | n2173;
  assign n2196 = (~n1140 & ~n2635) | (n1139_1 & (~n1140 | n2635));
  assign n2197 = n2068 | n2173;
  assign n2198 = (~n1140 & ~n2636) | (n1139_1 & (~n1140 | n2636));
  assign n2199 = n2069 | n2173;
  assign n2200 = (~n1140 & ~n2637) | (n1139_1 & (~n1140 | n2637));
  assign n2201 = n2070 | n2173;
  assign n2202 = (~n1140 & ~n2638) | (n1139_1 & (~n1140 | n2638));
  assign n2203 = n2071 | n2173;
  assign n2204 = (~n1140 & ~n2639) | (n1139_1 & (~n1140 | n2639));
  assign n2205 = n2072 | n2173;
  assign n2206 = (~n1140 & ~n2640) | (n1139_1 & (~n1140 | n2640));
  assign n2207 = n2073 | n2173;
  assign n2208 = (~n1140 & ~n2641) | (n1139_1 & (~n1140 | n2641));
  assign n2209 = n2074 | n2173;
  assign n2210 = (~n1140 & ~n2642) | (n1139_1 & (~n1140 | n2642));
  assign n2211 = n2075 | n2173;
  assign n2212 = (~n1140 & ~n2643) | (n1139_1 & (~n1140 | n2643));
  assign n2213 = n2076 | n2173;
  assign n2214 = (~n1140 & ~n2644) | (n1139_1 & (~n1140 | n2644));
  assign n2215 = n2077 | n2173;
  assign n2216 = (~n1140 & ~n2645) | (n1139_1 & (~n1140 | n2645));
  assign n2217 = n2078 | n2173;
  assign n2218 = (~n1140 & ~n2646) | (n1139_1 & (~n1140 | n2646));
  assign n2219 = n2079 | n2173;
  assign n2220 = (~n1140 & ~n2647) | (n1139_1 & (~n1140 | n2647));
  assign n2221 = n2080 | n2173;
  assign n2222 = (~n1140 & ~n2648) | (n1139_1 & (~n1140 | n2648));
  assign n2223 = n2081 | n2173;
  assign n2224 = (~n1140 & ~n2649) | (n1139_1 & (~n1140 | n2649));
  assign n2225 = n2082 | n2173;
  assign n2226 = (~n1140 & ~n2650) | (n1139_1 & (~n1140 | n2650));
  assign n2227 = n2083 | n2173;
  assign n2228 = (~n1140 & ~n2651) | (n1139_1 & (~n1140 | n2651));
  assign n2229 = n2084 | n2173;
  assign n2230 = (~n1140 & ~n2652) | (n1139_1 & (~n1140 | n2652));
  assign n2231 = n2085 | n2173;
  assign n2232 = (~n1140 & ~n2653) | (n1139_1 & (~n1140 | n2653));
  assign n2233 = n2086 | n2173;
  assign n2234 = (~n1140 & ~n2654) | (n1139_1 & (~n1140 | n2654));
  assign n2235 = n2087 | n2173;
  assign n2236 = (~n1140 & ~n2655) | (n1139_1 & (~n1140 | n2655));
  assign n2237 = n2088 | n2173;
  assign n2238 = (~n1140 & ~n2656) | (n1139_1 & (~n1140 | n2656));
  assign n2239 = n2089 | n2173;
  assign n2240 = (~n1140 & ~n2657) | (n1139_1 & (~n1140 | n2657));
  assign n2241 = n2090 | n2173;
  assign n2242 = (~n1140 & ~n2658) | (n1139_1 & (~n1140 | n2658));
  assign n2243 = n2091 | n2173;
  assign n2244 = (~n1140 & ~n2659) | (n1139_1 & (~n1140 | n2659));
  assign n2245 = n2092 | n2173;
  assign n2246 = (~n1140 & ~n2660) | (n1139_1 & (~n1140 | n2660));
  assign n2247 = n2093 | n2173;
  assign n2248 = (~n1140 & ~n2661) | (n1139_1 & (~n1140 | n2661));
  assign n2249 = n2094 | n2173;
  assign n2250 = (~n1140 & ~n2662) | (n1139_1 & (~n1140 | n2662));
  assign n2251 = n2095 | n2173;
  assign n2252 = (~n1140 & ~n2663) | (n1139_1 & (~n1140 | n2663));
  assign n2253 = n2096 | n2173;
  assign n2254 = (~n1140 & ~n2664) | (n1139_1 & (~n1140 | n2664));
  assign n2255 = n2097 | n2173;
  assign n2256 = (~n1140 & ~n2665) | (n1139_1 & (~n1140 | n2665));
  assign n2257 = n2098 | n2173;
  assign n2258 = (~n1140 & ~n2666) | (n1139_1 & (~n1140 | n2666));
  assign n2259 = n2099 | n2173;
  assign n2260 = (~n1140 & ~n2667) | (n1139_1 & (~n1140 | n2667));
  assign n2261 = n2100 | n2173;
  assign n2262 = (~n1140 & ~n2668) | (n1139_1 & (~n1140 | n2668));
  assign n2263 = n2101 | n2173;
  assign n2264 = (~n1140 & ~n2669) | (n1139_1 & (~n1140 | n2669));
  assign n2265 = n2102 | n2173;
  assign n2266 = (~n1140 & ~n2670) | (n1139_1 & (~n1140 | n2670));
  assign n2267 = n2103 | n2173;
  assign n2268 = (~n1140 & ~n2671) | (n1139_1 & (~n1140 | n2671));
  assign n2269 = n2104 | n2173;
  assign n2270 = (~n1140 & ~n2672) | (n1139_1 & (~n1140 | n2672));
  assign n2271 = n2105 | n2173;
  assign n2272 = (~n1140 & ~n2673) | (n1139_1 & (~n1140 | n2673));
  assign n2273 = n2106 | n2173;
  assign n2274 = (~n1140 & ~n2674) | (n1139_1 & (~n1140 | n2674));
  assign n2275 = n2107 | n2173;
  assign n2276 = (~n1140 & ~n2675) | (n1139_1 & (~n1140 | n2675));
  assign n2277 = n2108 | n2173;
  assign n2278 = (~n1140 & ~n2676) | (n1139_1 & (~n1140 | n2676));
  assign n2279 = n2109 | n2173;
  assign n2280 = (~n1140 & ~n2677) | (n1139_1 & (~n1140 | n2677));
  assign n2281 = n2110 | n2173;
  assign n2282 = (~n1140 & ~n2678) | (n1139_1 & (~n1140 | n2678));
  assign n2283 = n2111 | n2173;
  assign n2284 = (~n1140 & ~n2679) | (n1139_1 & (~n1140 | n2679));
  assign n2285 = n2112 | n2173;
  assign n2286 = (~n1140 & ~n2680) | (n1139_1 & (~n1140 | n2680));
  assign n2287 = n2113 | n2173;
  assign n2288 = (~n1140 & ~n2681) | (n1139_1 & (~n1140 | n2681));
  assign n2289 = n2114 | n2173;
  assign n2290 = (~n1140 & ~n2682) | (n1139_1 & (~n1140 | n2682));
  assign n2291 = n2115 | n2173;
  assign n2292 = (~n1140 & ~n2683) | (n1139_1 & (~n1140 | n2683));
  assign n2293 = n2116 | n2173;
  assign n2294 = (~n1140 & ~n2684) | (n1139_1 & (~n1140 | n2684));
  assign n2295 = n2117 | n2173;
  assign n2296 = (~n1140 & ~n2685) | (n1139_1 & (~n1140 | n2685));
  assign n2297 = n2118 | n2173;
  assign n2298 = (~n1140 & ~n2686) | (n1139_1 & (~n1140 | n2686));
  assign n2299 = n2119 | n2173;
  assign n2300 = (~n1140 & ~n2687) | (n1139_1 & (~n1140 | n2687));
  assign n2301 = n2120 | n2173;
  assign n2302 = (~n1140 & ~n2688) | (n1139_1 & (~n1140 | n2688));
  assign n2303 = n2121 | n2173;
  assign n2304 = (~n1140 & ~n2689) | (n1139_1 & (~n1140 | n2689));
  assign n2305 = n2122 | n2173;
  assign n2306 = (~n1140 & ~n2690) | (n1139_1 & (~n1140 | n2690));
  assign n2307 = n2123 | n2173;
  assign n2308 = (~n1140 & ~n2691) | (n1139_1 & (~n1140 | n2691));
  assign n2309 = n2124 | n2173;
  assign n2310 = (~n1140 & ~n2692) | (n1139_1 & (~n1140 | n2692));
  assign n2311 = n2125 | n2173;
  assign n2312 = (~n1140 & ~n2693) | (n1139_1 & (~n1140 | n2693));
  assign n2313 = n2126 | n2173;
  assign n2314 = (~n1140 & ~n2694) | (n1139_1 & (~n1140 | n2694));
  assign n2315 = n2127 | n2173;
  assign n2316 = (~n1140 & ~n2695) | (n1139_1 & (~n1140 | n2695));
  assign n2317 = n2128 | n2173;
  assign n2318 = (~n1140 & ~n2696) | (n1139_1 & (~n1140 | n2696));
  assign n2319 = n2129 | n2173;
  assign n2320 = (~n1140 & ~n2697) | (n1139_1 & (~n1140 | n2697));
  assign n2321 = n2130 | n2173;
  assign n2322 = (~n1140 & ~n2698) | (n1139_1 & (~n1140 | n2698));
  assign n2323 = n2131 | n2173;
  assign n2324 = (~n1140 & ~n2699) | (n1139_1 & (~n1140 | n2699));
  assign n2325 = n2132 | n2173;
  assign n2326 = (~n1140 & ~n2700) | (n1139_1 & (~n1140 | n2700));
  assign n2327 = n2133 | n2173;
  assign n2328 = (~n1140 & ~n2701) | (n1139_1 & (~n1140 | n2701));
  assign n2329 = n2134 | n2173;
  assign n2330 = (~n1140 & ~n2702) | (n1139_1 & (~n1140 | n2702));
  assign n2331 = n2135 | n2173;
  assign n2332 = (~n1140 & ~n2703) | (n1139_1 & (~n1140 | n2703));
  assign n2333 = n2136 | n2173;
  assign n2334 = (~n1140 & ~n2704) | (n1139_1 & (~n1140 | n2704));
  assign n2335 = n2137 | n2173;
  assign n2336 = (~n1140 & ~n2705) | (n1139_1 & (~n1140 | n2705));
  assign n2337 = n2138 | n2173;
  assign n2338 = (~n1140 & ~n2706) | (n1139_1 & (~n1140 | n2706));
  assign n2339 = n2139 | n2173;
  assign n2340 = (~n1140 & ~n2707) | (n1139_1 & (~n1140 | n2707));
  assign n2341 = n2140 | n2173;
  assign n2342 = (~n1140 & ~n2708) | (n1139_1 & (~n1140 | n2708));
  assign n2343 = n2141 | n2173;
  assign n2344 = (~n1140 & ~n2709) | (n1139_1 & (~n1140 | n2709));
  assign n2345 = n2142 | n2173;
  assign n2346 = (~n1140 & ~n2710) | (n1139_1 & (~n1140 | n2710));
  assign n2347 = n2143 | n2173;
  assign n2348 = (~n1140 & ~n2711) | (n1139_1 & (~n1140 | n2711));
  assign n2349 = n2144 | n2173;
  assign n2350 = (~n1140 & ~n2712) | (n1139_1 & (~n1140 | n2712));
  assign n2351 = n2145 | n2173;
  assign n2352 = (~n1140 & ~n2713) | (n1139_1 & (~n1140 | n2713));
  assign n2353 = n2146 | n2173;
  assign n2354 = (~n1140 & ~n2714) | (n1139_1 & (~n1140 | n2714));
  assign n2355 = n2147 | n2173;
  assign n2356 = (~n1140 & ~n2715) | (n1139_1 & (~n1140 | n2715));
  assign n2357 = n2148 | n2173;
  assign n2358 = (~n1140 & ~n2716) | (n1139_1 & (~n1140 | n2716));
  assign n2359 = n2149 | n2173;
  assign n2360 = (~n1140 & ~n2717) | (n1139_1 & (~n1140 | n2717));
  assign n2361 = n2150 | n2173;
  assign n2362 = (~n1140 & ~n2718) | (n1139_1 & (~n1140 | n2718));
  assign n2363 = n2151 | n2173;
  assign n2364 = (~n1140 & ~n2719) | (n1139_1 & (~n1140 | n2719));
  assign n2365 = n2152 | n2173;
  assign n2366 = (~n1140 & ~n2720) | (n1139_1 & (~n1140 | n2720));
  assign n2367 = n2153 | n2173;
  assign n2368 = (~n1140 & ~n2721) | (n1139_1 & (~n1140 | n2721));
  assign n2369 = n2154 | n2173;
  assign n2370 = (~n1140 & ~n2722) | (n1139_1 & (~n1140 | n2722));
  assign n2371 = n2155 | n2173;
  assign n2372 = (~n1140 & ~n2723) | (n1139_1 & (~n1140 | n2723));
  assign n2373 = n2156 | n2173;
  assign n2374 = (~n1140 & ~n2724) | (n1139_1 & (~n1140 | n2724));
  assign n2375 = n2157 | n2173;
  assign n2376 = (~n1140 & ~n2725) | (n1139_1 & (~n1140 | n2725));
  assign n2377 = n2158 | n2173;
  assign n2378 = (~n1140 & ~n2726) | (n1139_1 & (~n1140 | n2726));
  assign n2379 = n2159 | n2173;
  assign n2380 = (~n1140 & ~n2727) | (n1139_1 & (~n1140 | n2727));
  assign n2381 = n2160 | n2173;
  assign n2382 = (~n1140 & ~n2728) | (n1139_1 & (~n1140 | n2728));
  assign n2383 = n2161 | n2173;
  assign n2384 = (~n1140 & ~n2729) | (n1139_1 & (~n1140 | n2729));
  assign n2385 = n2162 | n2173;
  assign n2386 = (~n1140 & ~n2730) | (n1139_1 & (~n1140 | n2730));
  assign n2387 = n2163 | n2173;
  assign n2388 = (~n1140 & ~n2731) | (n1139_1 & (~n1140 | n2731));
  assign n2389 = n2164 | n2173;
  assign n2390 = (~n1140 & ~n2732) | (n1139_1 & (~n1140 | n2732));
  assign n2391 = n2165 | n2173;
  assign n2392 = (~n1140 & ~n2733) | (n1139_1 & (~n1140 | n2733));
  assign n2393 = n2166 | n2173;
  assign n2394 = (~n1140 & ~n2734) | (n1139_1 & (~n1140 | n2734));
  assign n2395 = n2167 | n2173;
  assign n2396 = (~n1140 & ~n2735) | (n1139_1 & (~n1140 | n2735));
  assign n2397 = n2168 | n2173;
  assign n2398 = (~n1140 & ~n2736) | (n1139_1 & (~n1140 | n2736));
  assign n2399 = n2169 | n2173;
  assign n2400 = (~n1140 & ~n2737) | (n1139_1 & (~n1140 | n2737));
  assign n2401 = n2170 | n2173;
  assign n2402 = (~n1140 & ~n2738) | (n1139_1 & (~n1140 | n2738));
  assign n2403 = ~PKSi_118_ | ~PKSi_4_;
  assign n2404 = (~n1140 & n2627) | (n1139_1 & (~n1140 | ~n2627));
  assign n2405 = ~PKSi_102_ | ~PKSi_23_;
  assign n2406 = (~n1140 & n2628) | (n1139_1 & (~n1140 | ~n2628));
  assign n2407 = ~PKSi_98_ | ~PKSi_6_;
  assign n2408 = (~n1140 & n2629) | (n1139_1 & (~n1140 | ~n2629));
  assign n2409 = ~PKSi_119_ | ~PKSi_15_;
  assign n2410 = (~n1140 & n2630) | (n1139_1 & (~n1140 | ~n2630));
  assign n2411 = ~PKSi_106_ | ~PKSi_5_;
  assign n2412 = (~n1140 & n2631) | (n1139_1 & (~n1140 | ~n2631));
  assign n2413 = ~PKSi_112_ | ~PKSi_9_;
  assign n2414 = (~n1140 & n2632) | (n1139_1 & (~n1140 | ~n2632));
  assign n2415 = ~PKSi_19_ | ~N_N2986;
  assign n2416 = (~n1140 & n2633) | (n1139_1 & (~n1140 | ~n2633));
  assign n2417 = ~PKSi_117_ | ~PKSi_17_;
  assign n2418 = (~n1140 & n2634) | (n1139_1 & (~n1140 | ~n2634));
  assign n2419 = ~PKSi_99_ | ~N_N2853;
  assign n2420 = (~n1140 & n2635) | (n1139_1 & (~n1140 | ~n2635));
  assign n2421 = ~PKSi_11_ | ~N_N2982;
  assign n2422 = (~n1140 & n2636) | (n1139_1 & (~n1140 | ~n2636));
  assign n2423 = ~PKSi_110_ | ~PKSi_2_;
  assign n2424 = (~n1140 & n2637) | (n1139_1 & (~n1140 | ~n2637));
  assign n2425 = ~PKSi_103_ | ~PKSi_14_;
  assign n2426 = (~n1140 & n2638) | (n1139_1 & (~n1140 | ~n2638));
  assign n2427 = ~PKSi_96_ | ~PKSi_22_;
  assign n2428 = (~n1140 & n2639) | (n1139_1 & (~n1140 | ~n2639));
  assign n2429 = ~PKSi_115_ | ~PKSi_0_;
  assign n2430 = (~n1140 & n2640) | (n1139_1 & (~n1140 | ~n2640));
  assign n2431 = ~PKSi_8_ | ~N_N2976;
  assign n2432 = (~n1140 & n2641) | (n1139_1 & (~n1140 | ~n2641));
  assign n2433 = ~PKSi_108_ | ~PKSi_18_;
  assign n2434 = (~n1140 & n2642) | (n1139_1 & (~n1140 | ~n2642));
  assign n2435 = ~PKSi_105_ | ~PKSi_1_;
  assign n2436 = (~n1140 & n2643) | (n1139_1 & (~n1140 | ~n2643));
  assign n2437 = ~PKSi_114_ | ~N_N2843;
  assign n2438 = (~n1140 & n2644) | (n1139_1 & (~n1140 | ~n2644));
  assign n2439 = ~PKSi_100_ | ~PKSi_13_;
  assign n2440 = (~n1140 & n2645) | (n1139_1 & (~n1140 | ~n2645));
  assign n2441 = ~PKSi_107_ | ~PKSi_21_;
  assign n2442 = (~n1140 & n2646) | (n1139_1 & (~n1140 | ~n2646));
  assign n2443 = ~PKSi_109_ | ~PKSi_10_;
  assign n2444 = (~n1140 & n2647) | (n1139_1 & (~n1140 | ~n2647));
  assign n2445 = ~PKSi_116_ | ~N_N2838;
  assign n2446 = (~n1140 & n2648) | (n1139_1 & (~n1140 | ~n2648));
  assign n2447 = ~PKSi_104_ | ~PKSi_12_;
  assign n2448 = (~n1140 & n2649) | (n1139_1 & (~n1140 | ~n2649));
  assign n2449 = ~PKSi_97_ | ~PKSi_3_;
  assign n2450 = (~n1140 & n2650) | (n1139_1 & (~n1140 | ~n2650));
  assign n2451 = ~PKSi_113_ | ~N_N2834;
  assign n2452 = (~n1140 & n2651) | (n1139_1 & (~n1140 | ~n2651));
  assign n2453 = ~PKSi_16_ | ~N_N2964;
  assign n2454 = (~n1140 & n2652) | (n1139_1 & (~n1140 | ~n2652));
  assign n2455 = ~PKSi_101_ | ~PKSi_20_;
  assign n2456 = (~n1140 & n2653) | (n1139_1 & (~n1140 | ~n2653));
  assign n2457 = ~PKSi_111_ | ~PKSi_7_;
  assign n2458 = (~n1140 & n2654) | (n1139_1 & (~n1140 | ~n2654));
  assign n2459 = ~PKSi_142_ | ~PKSi_28_;
  assign n2460 = (~n1140 & n2655) | (n1139_1 & (~n1140 | ~n2655));
  assign n2461 = ~PKSi_126_ | ~PKSi_47_;
  assign n2462 = (~n1140 & n2656) | (n1139_1 & (~n1140 | ~n2656));
  assign n2463 = ~PKSi_122_ | ~PKSi_30_;
  assign n2464 = (~n1140 & n2657) | (n1139_1 & (~n1140 | ~n2657));
  assign n2465 = ~\[282]  | ~PKSi_39_;
  assign n2466 = (~n1140 & n2658) | (n1139_1 & (~n1140 | ~n2658));
  assign n2467 = ~PKSi_130_ | ~PKSi_29_;
  assign n2468 = (~n1140 & n2659) | (n1139_1 & (~n1140 | ~n2659));
  assign n2469 = ~PKSi_136_ | ~PKSi_33_;
  assign n2470 = (~n1140 & n2660) | (n1139_1 & (~n1140 | ~n2660));
  assign n2471 = ~PKSi_43_ | ~N_N2954;
  assign n2472 = (~n1140 & n2661) | (n1139_1 & (~n1140 | ~n2661));
  assign n2473 = ~PKSi_141_ | ~PKSi_41_;
  assign n2474 = (~n1140 & n2662) | (n1139_1 & (~n1140 | ~n2662));
  assign n2475 = ~PKSi_123_ | ~N_N2821;
  assign n2476 = (~n1140 & n2663) | (n1139_1 & (~n1140 | ~n2663));
  assign n2477 = ~PKSi_35_ | ~N_N2950;
  assign n2478 = (~n1140 & n2664) | (n1139_1 & (~n1140 | ~n2664));
  assign n2479 = ~PKSi_134_ | ~PKSi_26_;
  assign n2480 = (~n1140 & n2665) | (n1139_1 & (~n1140 | ~n2665));
  assign n2481 = ~PKSi_127_ | ~PKSi_38_;
  assign n2482 = (~n1140 & n2666) | (n1139_1 & (~n1140 | ~n2666));
  assign n2483 = ~PKSi_120_ | ~PKSi_46_;
  assign n2484 = (~n1140 & n2667) | (n1139_1 & (~n1140 | ~n2667));
  assign n2485 = ~PKSi_24_ | ~N_N2945;
  assign n2486 = (~n1140 & n2668) | (n1139_1 & (~n1140 | ~n2668));
  assign n2487 = ~PKSi_32_ | ~N_N2943;
  assign n2488 = (~n1140 & n2669) | (n1139_1 & (~n1140 | ~n2669));
  assign n2489 = ~PKSi_132_ | ~PKSi_42_;
  assign n2490 = (~n1140 & n2670) | (n1139_1 & (~n1140 | ~n2670));
  assign n2491 = ~PKSi_129_ | ~PKSi_25_;
  assign n2492 = (~n1140 & n2671) | (n1139_1 & (~n1140 | ~n2671));
  assign n2493 = ~PKSi_138_ | ~N_N2811;
  assign n2494 = (~n1140 & n2672) | (n1139_1 & (~n1140 | ~n2672));
  assign n2495 = ~PKSi_124_ | ~PKSi_37_;
  assign n2496 = (~n1140 & n2673) | (n1139_1 & (~n1140 | ~n2673));
  assign n2497 = ~PKSi_131_ | ~PKSi_45_;
  assign n2498 = (~n1140 & n2674) | (n1139_1 & (~n1140 | ~n2674));
  assign n2499 = ~PKSi_133_ | ~PKSi_34_;
  assign n2500 = (~n1140 & n2675) | (n1139_1 & (~n1140 | ~n2675));
  assign n2501 = ~PKSi_140_ | ~N_N2806;
  assign n2502 = (~n1140 & n2676) | (n1139_1 & (~n1140 | ~n2676));
  assign n2503 = ~PKSi_128_ | ~PKSi_36_;
  assign n2504 = (~n1140 & n2677) | (n1139_1 & (~n1140 | ~n2677));
  assign n2505 = ~PKSi_121_ | ~PKSi_27_;
  assign n2506 = (~n1140 & n2678) | (n1139_1 & (~n1140 | ~n2678));
  assign n2507 = ~PKSi_137_ | ~N_N2802;
  assign n2508 = (~n1140 & n2679) | (n1139_1 & (~n1140 | ~n2679));
  assign n2509 = ~PKSi_40_ | ~N_N2931;
  assign n2510 = (~n1140 & n2680) | (n1139_1 & (~n1140 | ~n2680));
  assign n2511 = ~PKSi_125_ | ~PKSi_44_;
  assign n2512 = (~n1140 & n2681) | (n1139_1 & (~n1140 | ~n2681));
  assign n2513 = ~PKSi_135_ | ~PKSi_31_;
  assign n2514 = (~n1140 & n2682) | (n1139_1 & (~n1140 | ~n2682));
  assign n2515 = ~PKSi_166_ | ~PKSi_52_;
  assign n2516 = (~n1140 & n2683) | (n1139_1 & (~n1140 | ~n2683));
  assign n2517 = ~PKSi_150_ | ~PKSi_71_;
  assign n2518 = (~n1140 & n2684) | (n1139_1 & (~n1140 | ~n2684));
  assign n2519 = ~PKSi_146_ | ~PKSi_54_;
  assign n2520 = (~n1140 & n2685) | (n1139_1 & (~n1140 | ~n2685));
  assign n2521 = ~PKSi_167_ | ~PKSi_63_;
  assign n2522 = (~n1140 & n2686) | (n1139_1 & (~n1140 | ~n2686));
  assign n2523 = ~PKSi_154_ | ~PKSi_53_;
  assign n2524 = (~n1140 & n2687) | (n1139_1 & (~n1140 | ~n2687));
  assign n2525 = ~PKSi_160_ | ~PKSi_57_;
  assign n2526 = (~n1140 & n2688) | (n1139_1 & (~n1140 | ~n2688));
  assign n2527 = ~PKSi_67_ | ~N_N2921;
  assign n2528 = (~n1140 & n2689) | (n1139_1 & (~n1140 | ~n2689));
  assign n2529 = ~PKSi_165_ | ~PKSi_65_;
  assign n2530 = (~n1140 & n2690) | (n1139_1 & (~n1140 | ~n2690));
  assign n2531 = ~PKSi_147_ | ~N_N2789;
  assign n2532 = (~n1140 & n2691) | (n1139_1 & (~n1140 | ~n2691));
  assign n2533 = ~PKSi_59_ | ~N_N2917;
  assign n2534 = (~n1140 & n2692) | (n1139_1 & (~n1140 | ~n2692));
  assign n2535 = ~PKSi_158_ | ~PKSi_50_;
  assign n2536 = (~n1140 & n2693) | (n1139_1 & (~n1140 | ~n2693));
  assign n2537 = ~PKSi_151_ | ~PKSi_62_;
  assign n2538 = (~n1140 & n2694) | (n1139_1 & (~n1140 | ~n2694));
  assign n2539 = ~PKSi_144_ | ~PKSi_70_;
  assign n2540 = (~n1140 & n2695) | (n1139_1 & (~n1140 | ~n2695));
  assign n2541 = ~PKSi_163_ | ~PKSi_48_;
  assign n2542 = (~n1140 & n2696) | (n1139_1 & (~n1140 | ~n2696));
  assign n2543 = ~PKSi_153_ | ~PKSi_56_;
  assign n2544 = (~n1140 & n2697) | (n1139_1 & (~n1140 | ~n2697));
  assign n2545 = ~PKSi_156_ | ~PKSi_66_;
  assign n2546 = (~n1140 & n2698) | (n1139_1 & (~n1140 | ~n2698));
  assign n2547 = ~PKSi_49_ | ~N_N2909;
  assign n2548 = (~n1140 & n2699) | (n1139_1 & (~n1140 | ~n2699));
  assign n2549 = ~PKSi_162_ | ~N_N2779;
  assign n2550 = (~n1140 & n2700) | (n1139_1 & (~n1140 | ~n2700));
  assign n2551 = ~PKSi_148_ | ~PKSi_61_;
  assign n2552 = (~n1140 & n2701) | (n1139_1 & (~n1140 | ~n2701));
  assign n2553 = ~PKSi_155_ | ~PKSi_69_;
  assign n2554 = (~n1140 & n2702) | (n1139_1 & (~n1140 | ~n2702));
  assign n2555 = ~PKSi_157_ | ~PKSi_58_;
  assign n2556 = (~n1140 & n2703) | (n1139_1 & (~n1140 | ~n2703));
  assign n2557 = ~PKSi_164_ | ~N_N2774;
  assign n2558 = (~n1140 & n2704) | (n1139_1 & (~n1140 | ~n2704));
  assign n2559 = ~PKSi_152_ | ~PKSi_60_;
  assign n2560 = (~n1140 & n2705) | (n1139_1 & (~n1140 | ~n2705));
  assign n2561 = ~PKSi_145_ | ~PKSi_51_;
  assign n2562 = (~n1140 & n2706) | (n1139_1 & (~n1140 | ~n2706));
  assign n2563 = ~PKSi_161_ | ~N_N2770;
  assign n2564 = (~n1140 & n2707) | (n1139_1 & (~n1140 | ~n2707));
  assign n2565 = ~PKSi_64_ | ~N_N2899;
  assign n2566 = (~n1140 & n2708) | (n1139_1 & (~n1140 | ~n2708));
  assign n2567 = ~PKSi_149_ | ~PKSi_68_;
  assign n2568 = (~n1140 & n2709) | (n1139_1 & (~n1140 | ~n2709));
  assign n2569 = ~PKSi_159_ | ~PKSi_55_;
  assign n2570 = (~n1140 & n2710) | (n1139_1 & (~n1140 | ~n2710));
  assign n2571 = ~PKSi_190_ | ~PKSi_76_;
  assign n2572 = (~n1140 & n2711) | (n1139_1 & (~n1140 | ~n2711));
  assign n2573 = ~PKSi_174_ | ~PKSi_95_;
  assign n2574 = (~n1140 & n2712) | (n1139_1 & (~n1140 | ~n2712));
  assign n2575 = ~PKSi_170_ | ~PKSi_78_;
  assign n2576 = (~n1140 & n2713) | (n1139_1 & (~n1140 | ~n2713));
  assign n2577 = ~\[234]  | ~PKSi_87_;
  assign n2578 = (~n1140 & n2714) | (n1139_1 & (~n1140 | ~n2714));
  assign n2579 = ~PKSi_178_ | ~PKSi_77_;
  assign n2580 = (~n1140 & n2715) | (n1139_1 & (~n1140 | ~n2715));
  assign n2581 = ~PKSi_184_ | ~PKSi_81_;
  assign n2582 = (~n1140 & n2716) | (n1139_1 & (~n1140 | ~n2716));
  assign n2583 = ~PKSi_91_ | ~N_N2889;
  assign n2584 = (~n1140 & n2717) | (n1139_1 & (~n1140 | ~n2717));
  assign n2585 = ~PKSi_189_ | ~PKSi_89_;
  assign n2586 = (~n1140 & n2718) | (n1139_1 & (~n1140 | ~n2718));
  assign n2587 = ~PKSi_171_ | ~N_N2757;
  assign n2588 = (~n1140 & n2719) | (n1139_1 & (~n1140 | ~n2719));
  assign n2589 = ~PKSi_83_ | ~N_N2885;
  assign n2590 = (~n1140 & n2720) | (n1139_1 & (~n1140 | ~n2720));
  assign n2591 = ~PKSi_182_ | ~PKSi_74_;
  assign n2592 = (~n1140 & n2721) | (n1139_1 & (~n1140 | ~n2721));
  assign n2593 = ~PKSi_175_ | ~PKSi_86_;
  assign n2594 = (~n1140 & n2722) | (n1139_1 & (~n1140 | ~n2722));
  assign n2595 = ~PKSi_94_ | ~N_N2881;
  assign n2596 = (~n1140 & n2723) | (n1139_1 & (~n1140 | ~n2723));
  assign n2597 = ~PKSi_72_ | ~N_N2879;
  assign n2598 = (~n1140 & n2724) | (n1139_1 & (~n1140 | ~n2724));
  assign n2599 = ~PKSi_80_ | ~N_N2877;
  assign n2600 = (~n1140 & n2725) | (n1139_1 & (~n1140 | ~n2725));
  assign n2601 = ~PKSi_180_ | ~N_N2749;
  assign n2602 = (~n1140 & n2726) | (n1139_1 & (~n1140 | ~n2726));
  assign n2603 = ~PKSi_177_ | ~PKSi_73_;
  assign n2604 = (~n1140 & n2727) | (n1139_1 & (~n1140 | ~n2727));
  assign n2605 = ~PKSi_186_ | ~N_N2746;
  assign n2606 = (~n1140 & n2728) | (n1139_1 & (~n1140 | ~n2728));
  assign n2607 = ~PKSi_172_ | ~PKSi_85_;
  assign n2608 = (~n1140 & n2729) | (n1139_1 & (~n1140 | ~n2729));
  assign n2609 = ~PKSi_179_ | ~PKSi_93_;
  assign n2610 = (~n1140 & n2730) | (n1139_1 & (~n1140 | ~n2730));
  assign n2611 = ~\[253]  | ~PKSi_82_;
  assign n2612 = (~n1140 & n2731) | (n1139_1 & (~n1140 | ~n2731));
  assign n2613 = ~PKSi_188_ | ~N_N2741;
  assign n2614 = (~n1140 & n2732) | (n1139_1 & (~n1140 | ~n2732));
  assign n2615 = ~PKSi_176_ | ~PKSi_84_;
  assign n2616 = (~n1140 & n2733) | (n1139_1 & (~n1140 | ~n2733));
  assign n2617 = ~PKSi_169_ | ~PKSi_75_;
  assign n2618 = (~n1140 & n2734) | (n1139_1 & (~n1140 | ~n2734));
  assign n2619 = ~PKSi_185_ | ~N_N2737;
  assign n2620 = (~n1140 & n2735) | (n1139_1 & (~n1140 | ~n2735));
  assign n2621 = ~\[333]  | ~N_N2865;
  assign n2622 = (~n1140 & n2736) | (n1139_1 & (~n1140 | ~n2736));
  assign n2623 = ~PKSi_173_ | ~PKSi_92_;
  assign n2624 = (~n1140 & n2737) | (n1139_1 & (~n1140 | ~n2737));
  assign n2625 = ~PKSi_183_ | ~PKSi_79_;
  assign n2626 = (~n1140 & n2738) | (n1139_1 & (~n1140 | ~n2738));
  assign n2627 = PKSi_4_ | PKSi_118_;
  assign n2628 = PKSi_23_ | PKSi_102_;
  assign n2629 = PKSi_6_ | PKSi_98_;
  assign n2630 = PKSi_15_ | PKSi_119_;
  assign n2631 = PKSi_5_ | PKSi_106_;
  assign n2632 = PKSi_9_ | PKSi_112_;
  assign n2633 = PKSi_19_ | N_N2986;
  assign n2634 = PKSi_17_ | PKSi_117_;
  assign n2635 = N_N2853 | PKSi_99_;
  assign n2636 = PKSi_11_ | N_N2982;
  assign n2637 = PKSi_2_ | PKSi_110_;
  assign n2638 = PKSi_14_ | PKSi_103_;
  assign n2639 = PKSi_22_ | PKSi_96_;
  assign n2640 = PKSi_0_ | PKSi_115_;
  assign n2641 = PKSi_8_ | N_N2976;
  assign n2642 = PKSi_18_ | PKSi_108_;
  assign n2643 = PKSi_1_ | PKSi_105_;
  assign n2644 = N_N2843 | PKSi_114_;
  assign n2645 = PKSi_13_ | PKSi_100_;
  assign n2646 = PKSi_21_ | PKSi_107_;
  assign n2647 = PKSi_10_ | PKSi_109_;
  assign n2648 = N_N2838 | PKSi_116_;
  assign n2649 = PKSi_12_ | PKSi_104_;
  assign n2650 = PKSi_3_ | PKSi_97_;
  assign n2651 = N_N2834 | PKSi_113_;
  assign n2652 = PKSi_16_ | N_N2964;
  assign n2653 = PKSi_20_ | PKSi_101_;
  assign n2654 = PKSi_7_ | PKSi_111_;
  assign n2655 = PKSi_28_ | PKSi_142_;
  assign n2656 = PKSi_47_ | PKSi_126_;
  assign n2657 = PKSi_30_ | PKSi_122_;
  assign n2658 = PKSi_39_ | \[282] ;
  assign n2659 = PKSi_29_ | PKSi_130_;
  assign n2660 = PKSi_33_ | PKSi_136_;
  assign n2661 = PKSi_43_ | N_N2954;
  assign n2662 = PKSi_41_ | PKSi_141_;
  assign n2663 = N_N2821 | PKSi_123_;
  assign n2664 = PKSi_35_ | N_N2950;
  assign n2665 = PKSi_26_ | PKSi_134_;
  assign n2666 = PKSi_38_ | PKSi_127_;
  assign n2667 = PKSi_46_ | PKSi_120_;
  assign n2668 = PKSi_24_ | N_N2945;
  assign n2669 = PKSi_32_ | N_N2943;
  assign n2670 = PKSi_42_ | PKSi_132_;
  assign n2671 = PKSi_25_ | PKSi_129_;
  assign n2672 = N_N2811 | PKSi_138_;
  assign n2673 = PKSi_37_ | PKSi_124_;
  assign n2674 = PKSi_45_ | PKSi_131_;
  assign n2675 = PKSi_34_ | PKSi_133_;
  assign n2676 = N_N2806 | PKSi_140_;
  assign n2677 = PKSi_36_ | PKSi_128_;
  assign n2678 = PKSi_27_ | PKSi_121_;
  assign n2679 = N_N2802 | PKSi_137_;
  assign n2680 = PKSi_40_ | N_N2931;
  assign n2681 = PKSi_44_ | PKSi_125_;
  assign n2682 = PKSi_31_ | PKSi_135_;
  assign n2683 = PKSi_52_ | PKSi_166_;
  assign n2684 = PKSi_71_ | PKSi_150_;
  assign n2685 = PKSi_54_ | PKSi_146_;
  assign n2686 = PKSi_63_ | PKSi_167_;
  assign n2687 = PKSi_53_ | PKSi_154_;
  assign n2688 = PKSi_57_ | PKSi_160_;
  assign n2689 = PKSi_67_ | N_N2921;
  assign n2690 = PKSi_65_ | PKSi_165_;
  assign n2691 = N_N2789 | PKSi_147_;
  assign n2692 = PKSi_59_ | N_N2917;
  assign n2693 = PKSi_50_ | PKSi_158_;
  assign n2694 = PKSi_62_ | PKSi_151_;
  assign n2695 = PKSi_70_ | PKSi_144_;
  assign n2696 = PKSi_48_ | PKSi_163_;
  assign n2697 = PKSi_56_ | PKSi_153_;
  assign n2698 = PKSi_66_ | PKSi_156_;
  assign n2699 = PKSi_49_ | N_N2909;
  assign n2700 = N_N2779 | PKSi_162_;
  assign n2701 = PKSi_61_ | PKSi_148_;
  assign n2702 = PKSi_69_ | PKSi_155_;
  assign n2703 = PKSi_58_ | PKSi_157_;
  assign n2704 = N_N2774 | PKSi_164_;
  assign n2705 = PKSi_60_ | PKSi_152_;
  assign n2706 = PKSi_51_ | PKSi_145_;
  assign n2707 = N_N2770 | PKSi_161_;
  assign n2708 = PKSi_64_ | N_N2899;
  assign n2709 = PKSi_68_ | PKSi_149_;
  assign n2710 = PKSi_55_ | PKSi_159_;
  assign n2711 = PKSi_76_ | PKSi_190_;
  assign n2712 = PKSi_95_ | PKSi_174_;
  assign n2713 = PKSi_78_ | PKSi_170_;
  assign n2714 = PKSi_87_ | \[234] ;
  assign n2715 = PKSi_77_ | PKSi_178_;
  assign n2716 = PKSi_81_ | PKSi_184_;
  assign n2717 = PKSi_91_ | N_N2889;
  assign n2718 = PKSi_89_ | PKSi_189_;
  assign n2719 = N_N2757 | PKSi_171_;
  assign n2720 = PKSi_83_ | N_N2885;
  assign n2721 = PKSi_74_ | PKSi_182_;
  assign n2722 = PKSi_86_ | PKSi_175_;
  assign n2723 = PKSi_94_ | N_N2881;
  assign n2724 = PKSi_72_ | N_N2879;
  assign n2725 = PKSi_80_ | N_N2877;
  assign n2726 = N_N2749 | PKSi_180_;
  assign n2727 = PKSi_73_ | PKSi_177_;
  assign n2728 = N_N2746 | PKSi_186_;
  assign n2729 = PKSi_85_ | PKSi_172_;
  assign n2730 = PKSi_93_ | PKSi_179_;
  assign n2731 = PKSi_82_ | \[253] ;
  assign n2732 = N_N2741 | PKSi_188_;
  assign n2733 = PKSi_84_ | PKSi_176_;
  assign n2734 = PKSi_75_ | PKSi_169_;
  assign n2735 = N_N2737 | PKSi_185_;
  assign n2736 = \[333]  | N_N2865;
  assign n2737 = PKSi_92_ | PKSi_173_;
  assign n2738 = PKSi_79_ | PKSi_183_;
  assign n2739 = (Pcount_0_ & n2177) | (Pencrypt_0_ & (~Pcount_0_ | n2177));
  assign n2740 = Pcount_0_ | n2177;
  assign n2741 = Pcount_1_ | Pcount_2_;
  assign PKSi_191_ = \[234] ;
  assign PKSi_187_ = \[234] ;
  assign PKSi_181_ = \[253] ;
  assign PKSi_168_ = \[253] ;
  assign PKSi_143_ = \[282] ;
  assign PKSi_139_ = \[282] ;
  assign PKSi_90_ = \[333] ;
  assign PKSi_88_ = \[333] ;
  always @ (posedge clock) begin
    PKSi_79_ <= n921;
    PKSi_92_ <= n925_1;
    \[333]  <= n929_1;
    N_N2737 <= n934_1;
    PKSi_75_ <= n939_1;
    PKSi_84_ <= n943;
    N_N2741 <= n947;
    PKSi_82_ <= n952_1;
    PKSi_93_ <= n956_1;
    PKSi_85_ <= n960_1;
    N_N2746 <= n964_1;
    PKSi_73_ <= n969;
    N_N2749 <= n973;
    PKSi_80_ <= n978_1;
    PKSi_72_ <= n982_1;
    PKSi_94_ <= n986_1;
    PKSi_86_ <= n990_1;
    PKSi_74_ <= n994_1;
    PKSi_83_ <= n998_1;
    N_N2757 <= n1002_1;
    PKSi_89_ <= n1007;
    PKSi_91_ <= n1011;
    PKSi_81_ <= n1015;
    PKSi_77_ <= n1019;
    PKSi_87_ <= n1023;
    PKSi_78_ <= n1027;
    PKSi_95_ <= n1031;
    PKSi_76_ <= n1035;
    PKSi_55_ <= n1039;
    PKSi_68_ <= n1043;
    PKSi_64_ <= n1047;
    N_N2770 <= n1051;
    PKSi_51_ <= n1056_1;
    PKSi_60_ <= n1060_1;
    N_N2774 <= n1064_1;
    PKSi_58_ <= n1069;
    PKSi_69_ <= n1073;
    PKSi_61_ <= n1077;
    N_N2779 <= n1081;
    PKSi_49_ <= n1086_1;
    PKSi_66_ <= n1090_1;
    PKSi_56_ <= n1094_1;
    PKSi_48_ <= n1098_1;
    PKSi_70_ <= n1102_1;
    PKSi_62_ <= n1106_1;
    PKSi_50_ <= n1110_1;
    PKSi_59_ <= n1114_1;
    N_N2789 <= n1118_1;
    PKSi_65_ <= n1123;
    PKSi_67_ <= n1127;
    PKSi_57_ <= n1131;
    PKSi_53_ <= n1135;
    PKSi_63_ <= n1139;
    PKSi_54_ <= n1143;
    PKSi_71_ <= n1147;
    PKSi_52_ <= n1151;
    PKSi_31_ <= n1155;
    PKSi_44_ <= n1159;
    PKSi_40_ <= n1163;
    N_N2802 <= n1167_1;
    PKSi_27_ <= n1172;
    PKSi_36_ <= n1176;
    N_N2806 <= n1180;
    PKSi_34_ <= n1185;
    PKSi_45_ <= n1189;
    PKSi_37_ <= n1193;
    N_N2811 <= n1197;
    PKSi_25_ <= n1202;
    PKSi_42_ <= n1206;
    PKSi_32_ <= n1210;
    PKSi_24_ <= n1214;
    PKSi_46_ <= n1218;
    PKSi_38_ <= n1222;
    PKSi_26_ <= n1226;
    PKSi_35_ <= n1230;
    N_N2821 <= n1234;
    PKSi_41_ <= n1239;
    PKSi_43_ <= n1243;
    PKSi_33_ <= n1247;
    PKSi_29_ <= n1251;
    PKSi_39_ <= n1255;
    PKSi_30_ <= n1259;
    PKSi_47_ <= n1263;
    PKSi_28_ <= n1267;
    PKSi_7_ <= n1271;
    PKSi_20_ <= n1275;
    PKSi_16_ <= n1279;
    N_N2834 <= n1283;
    PKSi_3_ <= n1288;
    PKSi_12_ <= n1292_1;
    N_N2838 <= n1296_1;
    PKSi_10_ <= n1301_1;
    PKSi_21_ <= n1305_1;
    PKSi_13_ <= n1309_1;
    N_N2843 <= n1313_1;
    PKSi_1_ <= n1318_1;
    PKSi_18_ <= n1322_1;
    PKSi_8_ <= n1326_1;
    PKSi_0_ <= n1330_1;
    PKSi_22_ <= n1334_1;
    PKSi_14_ <= n1338_1;
    PKSi_2_ <= n1342_1;
    PKSi_11_ <= n1346_1;
    N_N2853 <= n1350_1;
    PKSi_17_ <= n1355_1;
    PKSi_19_ <= n1359_1;
    PKSi_9_ <= n1363_1;
    PKSi_5_ <= n1367_1;
    PKSi_15_ <= n1371_1;
    PKSi_6_ <= n1375_1;
    PKSi_23_ <= n1379_1;
    PKSi_4_ <= n1383_1;
    PKSi_183_ <= n1387_1;
    PKSi_173_ <= n1391_1;
    N_N2865 <= n1395_1;
    PKSi_185_ <= n1400_1;
    PKSi_169_ <= n1404_1;
    PKSi_176_ <= n1408_1;
    PKSi_188_ <= n1412_1;
    \[253]  <= n1416_1;
    PKSi_179_ <= n1421_1;
    PKSi_172_ <= n1425_1;
    PKSi_186_ <= n1429_1;
    PKSi_177_ <= n1433_1;
    PKSi_180_ <= n1437_1;
    N_N2877 <= n1441_1;
    N_N2879 <= n1446_1;
    N_N2881 <= n1451_1;
    PKSi_175_ <= n1456_1;
    PKSi_182_ <= n1460_1;
    N_N2885 <= n1464_1;
    PKSi_171_ <= n1469_1;
    PKSi_189_ <= n1473_1;
    N_N2889 <= n1477_1;
    PKSi_184_ <= n1482_1;
    PKSi_178_ <= n1486_1;
    \[234]  <= n1490_1;
    PKSi_170_ <= n1495_1;
    PKSi_174_ <= n1499_1;
    PKSi_190_ <= n1503_1;
    PKSi_159_ <= n1507_1;
    PKSi_149_ <= n1511_1;
    N_N2899 <= n1515;
    PKSi_161_ <= n1520_1;
    PKSi_145_ <= n1524_1;
    PKSi_152_ <= n1528_1;
    PKSi_164_ <= n1532_1;
    PKSi_157_ <= n1536_1;
    PKSi_155_ <= n1540_1;
    PKSi_148_ <= n1544_1;
    PKSi_162_ <= n1548_1;
    N_N2909 <= n1552_1;
    PKSi_156_ <= n1557_1;
    PKSi_153_ <= n1561_1;
    PKSi_163_ <= n1565_1;
    PKSi_144_ <= n1569_1;
    PKSi_151_ <= n1573_1;
    PKSi_158_ <= n1577_1;
    N_N2917 <= n1581_1;
    PKSi_147_ <= n1586_1;
    PKSi_165_ <= n1590_1;
    N_N2921 <= n1594_1;
    PKSi_160_ <= n1599_1;
    PKSi_154_ <= n1603_1;
    PKSi_167_ <= n1607_1;
    PKSi_146_ <= n1611_1;
    PKSi_150_ <= n1615_1;
    PKSi_166_ <= n1619_1;
    PKSi_135_ <= n1623_1;
    PKSi_125_ <= n1627_1;
    N_N2931 <= n1631_1;
    PKSi_137_ <= n1636_1;
    PKSi_121_ <= n1640_1;
    PKSi_128_ <= n1644_1;
    PKSi_140_ <= n1648_1;
    PKSi_133_ <= n1652_1;
    PKSi_131_ <= n1656_1;
    PKSi_124_ <= n1660_1;
    PKSi_138_ <= n1664_1;
    PKSi_129_ <= n1668_1;
    PKSi_132_ <= n1672_1;
    N_N2943 <= n1676_1;
    N_N2945 <= n1681_1;
    PKSi_120_ <= n1686_1;
    PKSi_127_ <= n1690_1;
    PKSi_134_ <= n1694_1;
    N_N2950 <= n1698_1;
    PKSi_123_ <= n1703_1;
    PKSi_141_ <= n1707_1;
    N_N2954 <= n1711_1;
    PKSi_136_ <= n1716_1;
    PKSi_130_ <= n1720_1;
    \[282]  <= n1724_1;
    PKSi_122_ <= n1729_1;
    PKSi_126_ <= n1733_1;
    PKSi_142_ <= n1737_1;
    PKSi_111_ <= n1741_1;
    PKSi_101_ <= n1745;
    N_N2964 <= n1749;
    PKSi_113_ <= n1754_1;
    PKSi_97_ <= n1758_1;
    PKSi_104_ <= n1762_1;
    PKSi_116_ <= n1766_1;
    PKSi_109_ <= n1770_1;
    PKSi_107_ <= n1774_1;
    PKSi_100_ <= n1778_1;
    PKSi_114_ <= n1782_1;
    PKSi_105_ <= n1786_1;
    PKSi_108_ <= n1790_1;
    N_N2976 <= n1794_1;
    PKSi_115_ <= n1799;
    PKSi_96_ <= n1803;
    PKSi_103_ <= n1807;
    PKSi_110_ <= n1811;
    N_N2982 <= n1815;
    PKSi_99_ <= n1820_1;
    PKSi_117_ <= n1824_1;
    N_N2986 <= n1828_1;
    PKSi_112_ <= n1833;
    PKSi_106_ <= n1837;
    PKSi_119_ <= n1841;
    PKSi_98_ <= n1845;
    PKSi_102_ <= n1849;
    PKSi_118_ <= n1853;
  end
endmodule


