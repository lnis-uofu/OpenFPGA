`ifndef "BITSTREAM_andgate"
`define "BITSTREAM_andgate"


class bitstream_andgate extends bs_base_seq;
   `uvm_object_utils(bitstream_andgate)
   
   /**
    * Default constructor.
    */
   extern function new(string name="bitstream_andgate");
   /**
    * Sequence body
    */
   extern virtual task body();

endclass : bitstream_andgate

function bitstream_andgate::new(string name = "bitstream_andgate");

      super.new(name);

endfunction // new

task bitstream_andgate::body();
// ----- Configuration chain default input -----
		prog_cycle_task(16'b0000000000000000, 1'b1);
		prog_cycle_task(16'b0100000000000000, 1'b1);
		prog_cycle_task(16'b0010000000000000, 1'b1);
		prog_cycle_task(16'b0110000000000000, 1'b1);
		prog_cycle_task(16'b0001000000000000, 1'b1);
		prog_cycle_task(16'b0101000000000000, 1'b1);
		prog_cycle_task(16'b0011000000000000, 1'b1);
		prog_cycle_task(16'b0111000000000000, 1'b1);
		prog_cycle_task(16'b0000000000100000, 1'b1);
		prog_cycle_task(16'b0100000000100000, 1'b1);
		prog_cycle_task(16'b0010000000100000, 1'b1);
		prog_cycle_task(16'b0110000000100000, 1'b1);
		prog_cycle_task(16'b0001000000100000, 1'b1);
		prog_cycle_task(16'b0101000000100000, 1'b1);
		prog_cycle_task(16'b0011000000100000, 1'b0);
		prog_cycle_task(16'b0111000000100000, 1'b1);
		prog_cycle_task(16'b0000000000010000, 1'b1);
		prog_cycle_task(16'b0100000000010000, 1'b1);
		prog_cycle_task(16'b0010000000010000, 1'b1);
		prog_cycle_task(16'b0110000000010000, 1'b1);
		prog_cycle_task(16'b0001000000010000, 1'b1);
		prog_cycle_task(16'b0101000000010000, 1'b1);
		prog_cycle_task(16'b0011000000010000, 1'b1);
		prog_cycle_task(16'b0111000000010000, 1'b1);
		prog_cycle_task(16'b0000000000110000, 1'b1);
		prog_cycle_task(16'b0100000000110000, 1'b1);
		prog_cycle_task(16'b0010000000110000, 1'b1);
		prog_cycle_task(16'b0110000000110000, 1'b1);
		prog_cycle_task(16'b0001000000110000, 1'b1);
		prog_cycle_task(16'b0101000000110000, 1'b1);
		prog_cycle_task(16'b0011000000110000, 1'b1);
		prog_cycle_task(16'b0111000000110000, 1'b1);
		prog_cycle_task(16'b0000000000001000, 1'b1);
		prog_cycle_task(16'b1000000000001000, 1'b1);
		prog_cycle_task(16'b0100000000001000, 1'b1);
		prog_cycle_task(16'b1100000000001000, 1'b1);
		prog_cycle_task(16'b0010000000001000, 1'b1);
		prog_cycle_task(16'b1010000000001000, 1'b1);
		prog_cycle_task(16'b0110000000001000, 1'b1);
		prog_cycle_task(16'b1110000000001000, 1'b1);
		prog_cycle_task(16'b0001000000001000, 1'b1);
		prog_cycle_task(16'b1001000000001000, 1'b1);
		prog_cycle_task(16'b0101000000001000, 1'b1);
		prog_cycle_task(16'b1101000000001000, 1'b1);
		prog_cycle_task(16'b0011000000001000, 1'b1);
		prog_cycle_task(16'b1011000000001000, 1'b1);
		prog_cycle_task(16'b0111000000001000, 1'b1);
		prog_cycle_task(16'b1111000000001000, 1'b1);
		prog_cycle_task(16'b0000100000001000, 1'b1);
		prog_cycle_task(16'b1000100000001000, 1'b1);
		prog_cycle_task(16'b0100100000001000, 1'b1);
		prog_cycle_task(16'b1100100000001000, 1'b1);
		prog_cycle_task(16'b0010100000001000, 1'b1);
		prog_cycle_task(16'b1010100000001000, 1'b1);
		prog_cycle_task(16'b0110100000001000, 1'b0);
		prog_cycle_task(16'b1110100000001000, 1'b1);
		prog_cycle_task(16'b0001100000001000, 1'b1);
		prog_cycle_task(16'b1001100000001000, 1'b1);
		prog_cycle_task(16'b0101100000001000, 1'b0);
		prog_cycle_task(16'b1101100000001000, 1'b1);
		prog_cycle_task(16'b0011100000001000, 1'b1);
		prog_cycle_task(16'b1011100000001000, 1'b1);
		prog_cycle_task(16'b0111100000001000, 1'b1);
		prog_cycle_task(16'b1111100000001000, 1'b1);
		prog_cycle_task(16'b0000010000001000, 1'b1);
		prog_cycle_task(16'b1000010000001000, 1'b1);
		prog_cycle_task(16'b0100010000001000, 1'b1);
		prog_cycle_task(16'b1100010000001000, 1'b1);
		prog_cycle_task(16'b0000000000101000, 1'b1);
		prog_cycle_task(16'b1000000000101000, 1'b0);
		prog_cycle_task(16'b0100000000101000, 1'b0);
		prog_cycle_task(16'b1100000000101000, 1'b1);
		prog_cycle_task(16'b0010000000101000, 1'b0);
		prog_cycle_task(16'b1010000000101000, 1'b0);
		prog_cycle_task(16'b0001000000101000, 1'b1);
		prog_cycle_task(16'b1001000000101000, 1'b0);
		prog_cycle_task(16'b0101000000101000, 1'b0);
		prog_cycle_task(16'b1101000000101000, 1'b1);
		prog_cycle_task(16'b0011000000101000, 1'b0);
		prog_cycle_task(16'b1011000000101000, 1'b0);
		prog_cycle_task(16'b0000100000101000, 1'b1);
		prog_cycle_task(16'b1000100000101000, 1'b0);
		prog_cycle_task(16'b0100100000101000, 1'b0);
		prog_cycle_task(16'b1100100000101000, 1'b1);
		prog_cycle_task(16'b0010100000101000, 1'b0);
		prog_cycle_task(16'b1010100000101000, 1'b0);
		prog_cycle_task(16'b0001100000101000, 1'b1);
		prog_cycle_task(16'b1001100000101000, 1'b0);
		prog_cycle_task(16'b0101100000101000, 1'b0);
		prog_cycle_task(16'b1101100000101000, 1'b1);
		prog_cycle_task(16'b0011100000101000, 1'b0);
		prog_cycle_task(16'b1011100000101000, 1'b0);
		prog_cycle_task(16'b0000010000101000, 1'b1);
		prog_cycle_task(16'b1000010000101000, 1'b0);
		prog_cycle_task(16'b0100010000101000, 1'b0);
		prog_cycle_task(16'b1100010000101000, 1'b1);
		prog_cycle_task(16'b0010010000101000, 1'b0);
		prog_cycle_task(16'b1010010000101000, 1'b0);
		prog_cycle_task(16'b0001010000101000, 1'b1);
		prog_cycle_task(16'b1001010000101000, 1'b0);
		prog_cycle_task(16'b0101010000101000, 1'b0);
		prog_cycle_task(16'b1101010000101000, 1'b1);
		prog_cycle_task(16'b0011010000101000, 1'b0);
		prog_cycle_task(16'b1011010000101000, 1'b0);
		prog_cycle_task(16'b0000110000101000, 1'b1);
		prog_cycle_task(16'b1000110000101000, 1'b0);
		prog_cycle_task(16'b0100110000101000, 1'b0);
		prog_cycle_task(16'b1100110000101000, 1'b1);
		prog_cycle_task(16'b0010110000101000, 1'b0);
		prog_cycle_task(16'b1010110000101000, 1'b0);
		prog_cycle_task(16'b0001110000101000, 1'b1);
		prog_cycle_task(16'b1001110000101000, 1'b0);
		prog_cycle_task(16'b0101110000101000, 1'b0);
		prog_cycle_task(16'b1101110000101000, 1'b1);
		prog_cycle_task(16'b0011110000101000, 1'b0);
		prog_cycle_task(16'b1011110000101000, 1'b0);
		prog_cycle_task(16'b0000001000101000, 1'b1);
		prog_cycle_task(16'b1000001000101000, 1'b0);
		prog_cycle_task(16'b0100001000101000, 1'b0);
		prog_cycle_task(16'b1100001000101000, 1'b1);
		prog_cycle_task(16'b0010001000101000, 1'b0);
		prog_cycle_task(16'b1010001000101000, 1'b0);
		prog_cycle_task(16'b0001001000101000, 1'b1);
		prog_cycle_task(16'b1001001000101000, 1'b1);
		prog_cycle_task(16'b0000101000101000, 1'b1);
		prog_cycle_task(16'b1000101000101000, 1'b1);
		prog_cycle_task(16'b0000000000011000, 1'b1);
		prog_cycle_task(16'b0100000000011000, 1'b1);
		prog_cycle_task(16'b0010000000011000, 1'b1);
		prog_cycle_task(16'b0110000000011000, 1'b1);
		prog_cycle_task(16'b0001000000011000, 1'b1);
		prog_cycle_task(16'b0101000000011000, 1'b1);
		prog_cycle_task(16'b0011000000011000, 1'b1);
		prog_cycle_task(16'b0111000000011000, 1'b1);
		prog_cycle_task(16'b0000000000111000, 1'b1);
		prog_cycle_task(16'b1000000000111000, 1'b0);
		prog_cycle_task(16'b0100000000111000, 1'b0);
		prog_cycle_task(16'b1100000000111000, 1'b1);
		prog_cycle_task(16'b0010000000111000, 1'b0);
		prog_cycle_task(16'b1010000000111000, 1'b0);
		prog_cycle_task(16'b0001000000111000, 1'b1);
		prog_cycle_task(16'b1001000000111000, 1'b0);
		prog_cycle_task(16'b0101000000111000, 1'b0);
		prog_cycle_task(16'b1101000000111000, 1'b1);
		prog_cycle_task(16'b0011000000111000, 1'b0);
		prog_cycle_task(16'b1011000000111000, 1'b0);
		prog_cycle_task(16'b0000100000111000, 1'b1);
		prog_cycle_task(16'b1000100000111000, 1'b0);
		prog_cycle_task(16'b0100100000111000, 1'b0);
		prog_cycle_task(16'b1100100000111000, 1'b1);
		prog_cycle_task(16'b0010100000111000, 1'b0);
		prog_cycle_task(16'b1010100000111000, 1'b0);
		prog_cycle_task(16'b0001100000111000, 1'b1);
		prog_cycle_task(16'b1001100000111000, 1'b1);
		prog_cycle_task(16'b0000010000111000, 1'b1);
		prog_cycle_task(16'b1000010000111000, 1'b1);
		prog_cycle_task(16'b0001010000111000, 1'b1);
		prog_cycle_task(16'b1001010000111000, 1'b1);
		prog_cycle_task(16'b0000110000111000, 1'b1);
		prog_cycle_task(16'b1000110000111000, 1'b1);
		prog_cycle_task(16'b0001110000111000, 1'b1);
		prog_cycle_task(16'b1001110000111000, 1'b1);
		prog_cycle_task(16'b0000001000111000, 1'b1);
		prog_cycle_task(16'b1000001000111000, 1'b1);
		prog_cycle_task(16'b0001001000111000, 1'b1);
		prog_cycle_task(16'b1001001000111000, 1'b1);
		prog_cycle_task(16'b0000101000111000, 1'b1);
		prog_cycle_task(16'b1000101000111000, 1'b1);
		prog_cycle_task(16'b0001101000111000, 1'b1);
		prog_cycle_task(16'b1001101000111000, 1'b1);
		prog_cycle_task(16'b0000011000111000, 1'b1);
		prog_cycle_task(16'b1000011000111000, 1'b0);
		prog_cycle_task(16'b0100011000111000, 1'b0);
		prog_cycle_task(16'b1100011000111000, 1'b1);
		prog_cycle_task(16'b0010011000111000, 1'b0);
		prog_cycle_task(16'b1010011000111000, 1'b0);
		prog_cycle_task(16'b0001011000111000, 1'b1);
		prog_cycle_task(16'b1001011000111000, 1'b0);
		prog_cycle_task(16'b0101011000111000, 1'b0);
		prog_cycle_task(16'b1101011000111000, 1'b1);
		prog_cycle_task(16'b0011011000111000, 1'b0);
		prog_cycle_task(16'b1011011000111000, 1'b0);
		prog_cycle_task(16'b0000111000111000, 1'b1);
		prog_cycle_task(16'b1000111000111000, 1'b0);
		prog_cycle_task(16'b0100111000111000, 1'b0);
		prog_cycle_task(16'b1100111000111000, 1'b1);
		prog_cycle_task(16'b0010111000111000, 1'b0);
		prog_cycle_task(16'b1010111000111000, 1'b0);
		prog_cycle_task(16'b0000000000000100, 1'b1);
		prog_cycle_task(16'b1000000000000100, 1'b0);
		prog_cycle_task(16'b0100000000000100, 1'b0);
		prog_cycle_task(16'b1100000000000100, 1'b1);
		prog_cycle_task(16'b0010000000000100, 1'b0);
		prog_cycle_task(16'b1010000000000100, 1'b0);
		prog_cycle_task(16'b0001000000000100, 1'b1);
		prog_cycle_task(16'b1001000000000100, 1'b0);
		prog_cycle_task(16'b0101000000000100, 1'b0);
		prog_cycle_task(16'b1101000000000100, 1'b1);
		prog_cycle_task(16'b0011000000000100, 1'b0);
		prog_cycle_task(16'b1011000000000100, 1'b0);
		prog_cycle_task(16'b0000100000000100, 1'b1);
		prog_cycle_task(16'b1000100000000100, 1'b0);
		prog_cycle_task(16'b0100100000000100, 1'b0);
		prog_cycle_task(16'b1100100000000100, 1'b1);
		prog_cycle_task(16'b0010100000000100, 1'b0);
		prog_cycle_task(16'b1010100000000100, 1'b0);
		prog_cycle_task(16'b0001100000000100, 1'b1);
		prog_cycle_task(16'b1001100000000100, 1'b0);
		prog_cycle_task(16'b0101100000000100, 1'b0);
		prog_cycle_task(16'b1101100000000100, 1'b1);
		prog_cycle_task(16'b0011100000000100, 1'b0);
		prog_cycle_task(16'b1011100000000100, 1'b0);
		prog_cycle_task(16'b0000010000000100, 1'b1);
		prog_cycle_task(16'b1000010000000100, 1'b0);
		prog_cycle_task(16'b0100010000000100, 1'b0);
		prog_cycle_task(16'b1100010000000100, 1'b1);
		prog_cycle_task(16'b0010010000000100, 1'b0);
		prog_cycle_task(16'b1010010000000100, 1'b0);
		prog_cycle_task(16'b0001010000000100, 1'b1);
		prog_cycle_task(16'b1001010000000100, 1'b0);
		prog_cycle_task(16'b0101010000000100, 1'b0);
		prog_cycle_task(16'b1101010000000100, 1'b1);
		prog_cycle_task(16'b0011010000000100, 1'b0);
		prog_cycle_task(16'b1011010000000100, 1'b0);
		prog_cycle_task(16'b0000110000000100, 1'b1);
		prog_cycle_task(16'b1000110000000100, 1'b0);
		prog_cycle_task(16'b0100110000000100, 1'b0);
		prog_cycle_task(16'b1100110000000100, 1'b1);
		prog_cycle_task(16'b0010110000000100, 1'b0);
		prog_cycle_task(16'b1010110000000100, 1'b0);
		prog_cycle_task(16'b0001110000000100, 1'b1);
		prog_cycle_task(16'b1001110000000100, 1'b0);
		prog_cycle_task(16'b0101110000000100, 1'b0);
		prog_cycle_task(16'b1101110000000100, 1'b1);
		prog_cycle_task(16'b0011110000000100, 1'b0);
		prog_cycle_task(16'b1011110000000100, 1'b0);
		prog_cycle_task(16'b0000001000000100, 1'b1);
		prog_cycle_task(16'b1000001000000100, 1'b0);
		prog_cycle_task(16'b0100001000000100, 1'b0);
		prog_cycle_task(16'b1100001000000100, 1'b1);
		prog_cycle_task(16'b0010001000000100, 1'b0);
		prog_cycle_task(16'b1010001000000100, 1'b0);
		prog_cycle_task(16'b0001001000000100, 1'b1);
		prog_cycle_task(16'b1001001000000100, 1'b1);
		prog_cycle_task(16'b0000101000000100, 1'b1);
		prog_cycle_task(16'b1000101000000100, 1'b1);
		prog_cycle_task(16'b0000000000100100, 1'b1);
		prog_cycle_task(16'b0100000000100100, 1'b1);
		prog_cycle_task(16'b0010000000100100, 1'b1);
		prog_cycle_task(16'b0110000000100100, 1'b1);
		prog_cycle_task(16'b0001000000100100, 1'b1);
		prog_cycle_task(16'b0101000000100100, 1'b1);
		prog_cycle_task(16'b0011000000100100, 1'b1);
		prog_cycle_task(16'b0111000000100100, 1'b1);
		prog_cycle_task(16'b0000000000010100, 1'b1);
		prog_cycle_task(16'b1000000000010100, 1'b1);
		prog_cycle_task(16'b0100000000010100, 1'b1);
		prog_cycle_task(16'b1100000000010100, 1'b1);
		prog_cycle_task(16'b0010000000010100, 1'b1);
		prog_cycle_task(16'b1010000000010100, 1'b1);
		prog_cycle_task(16'b0110000000010100, 1'b1);
		prog_cycle_task(16'b1110000000010100, 1'b1);
		prog_cycle_task(16'b0001000000010100, 1'b1);
		prog_cycle_task(16'b1001000000010100, 1'b1);
		prog_cycle_task(16'b0101000000010100, 1'b1);
		prog_cycle_task(16'b1101000000010100, 1'b1);
		prog_cycle_task(16'b0011000000010100, 1'b1);
		prog_cycle_task(16'b1011000000010100, 1'b1);
		prog_cycle_task(16'b0111000000010100, 1'b1);
		prog_cycle_task(16'b1111000000010100, 1'b1);
		prog_cycle_task(16'b0000100000010100, 1'b1);
		prog_cycle_task(16'b1000100000010100, 1'b1);
		prog_cycle_task(16'b0100100000010100, 1'b1);
		prog_cycle_task(16'b1100100000010100, 1'b1);
		prog_cycle_task(16'b0010100000010100, 1'b1);
		prog_cycle_task(16'b1010100000010100, 1'b1);
		prog_cycle_task(16'b0110100000010100, 1'b1);
		prog_cycle_task(16'b1110100000010100, 1'b1);
		prog_cycle_task(16'b0001100000010100, 1'b1);
		prog_cycle_task(16'b1001100000010100, 1'b1);
		prog_cycle_task(16'b0101100000010100, 1'b1);
		prog_cycle_task(16'b1101100000010100, 1'b1);
		prog_cycle_task(16'b0011100000010100, 1'b1);
		prog_cycle_task(16'b1011100000010100, 1'b1);
		prog_cycle_task(16'b0111100000010100, 1'b1);
		prog_cycle_task(16'b1111100000010100, 1'b1);
		prog_cycle_task(16'b0000010000010100, 1'b1);
		prog_cycle_task(16'b1000010000010100, 1'b1);
		prog_cycle_task(16'b0100010000010100, 1'b1);
		prog_cycle_task(16'b1100010000010100, 1'b1);
		prog_cycle_task(16'b0000000000110100, 1'b1);
		prog_cycle_task(16'b1000000000110100, 1'b0);
		prog_cycle_task(16'b0100000000110100, 1'b0);
		prog_cycle_task(16'b1100000000110100, 1'b1);
		prog_cycle_task(16'b0010000000110100, 1'b0);
		prog_cycle_task(16'b1010000000110100, 1'b0);
		prog_cycle_task(16'b0001000000110100, 1'b1);
		prog_cycle_task(16'b1001000000110100, 1'b0);
		prog_cycle_task(16'b0101000000110100, 1'b0);
		prog_cycle_task(16'b1101000000110100, 1'b1);
		prog_cycle_task(16'b0011000000110100, 1'b0);
		prog_cycle_task(16'b1011000000110100, 1'b0);
		prog_cycle_task(16'b0000100000110100, 1'b1);
		prog_cycle_task(16'b1000100000110100, 1'b0);
		prog_cycle_task(16'b0100100000110100, 1'b0);
		prog_cycle_task(16'b1100100000110100, 1'b1);
		prog_cycle_task(16'b0010100000110100, 1'b0);
		prog_cycle_task(16'b1010100000110100, 1'b0);
		prog_cycle_task(16'b0001100000110100, 1'b1);
		prog_cycle_task(16'b1001100000110100, 1'b1);
		prog_cycle_task(16'b0000010000110100, 1'b1);
		prog_cycle_task(16'b1000010000110100, 1'b1);
		prog_cycle_task(16'b0001010000110100, 1'b1);
		prog_cycle_task(16'b1001010000110100, 1'b1);
		prog_cycle_task(16'b0000110000110100, 1'b1);
		prog_cycle_task(16'b1000110000110100, 1'b1);
		prog_cycle_task(16'b0001110000110100, 1'b1);
		prog_cycle_task(16'b1001110000110100, 1'b1);
		prog_cycle_task(16'b0000001000110100, 1'b1);
		prog_cycle_task(16'b1000001000110100, 1'b1);
		prog_cycle_task(16'b0001001000110100, 1'b1);
		prog_cycle_task(16'b1001001000110100, 1'b1);
		prog_cycle_task(16'b0000101000110100, 1'b1);
		prog_cycle_task(16'b1000101000110100, 1'b0);
		prog_cycle_task(16'b0100101000110100, 1'b0);
		prog_cycle_task(16'b1100101000110100, 1'b1);
		prog_cycle_task(16'b0010101000110100, 1'b0);
		prog_cycle_task(16'b1010101000110100, 1'b0);
		prog_cycle_task(16'b0001101000110100, 1'b1);
		prog_cycle_task(16'b1001101000110100, 1'b0);
		prog_cycle_task(16'b0101101000110100, 1'b0);
		prog_cycle_task(16'b1101101000110100, 1'b1);
		prog_cycle_task(16'b0011101000110100, 1'b0);
		prog_cycle_task(16'b1011101000110100, 1'b0);
		prog_cycle_task(16'b0000011000110100, 1'b1);
		prog_cycle_task(16'b1000011000110100, 1'b0);
		prog_cycle_task(16'b0100011000110100, 1'b0);
		prog_cycle_task(16'b1100011000110100, 1'b1);
		prog_cycle_task(16'b0010011000110100, 1'b0);
		prog_cycle_task(16'b1010011000110100, 1'b0);
		prog_cycle_task(16'b0000000000001100, 1'b1);
		prog_cycle_task(16'b1000000000001100, 1'b0);
		prog_cycle_task(16'b0100000000001100, 1'b0);
		prog_cycle_task(16'b1100000000001100, 1'b1);
		prog_cycle_task(16'b0010000000001100, 1'b0);
		prog_cycle_task(16'b1010000000001100, 1'b0);
		prog_cycle_task(16'b0001000000001100, 1'b1);
		prog_cycle_task(16'b1001000000001100, 1'b1);
		prog_cycle_task(16'b0000100000001100, 1'b1);
		prog_cycle_task(16'b1000100000001100, 1'b0);
		prog_cycle_task(16'b0100100000001100, 1'b0);
		prog_cycle_task(16'b1100100000001100, 1'b1);
		prog_cycle_task(16'b0010100000001100, 1'b0);
		prog_cycle_task(16'b1010100000001100, 1'b0);
		prog_cycle_task(16'b0001100000001100, 1'b1);
		prog_cycle_task(16'b1001100000001100, 1'b0);
		prog_cycle_task(16'b0101100000001100, 1'b0);
		prog_cycle_task(16'b1101100000001100, 1'b1);
		prog_cycle_task(16'b0011100000001100, 1'b0);
		prog_cycle_task(16'b1011100000001100, 1'b0);
		prog_cycle_task(16'b0000010000001100, 1'b1);
		prog_cycle_task(16'b1000010000001100, 1'b0);
		prog_cycle_task(16'b0100010000001100, 1'b0);
		prog_cycle_task(16'b1100010000001100, 1'b1);
		prog_cycle_task(16'b0010010000001100, 1'b0);
		prog_cycle_task(16'b1010010000001100, 1'b0);
		prog_cycle_task(16'b0001010000001100, 1'b1);
		prog_cycle_task(16'b1001010000001100, 1'b0);
		prog_cycle_task(16'b0101010000001100, 1'b0);
		prog_cycle_task(16'b1101010000001100, 1'b1);
		prog_cycle_task(16'b0011010000001100, 1'b0);
		prog_cycle_task(16'b1011010000001100, 1'b0);
		prog_cycle_task(16'b0000110000001100, 1'b1);
		prog_cycle_task(16'b1000110000001100, 1'b0);
		prog_cycle_task(16'b0100110000001100, 1'b0);
		prog_cycle_task(16'b1100110000001100, 1'b1);
		prog_cycle_task(16'b0010110000001100, 1'b0);
		prog_cycle_task(16'b1010110000001100, 1'b0);
		prog_cycle_task(16'b0001110000001100, 1'b1);
		prog_cycle_task(16'b1001110000001100, 1'b0);
		prog_cycle_task(16'b0101110000001100, 1'b0);
		prog_cycle_task(16'b1101110000001100, 1'b1);
		prog_cycle_task(16'b0011110000001100, 1'b0);
		prog_cycle_task(16'b1011110000001100, 1'b0);
		prog_cycle_task(16'b0000001000001100, 1'b1);
		prog_cycle_task(16'b1000001000001100, 1'b0);
		prog_cycle_task(16'b0100001000001100, 1'b0);
		prog_cycle_task(16'b1100001000001100, 1'b1);
		prog_cycle_task(16'b0010001000001100, 1'b0);
		prog_cycle_task(16'b1010001000001100, 1'b0);
		prog_cycle_task(16'b0001001000001100, 1'b1);
		prog_cycle_task(16'b1001001000001100, 1'b0);
		prog_cycle_task(16'b0101001000001100, 1'b0);
		prog_cycle_task(16'b1101001000001100, 1'b1);
		prog_cycle_task(16'b0011001000001100, 1'b0);
		prog_cycle_task(16'b1011001000001100, 1'b0);
		prog_cycle_task(16'b0000000000101100, 1'b1);
		prog_cycle_task(16'b0100000000101100, 1'b1);
		prog_cycle_task(16'b0010000000101100, 1'b1);
		prog_cycle_task(16'b0110000000101100, 1'b1);
		prog_cycle_task(16'b0001000000101100, 1'b1);
		prog_cycle_task(16'b0101000000101100, 1'b1);
		prog_cycle_task(16'b0011000000101100, 1'b1);
		prog_cycle_task(16'b0111000000101100, 1'b1);
		prog_cycle_task(16'b0000000000011100, 1'b1);
		prog_cycle_task(16'b1000000000011100, 1'b1);
		prog_cycle_task(16'b0100000000011100, 1'b1);
		prog_cycle_task(16'b1100000000011100, 1'b1);
		prog_cycle_task(16'b0010000000011100, 1'b1);
		prog_cycle_task(16'b1010000000011100, 1'b1);
		prog_cycle_task(16'b0110000000011100, 1'b1);
		prog_cycle_task(16'b1110000000011100, 1'b1);
		prog_cycle_task(16'b0001000000011100, 1'b1);
		prog_cycle_task(16'b1001000000011100, 1'b1);
		prog_cycle_task(16'b0101000000011100, 1'b1);
		prog_cycle_task(16'b1101000000011100, 1'b1);
		prog_cycle_task(16'b0011000000011100, 1'b1);
		prog_cycle_task(16'b1011000000011100, 1'b1);
		prog_cycle_task(16'b0111000000011100, 1'b1);
		prog_cycle_task(16'b1111000000011100, 1'b1);
		prog_cycle_task(16'b0000100000011100, 1'b1);
		prog_cycle_task(16'b1000100000011100, 1'b1);
		prog_cycle_task(16'b0100100000011100, 1'b1);
		prog_cycle_task(16'b1100100000011100, 1'b1);
		prog_cycle_task(16'b0010100000011100, 1'b1);
		prog_cycle_task(16'b1010100000011100, 1'b1);
		prog_cycle_task(16'b0110100000011100, 1'b1);
		prog_cycle_task(16'b1110100000011100, 1'b1);
		prog_cycle_task(16'b0001100000011100, 1'b1);
		prog_cycle_task(16'b1001100000011100, 1'b1);
		prog_cycle_task(16'b0101100000011100, 1'b1);
		prog_cycle_task(16'b1101100000011100, 1'b1);
		prog_cycle_task(16'b0011100000011100, 1'b1);
		prog_cycle_task(16'b1011100000011100, 1'b1);
		prog_cycle_task(16'b0111100000011100, 1'b1);
		prog_cycle_task(16'b1111100000011100, 1'b1);
		prog_cycle_task(16'b0000010000011100, 1'b1);
		prog_cycle_task(16'b1000010000011100, 1'b1);
		prog_cycle_task(16'b0100010000011100, 1'b1);
		prog_cycle_task(16'b1100010000011100, 1'b1);
		prog_cycle_task(16'b0000000000111100, 1'b1);
		prog_cycle_task(16'b1000000000111100, 1'b0);
		prog_cycle_task(16'b0100000000111100, 1'b0);
		prog_cycle_task(16'b1100000000111100, 1'b1);
		prog_cycle_task(16'b0010000000111100, 1'b0);
		prog_cycle_task(16'b1010000000111100, 1'b0);
		prog_cycle_task(16'b0001000000111100, 1'b1);
		prog_cycle_task(16'b1001000000111100, 1'b1);
		prog_cycle_task(16'b0000100000111100, 1'b1);
		prog_cycle_task(16'b1000100000111100, 1'b0);
		prog_cycle_task(16'b0100100000111100, 1'b0);
		prog_cycle_task(16'b1100100000111100, 1'b1);
		prog_cycle_task(16'b0010100000111100, 1'b0);
		prog_cycle_task(16'b1010100000111100, 1'b0);
		prog_cycle_task(16'b0001100000111100, 1'b1);
		prog_cycle_task(16'b1001100000111100, 1'b0);
		prog_cycle_task(16'b0101100000111100, 1'b0);
		prog_cycle_task(16'b1101100000111100, 1'b1);
		prog_cycle_task(16'b0011100000111100, 1'b0);
		prog_cycle_task(16'b1011100000111100, 1'b0);
		prog_cycle_task(16'b0000010000111100, 1'b1);
		prog_cycle_task(16'b1000010000111100, 1'b0);
		prog_cycle_task(16'b0100010000111100, 1'b0);
		prog_cycle_task(16'b1100010000111100, 1'b1);
		prog_cycle_task(16'b0010010000111100, 1'b0);
		prog_cycle_task(16'b1010010000111100, 1'b0);
		prog_cycle_task(16'b0001010000111100, 1'b1);
		prog_cycle_task(16'b1001010000111100, 1'b0);
		prog_cycle_task(16'b0101010000111100, 1'b0);
		prog_cycle_task(16'b1101010000111100, 1'b1);
		prog_cycle_task(16'b0011010000111100, 1'b0);
		prog_cycle_task(16'b1011010000111100, 1'b0);
		prog_cycle_task(16'b0000110000111100, 1'b1);
		prog_cycle_task(16'b1000110000111100, 1'b0);
		prog_cycle_task(16'b0100110000111100, 1'b0);
		prog_cycle_task(16'b1100110000111100, 1'b1);
		prog_cycle_task(16'b0010110000111100, 1'b0);
		prog_cycle_task(16'b1010110000111100, 1'b0);
		prog_cycle_task(16'b0001110000111100, 1'b1);
		prog_cycle_task(16'b1001110000111100, 1'b0);
		prog_cycle_task(16'b0101110000111100, 1'b0);
		prog_cycle_task(16'b1101110000111100, 1'b1);
		prog_cycle_task(16'b0011110000111100, 1'b0);
		prog_cycle_task(16'b1011110000111100, 1'b0);
		prog_cycle_task(16'b0000001000111100, 1'b1);
		prog_cycle_task(16'b1000001000111100, 1'b0);
		prog_cycle_task(16'b0100001000111100, 1'b0);
		prog_cycle_task(16'b1100001000111100, 1'b1);
		prog_cycle_task(16'b0010001000111100, 1'b0);
		prog_cycle_task(16'b1010001000111100, 1'b0);
		prog_cycle_task(16'b0001001000111100, 1'b1);
		prog_cycle_task(16'b1001001000111100, 1'b0);
		prog_cycle_task(16'b0101001000111100, 1'b0);
		prog_cycle_task(16'b1101001000111100, 1'b1);
		prog_cycle_task(16'b0011001000111100, 1'b0);
		prog_cycle_task(16'b1011001000111100, 1'b0);
		prog_cycle_task(16'b0000000000000010, 1'b1);
		prog_cycle_task(16'b0100000000000010, 1'b1);
		prog_cycle_task(16'b0010000000000010, 1'b1);
		prog_cycle_task(16'b0110000000000010, 1'b1);
		prog_cycle_task(16'b0001000000000010, 1'b1);
		prog_cycle_task(16'b0101000000000010, 1'b1);
		prog_cycle_task(16'b0011000000000010, 1'b1);
		prog_cycle_task(16'b0111000000000010, 1'b1);
		prog_cycle_task(16'b0000000000100010, 1'b1);
		prog_cycle_task(16'b1000000000100010, 1'b0);
		prog_cycle_task(16'b0100000000100010, 1'b0);
		prog_cycle_task(16'b1100000000100010, 1'b1);
		prog_cycle_task(16'b0010000000100010, 1'b0);
		prog_cycle_task(16'b1010000000100010, 1'b0);
		prog_cycle_task(16'b0001000000100010, 1'b1);
		prog_cycle_task(16'b1001000000100010, 1'b1);
		prog_cycle_task(16'b0000100000100010, 1'b1);
		prog_cycle_task(16'b1000100000100010, 1'b1);
		prog_cycle_task(16'b0001100000100010, 1'b1);
		prog_cycle_task(16'b1001100000100010, 1'b1);
		prog_cycle_task(16'b0000010000100010, 1'b1);
		prog_cycle_task(16'b1000010000100010, 1'b0);
		prog_cycle_task(16'b0100010000100010, 1'b0);
		prog_cycle_task(16'b1100010000100010, 1'b1);
		prog_cycle_task(16'b0010010000100010, 1'b0);
		prog_cycle_task(16'b1010010000100010, 1'b0);
		prog_cycle_task(16'b0001010000100010, 1'b1);
		prog_cycle_task(16'b1001010000100010, 1'b0);
		prog_cycle_task(16'b0101010000100010, 1'b0);
		prog_cycle_task(16'b1101010000100010, 1'b1);
		prog_cycle_task(16'b0011010000100010, 1'b0);
		prog_cycle_task(16'b1011010000100010, 1'b0);
		prog_cycle_task(16'b0000110000100010, 1'b1);
		prog_cycle_task(16'b1000110000100010, 1'b0);
		prog_cycle_task(16'b0100110000100010, 1'b0);
		prog_cycle_task(16'b1100110000100010, 1'b1);
		prog_cycle_task(16'b0010110000100010, 1'b0);
		prog_cycle_task(16'b1010110000100010, 1'b0);
		prog_cycle_task(16'b0001110000100010, 1'b1);
		prog_cycle_task(16'b1001110000100010, 1'b0);
		prog_cycle_task(16'b0101110000100010, 1'b0);
		prog_cycle_task(16'b1101110000100010, 1'b1);
		prog_cycle_task(16'b0011110000100010, 1'b0);
		prog_cycle_task(16'b1011110000100010, 1'b0);
		prog_cycle_task(16'b0000001000100010, 1'b0);
		prog_cycle_task(16'b1000001000100010, 1'b1);
		prog_cycle_task(16'b0100001000100010, 1'b0);
		prog_cycle_task(16'b1100001000100010, 1'b1);
		prog_cycle_task(16'b0010001000100010, 1'b0);
		prog_cycle_task(16'b1010001000100010, 1'b0);
		prog_cycle_task(16'b0001001000100010, 1'b1);
		prog_cycle_task(16'b1001001000100010, 1'b0);
		prog_cycle_task(16'b0101001000100010, 1'b0);
		prog_cycle_task(16'b1101001000100010, 1'b1);
		prog_cycle_task(16'b0011001000100010, 1'b0);
		prog_cycle_task(16'b1011001000100010, 1'b0);
		prog_cycle_task(16'b0000101000100010, 1'b1);
		prog_cycle_task(16'b1000101000100010, 1'b0);
		prog_cycle_task(16'b0100101000100010, 1'b0);
		prog_cycle_task(16'b1100101000100010, 1'b1);
		prog_cycle_task(16'b0010101000100010, 1'b0);
		prog_cycle_task(16'b1010101000100010, 1'b0);
		prog_cycle_task(16'b0000000000010010, 1'b1);
		prog_cycle_task(16'b1000000000010010, 1'b0);
		prog_cycle_task(16'b0100000000010010, 1'b0);
		prog_cycle_task(16'b1100000000010010, 1'b1);
		prog_cycle_task(16'b0010000000010010, 1'b0);
		prog_cycle_task(16'b1010000000010010, 1'b0);
		prog_cycle_task(16'b0001000000010010, 1'b1);
		prog_cycle_task(16'b1001000000010010, 1'b1);
		prog_cycle_task(16'b0000100000010010, 1'b1);
		prog_cycle_task(16'b1000100000010010, 1'b0);
		prog_cycle_task(16'b0100100000010010, 1'b0);
		prog_cycle_task(16'b1100100000010010, 1'b1);
		prog_cycle_task(16'b0010100000010010, 1'b0);
		prog_cycle_task(16'b1010100000010010, 1'b0);
		prog_cycle_task(16'b0001100000010010, 1'b1);
		prog_cycle_task(16'b1001100000010010, 1'b0);
		prog_cycle_task(16'b0101100000010010, 1'b0);
		prog_cycle_task(16'b1101100000010010, 1'b1);
		prog_cycle_task(16'b0011100000010010, 1'b0);
		prog_cycle_task(16'b1011100000010010, 1'b0);
		prog_cycle_task(16'b0000010000010010, 1'b1);
		prog_cycle_task(16'b1000010000010010, 1'b0);
		prog_cycle_task(16'b0100010000010010, 1'b0);
		prog_cycle_task(16'b1100010000010010, 1'b1);
		prog_cycle_task(16'b0010010000010010, 1'b0);
		prog_cycle_task(16'b1010010000010010, 1'b0);
		prog_cycle_task(16'b0001010000010010, 1'b1);
		prog_cycle_task(16'b1001010000010010, 1'b0);
		prog_cycle_task(16'b0101010000010010, 1'b0);
		prog_cycle_task(16'b1101010000010010, 1'b1);
		prog_cycle_task(16'b0011010000010010, 1'b0);
		prog_cycle_task(16'b1011010000010010, 1'b0);
		prog_cycle_task(16'b0000110000010010, 1'b1);
		prog_cycle_task(16'b1000110000010010, 1'b0);
		prog_cycle_task(16'b0100110000010010, 1'b0);
		prog_cycle_task(16'b1100110000010010, 1'b1);
		prog_cycle_task(16'b0010110000010010, 1'b0);
		prog_cycle_task(16'b1010110000010010, 1'b0);
		prog_cycle_task(16'b0001110000010010, 1'b1);
		prog_cycle_task(16'b1001110000010010, 1'b0);
		prog_cycle_task(16'b0101110000010010, 1'b0);
		prog_cycle_task(16'b1101110000010010, 1'b1);
		prog_cycle_task(16'b0011110000010010, 1'b0);
		prog_cycle_task(16'b1011110000010010, 1'b0);
		prog_cycle_task(16'b0000001000010010, 1'b1);
		prog_cycle_task(16'b1000001000010010, 1'b0);
		prog_cycle_task(16'b0100001000010010, 1'b0);
		prog_cycle_task(16'b1100001000010010, 1'b1);
		prog_cycle_task(16'b0010001000010010, 1'b0);
		prog_cycle_task(16'b1010001000010010, 1'b0);
		prog_cycle_task(16'b0001001000010010, 1'b1);
		prog_cycle_task(16'b1001001000010010, 1'b0);
		prog_cycle_task(16'b0101001000010010, 1'b0);
		prog_cycle_task(16'b1101001000010010, 1'b1);
		prog_cycle_task(16'b0011001000010010, 1'b0);
		prog_cycle_task(16'b1011001000010010, 1'b0);
		prog_cycle_task(16'b0000101000010010, 1'b1);
		prog_cycle_task(16'b1000101000010010, 1'b0);
		prog_cycle_task(16'b0100101000010010, 1'b0);
		prog_cycle_task(16'b1100101000010010, 1'b1);
		prog_cycle_task(16'b0010101000010010, 1'b0);
		prog_cycle_task(16'b1010101000010010, 1'b0);
		prog_cycle_task(16'b0000000000110010, 1'b1);
		prog_cycle_task(16'b1000000000110010, 1'b0);
		prog_cycle_task(16'b0100000000110010, 1'b0);
		prog_cycle_task(16'b1100000000110010, 1'b1);
		prog_cycle_task(16'b0010000000110010, 1'b0);
		prog_cycle_task(16'b1010000000110010, 1'b0);
		prog_cycle_task(16'b0001000000110010, 1'b1);
		prog_cycle_task(16'b1001000000110010, 1'b1);
		prog_cycle_task(16'b0000100000110010, 1'b1);
		prog_cycle_task(16'b1000100000110010, 1'b0);
		prog_cycle_task(16'b0100100000110010, 1'b0);
		prog_cycle_task(16'b1100100000110010, 1'b1);
		prog_cycle_task(16'b0010100000110010, 1'b0);
		prog_cycle_task(16'b1010100000110010, 1'b0);
		prog_cycle_task(16'b0001100000110010, 1'b1);
		prog_cycle_task(16'b1001100000110010, 1'b1);
		prog_cycle_task(16'b0000010000110010, 1'b1);
		prog_cycle_task(16'b1000010000110010, 1'b1);
		prog_cycle_task(16'b0000000000001010, 1'b0);
		prog_cycle_task(16'b1000000000001010, 1'b0);
		prog_cycle_task(16'b0100000000001010, 1'b0);
		prog_cycle_task(16'b1100000000001010, 1'b0);
		prog_cycle_task(16'b0010000000001010, 1'b0);
		prog_cycle_task(16'b1010000000001010, 1'b0);
		prog_cycle_task(16'b0110000000001010, 1'b0);
		prog_cycle_task(16'b1110000000001010, 1'b0);
		prog_cycle_task(16'b0001000000001010, 1'b0);
		prog_cycle_task(16'b1001000000001010, 1'b0);
		prog_cycle_task(16'b0101000000001010, 1'b0);
		prog_cycle_task(16'b1101000000001010, 1'b0);
		prog_cycle_task(16'b0011000000001010, 1'b0);
		prog_cycle_task(16'b1011000000001010, 1'b0);
		prog_cycle_task(16'b0111000000001010, 1'b0);
		prog_cycle_task(16'b1111000000001010, 1'b0);
		prog_cycle_task(16'b0000100000001010, 1'b0);
		prog_cycle_task(16'b1000100000001010, 1'b0);
		prog_cycle_task(16'b0100100000001010, 1'b1);
		prog_cycle_task(16'b0000010000001010, 1'b0);
		prog_cycle_task(16'b1000010000001010, 1'b0);
		prog_cycle_task(16'b0100010000001010, 1'b0);
		prog_cycle_task(16'b1100010000001010, 1'b0);
		prog_cycle_task(16'b0010010000001010, 1'b0);
		prog_cycle_task(16'b1010010000001010, 1'b0);
		prog_cycle_task(16'b0110010000001010, 1'b0);
		prog_cycle_task(16'b1110010000001010, 1'b0);
		prog_cycle_task(16'b0001010000001010, 1'b0);
		prog_cycle_task(16'b1001010000001010, 1'b0);
		prog_cycle_task(16'b0101010000001010, 1'b0);
		prog_cycle_task(16'b1101010000001010, 1'b0);
		prog_cycle_task(16'b0011010000001010, 1'b0);
		prog_cycle_task(16'b1011010000001010, 1'b0);
		prog_cycle_task(16'b0111010000001010, 1'b0);
		prog_cycle_task(16'b1111010000001010, 1'b0);
		prog_cycle_task(16'b0000110000001010, 1'b0);
		prog_cycle_task(16'b1000110000001010, 1'b0);
		prog_cycle_task(16'b0100110000001010, 1'b1);
		prog_cycle_task(16'b0000001000001010, 1'b0);
		prog_cycle_task(16'b1000001000001010, 1'b0);
		prog_cycle_task(16'b0100001000001010, 1'b0);
		prog_cycle_task(16'b1100001000001010, 1'b0);
		prog_cycle_task(16'b0010001000001010, 1'b0);
		prog_cycle_task(16'b1010001000001010, 1'b0);
		prog_cycle_task(16'b0110001000001010, 1'b0);
		prog_cycle_task(16'b1110001000001010, 1'b0);
		prog_cycle_task(16'b0001001000001010, 1'b0);
		prog_cycle_task(16'b1001001000001010, 1'b0);
		prog_cycle_task(16'b0101001000001010, 1'b0);
		prog_cycle_task(16'b1101001000001010, 1'b0);
		prog_cycle_task(16'b0011001000001010, 1'b0);
		prog_cycle_task(16'b1011001000001010, 1'b0);
		prog_cycle_task(16'b0111001000001010, 1'b0);
		prog_cycle_task(16'b1111001000001010, 1'b0);
		prog_cycle_task(16'b0000101000001010, 1'b0);
		prog_cycle_task(16'b1000101000001010, 1'b0);
		prog_cycle_task(16'b0100101000001010, 1'b1);
		prog_cycle_task(16'b0000011000001010, 1'b0);
		prog_cycle_task(16'b1000011000001010, 1'b0);
		prog_cycle_task(16'b0100011000001010, 1'b0);
		prog_cycle_task(16'b1100011000001010, 1'b0);
		prog_cycle_task(16'b0010011000001010, 1'b0);
		prog_cycle_task(16'b1010011000001010, 1'b0);
		prog_cycle_task(16'b0110011000001010, 1'b0);
		prog_cycle_task(16'b1110011000001010, 1'b0);
		prog_cycle_task(16'b0001011000001010, 1'b0);
		prog_cycle_task(16'b1001011000001010, 1'b0);
		prog_cycle_task(16'b0101011000001010, 1'b0);
		prog_cycle_task(16'b1101011000001010, 1'b0);
		prog_cycle_task(16'b0011011000001010, 1'b0);
		prog_cycle_task(16'b1011011000001010, 1'b0);
		prog_cycle_task(16'b0111011000001010, 1'b0);
		prog_cycle_task(16'b1111011000001010, 1'b0);
		prog_cycle_task(16'b0000111000001010, 1'b0);
		prog_cycle_task(16'b1000111000001010, 1'b0);
		prog_cycle_task(16'b0100111000001010, 1'b1);
		prog_cycle_task(16'b0000000100001010, 1'b0);
		prog_cycle_task(16'b1000000100001010, 1'b0);
		prog_cycle_task(16'b0100000100001010, 1'b1);
		prog_cycle_task(16'b1100000100001010, 1'b0);
		prog_cycle_task(16'b0010000100001010, 1'b0);
		prog_cycle_task(16'b1010000100001010, 1'b0);
		prog_cycle_task(16'b0110000100001010, 1'b0);
		prog_cycle_task(16'b1110000100001010, 1'b1);
		prog_cycle_task(16'b0000010100001010, 1'b0);
		prog_cycle_task(16'b1000010100001010, 1'b0);
		prog_cycle_task(16'b0100010100001010, 1'b1);
		prog_cycle_task(16'b1100010100001010, 1'b0);
		prog_cycle_task(16'b0010010100001010, 1'b0);
		prog_cycle_task(16'b1010010100001010, 1'b0);
		prog_cycle_task(16'b0110010100001010, 1'b0);
		prog_cycle_task(16'b1110010100001010, 1'b1);
		prog_cycle_task(16'b0000001100001010, 1'b0);
		prog_cycle_task(16'b1000001100001010, 1'b0);
		prog_cycle_task(16'b0100001100001010, 1'b1);
		prog_cycle_task(16'b1100001100001010, 1'b0);
		prog_cycle_task(16'b0010001100001010, 1'b0);
		prog_cycle_task(16'b1010001100001010, 1'b0);
		prog_cycle_task(16'b0110001100001010, 1'b0);
		prog_cycle_task(16'b1110001100001010, 1'b1);
		prog_cycle_task(16'b0000011100001010, 1'b0);
		prog_cycle_task(16'b1000011100001010, 1'b0);
		prog_cycle_task(16'b0100011100001010, 1'b1);
		prog_cycle_task(16'b1100011100001010, 1'b0);
		prog_cycle_task(16'b0010011100001010, 1'b0);
		prog_cycle_task(16'b1010011100001010, 1'b0);
		prog_cycle_task(16'b0110011100001010, 1'b0);
		prog_cycle_task(16'b1110011100001010, 1'b1);
		prog_cycle_task(16'b0000000010001010, 1'b0);
		prog_cycle_task(16'b1000000010001010, 1'b0);
		prog_cycle_task(16'b0100000010001010, 1'b1);
		prog_cycle_task(16'b1100000010001010, 1'b0);
		prog_cycle_task(16'b0010000010001010, 1'b0);
		prog_cycle_task(16'b1010000010001010, 1'b0);
		prog_cycle_task(16'b0110000010001010, 1'b0);
		prog_cycle_task(16'b1110000010001010, 1'b1);
		prog_cycle_task(16'b0000010010001010, 1'b0);
		prog_cycle_task(16'b1000010010001010, 1'b0);
		prog_cycle_task(16'b0100010010001010, 1'b1);
		prog_cycle_task(16'b1100010010001010, 1'b0);
		prog_cycle_task(16'b0010010010001010, 1'b0);
		prog_cycle_task(16'b1010010010001010, 1'b0);
		prog_cycle_task(16'b0110010010001010, 1'b0);
		prog_cycle_task(16'b1110010010001010, 1'b1);
		prog_cycle_task(16'b0000001010001010, 1'b0);
		prog_cycle_task(16'b1000001010001010, 1'b0);
		prog_cycle_task(16'b0100001010001010, 1'b1);
		prog_cycle_task(16'b1100001010001010, 1'b0);
		prog_cycle_task(16'b0010001010001010, 1'b0);
		prog_cycle_task(16'b1010001010001010, 1'b0);
		prog_cycle_task(16'b0110001010001010, 1'b0);
		prog_cycle_task(16'b1110001010001010, 1'b1);
		prog_cycle_task(16'b0000011010001010, 1'b0);
		prog_cycle_task(16'b1000011010001010, 1'b0);
		prog_cycle_task(16'b0100011010001010, 1'b1);
		prog_cycle_task(16'b1100011010001010, 1'b0);
		prog_cycle_task(16'b0010011010001010, 1'b0);
		prog_cycle_task(16'b1010011010001010, 1'b0);
		prog_cycle_task(16'b0110011010001010, 1'b0);
		prog_cycle_task(16'b1110011010001010, 1'b1);
		prog_cycle_task(16'b0000000110001010, 1'b0);
		prog_cycle_task(16'b1000000110001010, 1'b0);
		prog_cycle_task(16'b0100000110001010, 1'b1);
		prog_cycle_task(16'b1100000110001010, 1'b0);
		prog_cycle_task(16'b0010000110001010, 1'b0);
		prog_cycle_task(16'b1010000110001010, 1'b0);
		prog_cycle_task(16'b0110000110001010, 1'b0);
		prog_cycle_task(16'b1110000110001010, 1'b1);
		prog_cycle_task(16'b0000010110001010, 1'b0);
		prog_cycle_task(16'b1000010110001010, 1'b0);
		prog_cycle_task(16'b0100010110001010, 1'b1);
		prog_cycle_task(16'b1100010110001010, 1'b0);
		prog_cycle_task(16'b0010010110001010, 1'b0);
		prog_cycle_task(16'b1010010110001010, 1'b0);
		prog_cycle_task(16'b0110010110001010, 1'b0);
		prog_cycle_task(16'b1110010110001010, 1'b1);
		prog_cycle_task(16'b0000001110001010, 1'b0);
		prog_cycle_task(16'b1000001110001010, 1'b0);
		prog_cycle_task(16'b0100001110001010, 1'b1);
		prog_cycle_task(16'b1100001110001010, 1'b0);
		prog_cycle_task(16'b0010001110001010, 1'b0);
		prog_cycle_task(16'b1010001110001010, 1'b0);
		prog_cycle_task(16'b0110001110001010, 1'b0);
		prog_cycle_task(16'b1110001110001010, 1'b1);
		prog_cycle_task(16'b0000011110001010, 1'b0);
		prog_cycle_task(16'b1000011110001010, 1'b0);
		prog_cycle_task(16'b0100011110001010, 1'b1);
		prog_cycle_task(16'b1100011110001010, 1'b0);
		prog_cycle_task(16'b0010011110001010, 1'b0);
		prog_cycle_task(16'b1010011110001010, 1'b0);
		prog_cycle_task(16'b0110011110001010, 1'b0);
		prog_cycle_task(16'b1110011110001010, 1'b1);
		prog_cycle_task(16'b0000000001001010, 1'b0);
		prog_cycle_task(16'b1000000001001010, 1'b0);
		prog_cycle_task(16'b0100000001001010, 1'b1);
		prog_cycle_task(16'b1100000001001010, 1'b0);
		prog_cycle_task(16'b0010000001001010, 1'b0);
		prog_cycle_task(16'b1010000001001010, 1'b0);
		prog_cycle_task(16'b0110000001001010, 1'b0);
		prog_cycle_task(16'b1110000001001010, 1'b1);
		prog_cycle_task(16'b0000010001001010, 1'b0);
		prog_cycle_task(16'b1000010001001010, 1'b0);
		prog_cycle_task(16'b0100010001001010, 1'b1);
		prog_cycle_task(16'b1100010001001010, 1'b0);
		prog_cycle_task(16'b0010010001001010, 1'b0);
		prog_cycle_task(16'b1010010001001010, 1'b0);
		prog_cycle_task(16'b0110010001001010, 1'b0);
		prog_cycle_task(16'b1110010001001010, 1'b1);
		prog_cycle_task(16'b0000001001001010, 1'b0);
		prog_cycle_task(16'b1000001001001010, 1'b0);
		prog_cycle_task(16'b0100001001001010, 1'b1);
		prog_cycle_task(16'b1100001001001010, 1'b0);
		prog_cycle_task(16'b0010001001001010, 1'b0);
		prog_cycle_task(16'b1010001001001010, 1'b0);
		prog_cycle_task(16'b0110001001001010, 1'b0);
		prog_cycle_task(16'b1110001001001010, 1'b1);
		prog_cycle_task(16'b0000011001001010, 1'b0);
		prog_cycle_task(16'b1000011001001010, 1'b0);
		prog_cycle_task(16'b0100011001001010, 1'b1);
		prog_cycle_task(16'b1100011001001010, 1'b0);
		prog_cycle_task(16'b0010011001001010, 1'b0);
		prog_cycle_task(16'b1010011001001010, 1'b0);
		prog_cycle_task(16'b0110011001001010, 1'b0);
		prog_cycle_task(16'b1110011001001010, 1'b1);
		prog_cycle_task(16'b0000000000101010, 1'b1);
		prog_cycle_task(16'b1000000000101010, 1'b1);
		prog_cycle_task(16'b0100000000101010, 1'b1);
		prog_cycle_task(16'b1100000000101010, 1'b1);
		prog_cycle_task(16'b0010000000101010, 1'b1);
		prog_cycle_task(16'b1010000000101010, 1'b1);
		prog_cycle_task(16'b0110000000101010, 1'b1);
		prog_cycle_task(16'b1110000000101010, 1'b1);
		prog_cycle_task(16'b0001000000101010, 1'b1);
		prog_cycle_task(16'b1001000000101010, 1'b1);
		prog_cycle_task(16'b0101000000101010, 1'b1);
		prog_cycle_task(16'b1101000000101010, 1'b1);
		prog_cycle_task(16'b0011000000101010, 1'b1);
		prog_cycle_task(16'b1011000000101010, 1'b1);
		prog_cycle_task(16'b0111000000101010, 1'b1);
		prog_cycle_task(16'b1111000000101010, 1'b1);
		prog_cycle_task(16'b0000100000101010, 1'b1);
		prog_cycle_task(16'b1000100000101010, 1'b1);
		prog_cycle_task(16'b0100100000101010, 1'b1);
		prog_cycle_task(16'b1100100000101010, 1'b1);
		prog_cycle_task(16'b0010100000101010, 1'b0);
		prog_cycle_task(16'b1010100000101010, 1'b1);
		prog_cycle_task(16'b0110100000101010, 1'b1);
		prog_cycle_task(16'b1110100000101010, 1'b1);
		prog_cycle_task(16'b0001100000101010, 1'b1);
		prog_cycle_task(16'b1001100000101010, 1'b1);
		prog_cycle_task(16'b0101100000101010, 1'b1);
		prog_cycle_task(16'b1101100000101010, 1'b1);
		prog_cycle_task(16'b0011100000101010, 1'b1);
		prog_cycle_task(16'b1011100000101010, 1'b1);
		prog_cycle_task(16'b0111100000101010, 1'b1);
		prog_cycle_task(16'b1111100000101010, 1'b1);
		prog_cycle_task(16'b0000010000101010, 1'b1);
		prog_cycle_task(16'b1000010000101010, 1'b1);
		prog_cycle_task(16'b0100010000101010, 1'b1);
		prog_cycle_task(16'b1100010000101010, 1'b1);
		prog_cycle_task(16'b0000000000011010, 1'b1);
		prog_cycle_task(16'b1000000000011010, 1'b0);
		prog_cycle_task(16'b0100000000011010, 1'b0);
		prog_cycle_task(16'b1100000000011010, 1'b1);
		prog_cycle_task(16'b0010000000011010, 1'b0);
		prog_cycle_task(16'b1010000000011010, 1'b0);
		prog_cycle_task(16'b0001000000011010, 1'b0);
		prog_cycle_task(16'b1001000000011010, 1'b1);
		prog_cycle_task(16'b0000100000011010, 1'b1);
		prog_cycle_task(16'b1000100000011010, 1'b0);
		prog_cycle_task(16'b0100100000011010, 1'b0);
		prog_cycle_task(16'b1100100000011010, 1'b1);
		prog_cycle_task(16'b0010100000011010, 1'b0);
		prog_cycle_task(16'b1010100000011010, 1'b0);
		prog_cycle_task(16'b0001100000011010, 1'b1);
		prog_cycle_task(16'b1001100000011010, 1'b0);
		prog_cycle_task(16'b0101100000011010, 1'b0);
		prog_cycle_task(16'b1101100000011010, 1'b1);
		prog_cycle_task(16'b0011100000011010, 1'b0);
		prog_cycle_task(16'b1011100000011010, 1'b0);
		prog_cycle_task(16'b0000010000011010, 1'b1);
		prog_cycle_task(16'b1000010000011010, 1'b0);
		prog_cycle_task(16'b0100010000011010, 1'b0);
		prog_cycle_task(16'b1100010000011010, 1'b1);
		prog_cycle_task(16'b0010010000011010, 1'b0);
		prog_cycle_task(16'b1010010000011010, 1'b0);
		prog_cycle_task(16'b0001010000011010, 1'b1);
		prog_cycle_task(16'b1001010000011010, 1'b0);
		prog_cycle_task(16'b0101010000011010, 1'b0);
		prog_cycle_task(16'b1101010000011010, 1'b1);
		prog_cycle_task(16'b0011010000011010, 1'b0);
		prog_cycle_task(16'b1011010000011010, 1'b0);
		prog_cycle_task(16'b0000110000011010, 1'b1);
		prog_cycle_task(16'b1000110000011010, 1'b0);
		prog_cycle_task(16'b0100110000011010, 1'b0);
		prog_cycle_task(16'b1100110000011010, 1'b1);
		prog_cycle_task(16'b0010110000011010, 1'b0);
		prog_cycle_task(16'b1010110000011010, 1'b0);
		prog_cycle_task(16'b0001110000011010, 1'b1);
		prog_cycle_task(16'b1001110000011010, 1'b0);
		prog_cycle_task(16'b0101110000011010, 1'b0);
		prog_cycle_task(16'b1101110000011010, 1'b1);
		prog_cycle_task(16'b0011110000011010, 1'b0);
		prog_cycle_task(16'b1011110000011010, 1'b0);
		prog_cycle_task(16'b0000001000011010, 1'b1);
		prog_cycle_task(16'b1000001000011010, 1'b0);
		prog_cycle_task(16'b0100001000011010, 1'b0);
		prog_cycle_task(16'b1100001000011010, 1'b1);
		prog_cycle_task(16'b0010001000011010, 1'b0);
		prog_cycle_task(16'b1010001000011010, 1'b0);
		prog_cycle_task(16'b0001001000011010, 1'b0);
		prog_cycle_task(16'b1001001000011010, 1'b0);
		prog_cycle_task(16'b0101001000011010, 1'b1);
		prog_cycle_task(16'b1101001000011010, 1'b1);
		prog_cycle_task(16'b0011001000011010, 1'b0);
		prog_cycle_task(16'b1011001000011010, 1'b0);
		prog_cycle_task(16'b0000101000011010, 1'b1);
		prog_cycle_task(16'b1000101000011010, 1'b0);
		prog_cycle_task(16'b0100101000011010, 1'b0);
		prog_cycle_task(16'b1100101000011010, 1'b1);
		prog_cycle_task(16'b0010101000011010, 1'b0);
		prog_cycle_task(16'b1010101000011010, 1'b0);
		prog_cycle_task(16'b0000000000111010, 1'b0);
		prog_cycle_task(16'b1000000000111010, 1'b1);
		prog_cycle_task(16'b0100000000111010, 1'b0);
		prog_cycle_task(16'b1100000000111010, 1'b1);
		prog_cycle_task(16'b0010000000111010, 1'b0);
		prog_cycle_task(16'b1010000000111010, 1'b0);
		prog_cycle_task(16'b0001000000111010, 1'b0);
		prog_cycle_task(16'b1001000000111010, 1'b1);
		prog_cycle_task(16'b0101000000111010, 1'b0);
		prog_cycle_task(16'b1101000000111010, 1'b1);
		prog_cycle_task(16'b0011000000111010, 1'b0);
		prog_cycle_task(16'b1011000000111010, 1'b0);
		prog_cycle_task(16'b0000100000111010, 1'b1);
		prog_cycle_task(16'b1000100000111010, 1'b0);
		prog_cycle_task(16'b0100100000111010, 1'b0);
		prog_cycle_task(16'b1100100000111010, 1'b1);
		prog_cycle_task(16'b0010100000111010, 1'b0);
		prog_cycle_task(16'b1010100000111010, 1'b0);
		prog_cycle_task(16'b0001100000111010, 1'b0);
		prog_cycle_task(16'b1001100000111010, 1'b1);
		prog_cycle_task(16'b0101100000111010, 1'b0);
		prog_cycle_task(16'b1101100000111010, 1'b1);
		prog_cycle_task(16'b0011100000111010, 1'b0);
		prog_cycle_task(16'b1011100000111010, 1'b0);
		prog_cycle_task(16'b0000010000111010, 1'b1);
		prog_cycle_task(16'b1000010000111010, 1'b0);
		prog_cycle_task(16'b0100010000111010, 1'b0);
		prog_cycle_task(16'b1100010000111010, 1'b1);
		prog_cycle_task(16'b0010010000111010, 1'b0);
		prog_cycle_task(16'b1010010000111010, 1'b0);
		prog_cycle_task(16'b0001010000111010, 1'b0);
		prog_cycle_task(16'b1001010000111010, 1'b1);
		prog_cycle_task(16'b0101010000111010, 1'b0);
		prog_cycle_task(16'b1101010000111010, 1'b1);
		prog_cycle_task(16'b0011010000111010, 1'b0);
		prog_cycle_task(16'b1011010000111010, 1'b0);
		prog_cycle_task(16'b0000110000111010, 1'b1);
		prog_cycle_task(16'b1000110000111010, 1'b0);
		prog_cycle_task(16'b0100110000111010, 1'b0);
		prog_cycle_task(16'b1100110000111010, 1'b1);
		prog_cycle_task(16'b0010110000111010, 1'b0);
		prog_cycle_task(16'b1010110000111010, 1'b0);
		prog_cycle_task(16'b0001110000111010, 1'b0);
		prog_cycle_task(16'b1001110000111010, 1'b1);
		prog_cycle_task(16'b0101110000111010, 1'b0);
		prog_cycle_task(16'b1101110000111010, 1'b1);
		prog_cycle_task(16'b0011110000111010, 1'b0);
		prog_cycle_task(16'b1011110000111010, 1'b0);
		prog_cycle_task(16'b0000001000111010, 1'b1);
		prog_cycle_task(16'b1000001000111010, 1'b0);
		prog_cycle_task(16'b0100001000111010, 1'b0);
		prog_cycle_task(16'b1100001000111010, 1'b1);
		prog_cycle_task(16'b0010001000111010, 1'b0);
		prog_cycle_task(16'b1010001000111010, 1'b0);
		prog_cycle_task(16'b0001001000111010, 1'b0);
		prog_cycle_task(16'b1001001000111010, 1'b1);
		prog_cycle_task(16'b0000101000111010, 1'b1);
		prog_cycle_task(16'b1000101000111010, 1'b1);
		prog_cycle_task(16'b0000000000000110, 1'b0);
		prog_cycle_task(16'b1000000000000110, 1'b0);
		prog_cycle_task(16'b0100000000000110, 1'b0);
		prog_cycle_task(16'b1100000000000110, 1'b0);
		prog_cycle_task(16'b0010000000000110, 1'b0);
		prog_cycle_task(16'b1010000000000110, 1'b0);
		prog_cycle_task(16'b0110000000000110, 1'b0);
		prog_cycle_task(16'b1110000000000110, 1'b0);
		prog_cycle_task(16'b0001000000000110, 1'b0);
		prog_cycle_task(16'b1001000000000110, 1'b0);
		prog_cycle_task(16'b0101000000000110, 1'b0);
		prog_cycle_task(16'b1101000000000110, 1'b0);
		prog_cycle_task(16'b0011000000000110, 1'b0);
		prog_cycle_task(16'b1011000000000110, 1'b0);
		prog_cycle_task(16'b0111000000000110, 1'b0);
		prog_cycle_task(16'b1111000000000110, 1'b0);
		prog_cycle_task(16'b0000100000000110, 1'b0);
		prog_cycle_task(16'b1000100000000110, 1'b0);
		prog_cycle_task(16'b0100100000000110, 1'b1);
		prog_cycle_task(16'b0000010000000110, 1'b0);
		prog_cycle_task(16'b1000010000000110, 1'b0);
		prog_cycle_task(16'b0100010000000110, 1'b0);
		prog_cycle_task(16'b1100010000000110, 1'b0);
		prog_cycle_task(16'b0010010000000110, 1'b0);
		prog_cycle_task(16'b1010010000000110, 1'b0);
		prog_cycle_task(16'b0110010000000110, 1'b0);
		prog_cycle_task(16'b1110010000000110, 1'b0);
		prog_cycle_task(16'b0001010000000110, 1'b0);
		prog_cycle_task(16'b1001010000000110, 1'b0);
		prog_cycle_task(16'b0101010000000110, 1'b0);
		prog_cycle_task(16'b1101010000000110, 1'b0);
		prog_cycle_task(16'b0011010000000110, 1'b0);
		prog_cycle_task(16'b1011010000000110, 1'b0);
		prog_cycle_task(16'b0111010000000110, 1'b0);
		prog_cycle_task(16'b1111010000000110, 1'b0);
		prog_cycle_task(16'b0000110000000110, 1'b0);
		prog_cycle_task(16'b1000110000000110, 1'b0);
		prog_cycle_task(16'b0100110000000110, 1'b1);
		prog_cycle_task(16'b0000001000000110, 1'b0);
		prog_cycle_task(16'b1000001000000110, 1'b0);
		prog_cycle_task(16'b0100001000000110, 1'b0);
		prog_cycle_task(16'b1100001000000110, 1'b0);
		prog_cycle_task(16'b0010001000000110, 1'b0);
		prog_cycle_task(16'b1010001000000110, 1'b0);
		prog_cycle_task(16'b0110001000000110, 1'b0);
		prog_cycle_task(16'b1110001000000110, 1'b0);
		prog_cycle_task(16'b0001001000000110, 1'b0);
		prog_cycle_task(16'b1001001000000110, 1'b0);
		prog_cycle_task(16'b0101001000000110, 1'b0);
		prog_cycle_task(16'b1101001000000110, 1'b0);
		prog_cycle_task(16'b0011001000000110, 1'b0);
		prog_cycle_task(16'b1011001000000110, 1'b0);
		prog_cycle_task(16'b0111001000000110, 1'b0);
		prog_cycle_task(16'b1111001000000110, 1'b0);
		prog_cycle_task(16'b0000101000000110, 1'b0);
		prog_cycle_task(16'b1000101000000110, 1'b0);
		prog_cycle_task(16'b0100101000000110, 1'b1);
		prog_cycle_task(16'b0000011000000110, 1'b1);
		prog_cycle_task(16'b1000011000000110, 1'b0);
		prog_cycle_task(16'b0100011000000110, 1'b1);
		prog_cycle_task(16'b1100011000000110, 1'b0);
		prog_cycle_task(16'b0010011000000110, 1'b1);
		prog_cycle_task(16'b1010011000000110, 1'b0);
		prog_cycle_task(16'b0110011000000110, 1'b1);
		prog_cycle_task(16'b1110011000000110, 1'b0);
		prog_cycle_task(16'b0001011000000110, 1'b0);
		prog_cycle_task(16'b1001011000000110, 1'b0);
		prog_cycle_task(16'b0101011000000110, 1'b0);
		prog_cycle_task(16'b1101011000000110, 1'b0);
		prog_cycle_task(16'b0011011000000110, 1'b0);
		prog_cycle_task(16'b1011011000000110, 1'b0);
		prog_cycle_task(16'b0111011000000110, 1'b0);
		prog_cycle_task(16'b1111011000000110, 1'b0);
		prog_cycle_task(16'b0000111000000110, 1'b0);
		prog_cycle_task(16'b1000111000000110, 1'b1);
		prog_cycle_task(16'b0100111000000110, 1'b0);
		prog_cycle_task(16'b0000000100000110, 1'b0);
		prog_cycle_task(16'b1000000100000110, 1'b0);
		prog_cycle_task(16'b0100000100000110, 1'b1);
		prog_cycle_task(16'b1100000100000110, 1'b0);
		prog_cycle_task(16'b0010000100000110, 1'b0);
		prog_cycle_task(16'b1010000100000110, 1'b0);
		prog_cycle_task(16'b0110000100000110, 1'b0);
		prog_cycle_task(16'b1110000100000110, 1'b1);
		prog_cycle_task(16'b0000010100000110, 1'b0);
		prog_cycle_task(16'b1000010100000110, 1'b0);
		prog_cycle_task(16'b0100010100000110, 1'b1);
		prog_cycle_task(16'b1100010100000110, 1'b0);
		prog_cycle_task(16'b0010010100000110, 1'b0);
		prog_cycle_task(16'b1010010100000110, 1'b0);
		prog_cycle_task(16'b0110010100000110, 1'b0);
		prog_cycle_task(16'b1110010100000110, 1'b1);
		prog_cycle_task(16'b0000001100000110, 1'b0);
		prog_cycle_task(16'b1000001100000110, 1'b0);
		prog_cycle_task(16'b0100001100000110, 1'b1);
		prog_cycle_task(16'b1100001100000110, 1'b0);
		prog_cycle_task(16'b0010001100000110, 1'b0);
		prog_cycle_task(16'b1010001100000110, 1'b0);
		prog_cycle_task(16'b0110001100000110, 1'b0);
		prog_cycle_task(16'b1110001100000110, 1'b1);
		prog_cycle_task(16'b0000011100000110, 1'b0);
		prog_cycle_task(16'b1000011100000110, 1'b0);
		prog_cycle_task(16'b0100011100000110, 1'b1);
		prog_cycle_task(16'b1100011100000110, 1'b0);
		prog_cycle_task(16'b0010011100000110, 1'b0);
		prog_cycle_task(16'b1010011100000110, 1'b0);
		prog_cycle_task(16'b0110011100000110, 1'b0);
		prog_cycle_task(16'b1110011100000110, 1'b1);
		prog_cycle_task(16'b0000000010000110, 1'b0);
		prog_cycle_task(16'b1000000010000110, 1'b0);
		prog_cycle_task(16'b0100000010000110, 1'b1);
		prog_cycle_task(16'b1100000010000110, 1'b0);
		prog_cycle_task(16'b0010000010000110, 1'b0);
		prog_cycle_task(16'b1010000010000110, 1'b0);
		prog_cycle_task(16'b0110000010000110, 1'b0);
		prog_cycle_task(16'b1110000010000110, 1'b1);
		prog_cycle_task(16'b0000010010000110, 1'b0);
		prog_cycle_task(16'b1000010010000110, 1'b0);
		prog_cycle_task(16'b0100010010000110, 1'b1);
		prog_cycle_task(16'b1100010010000110, 1'b0);
		prog_cycle_task(16'b0010010010000110, 1'b0);
		prog_cycle_task(16'b1010010010000110, 1'b0);
		prog_cycle_task(16'b0110010010000110, 1'b0);
		prog_cycle_task(16'b1110010010000110, 1'b1);
		prog_cycle_task(16'b0000001010000110, 1'b0);
		prog_cycle_task(16'b1000001010000110, 1'b0);
		prog_cycle_task(16'b0100001010000110, 1'b1);
		prog_cycle_task(16'b1100001010000110, 1'b0);
		prog_cycle_task(16'b0010001010000110, 1'b0);
		prog_cycle_task(16'b1010001010000110, 1'b0);
		prog_cycle_task(16'b0110001010000110, 1'b0);
		prog_cycle_task(16'b1110001010000110, 1'b1);
		prog_cycle_task(16'b0000011010000110, 1'b0);
		prog_cycle_task(16'b1000011010000110, 1'b0);
		prog_cycle_task(16'b0100011010000110, 1'b1);
		prog_cycle_task(16'b1100011010000110, 1'b0);
		prog_cycle_task(16'b0010011010000110, 1'b0);
		prog_cycle_task(16'b1010011010000110, 1'b0);
		prog_cycle_task(16'b0110011010000110, 1'b0);
		prog_cycle_task(16'b1110011010000110, 1'b1);
		prog_cycle_task(16'b0000000110000110, 1'b0);
		prog_cycle_task(16'b1000000110000110, 1'b0);
		prog_cycle_task(16'b0100000110000110, 1'b1);
		prog_cycle_task(16'b1100000110000110, 1'b0);
		prog_cycle_task(16'b0010000110000110, 1'b0);
		prog_cycle_task(16'b1010000110000110, 1'b0);
		prog_cycle_task(16'b0110000110000110, 1'b0);
		prog_cycle_task(16'b1110000110000110, 1'b1);
		prog_cycle_task(16'b0000010110000110, 1'b0);
		prog_cycle_task(16'b1000010110000110, 1'b0);
		prog_cycle_task(16'b0100010110000110, 1'b1);
		prog_cycle_task(16'b1100010110000110, 1'b0);
		prog_cycle_task(16'b0010010110000110, 1'b0);
		prog_cycle_task(16'b1010010110000110, 1'b0);
		prog_cycle_task(16'b0110010110000110, 1'b0);
		prog_cycle_task(16'b1110010110000110, 1'b1);
		prog_cycle_task(16'b0000001110000110, 1'b0);
		prog_cycle_task(16'b1000001110000110, 1'b0);
		prog_cycle_task(16'b0100001110000110, 1'b1);
		prog_cycle_task(16'b1100001110000110, 1'b0);
		prog_cycle_task(16'b0010001110000110, 1'b0);
		prog_cycle_task(16'b1010001110000110, 1'b0);
		prog_cycle_task(16'b0110001110000110, 1'b0);
		prog_cycle_task(16'b1110001110000110, 1'b1);
		prog_cycle_task(16'b0000011110000110, 1'b0);
		prog_cycle_task(16'b1000011110000110, 1'b0);
		prog_cycle_task(16'b0100011110000110, 1'b1);
		prog_cycle_task(16'b1100011110000110, 1'b0);
		prog_cycle_task(16'b0010011110000110, 1'b0);
		prog_cycle_task(16'b1010011110000110, 1'b0);
		prog_cycle_task(16'b0110011110000110, 1'b0);
		prog_cycle_task(16'b1110011110000110, 1'b1);
		prog_cycle_task(16'b0000000001000110, 1'b0);
		prog_cycle_task(16'b1000000001000110, 1'b0);
		prog_cycle_task(16'b0100000001000110, 1'b1);
		prog_cycle_task(16'b1100000001000110, 1'b0);
		prog_cycle_task(16'b0010000001000110, 1'b0);
		prog_cycle_task(16'b1010000001000110, 1'b1);
		prog_cycle_task(16'b0110000001000110, 1'b0);
		prog_cycle_task(16'b1110000001000110, 1'b0);
		prog_cycle_task(16'b0000010001000110, 1'b0);
		prog_cycle_task(16'b1000010001000110, 1'b0);
		prog_cycle_task(16'b0100010001000110, 1'b1);
		prog_cycle_task(16'b1100010001000110, 1'b0);
		prog_cycle_task(16'b0010010001000110, 1'b0);
		prog_cycle_task(16'b1010010001000110, 1'b0);
		prog_cycle_task(16'b0110010001000110, 1'b0);
		prog_cycle_task(16'b1110010001000110, 1'b1);
		prog_cycle_task(16'b0000001001000110, 1'b0);
		prog_cycle_task(16'b1000001001000110, 1'b0);
		prog_cycle_task(16'b0100001001000110, 1'b1);
		prog_cycle_task(16'b1100001001000110, 1'b0);
		prog_cycle_task(16'b0010001001000110, 1'b0);
		prog_cycle_task(16'b1010001001000110, 1'b0);
		prog_cycle_task(16'b0110001001000110, 1'b0);
		prog_cycle_task(16'b1110001001000110, 1'b1);
		prog_cycle_task(16'b0000011001000110, 1'b1);
		prog_cycle_task(16'b1000011001000110, 1'b0);
		prog_cycle_task(16'b0100011001000110, 1'b0);
		prog_cycle_task(16'b1100011001000110, 1'b0);
		prog_cycle_task(16'b0010011001000110, 1'b1);
		prog_cycle_task(16'b1010011001000110, 1'b0);
		prog_cycle_task(16'b0110011001000110, 1'b0);
		prog_cycle_task(16'b1110011001000110, 1'b0);
		prog_cycle_task(16'b0000000000100110, 1'b1);
		prog_cycle_task(16'b1000000000100110, 1'b0);
		prog_cycle_task(16'b0100000000100110, 1'b0);
		prog_cycle_task(16'b1100000000100110, 1'b1);
		prog_cycle_task(16'b0010000000100110, 1'b0);
		prog_cycle_task(16'b1010000000100110, 1'b0);
		prog_cycle_task(16'b0001000000100110, 1'b1);
		prog_cycle_task(16'b1001000000100110, 1'b0);
		prog_cycle_task(16'b0101000000100110, 1'b0);
		prog_cycle_task(16'b1101000000100110, 1'b1);
		prog_cycle_task(16'b0011000000100110, 1'b0);
		prog_cycle_task(16'b1011000000100110, 1'b0);
		prog_cycle_task(16'b0000100000100110, 1'b1);
		prog_cycle_task(16'b1000100000100110, 1'b0);
		prog_cycle_task(16'b0100100000100110, 1'b0);
		prog_cycle_task(16'b1100100000100110, 1'b1);
		prog_cycle_task(16'b0010100000100110, 1'b0);
		prog_cycle_task(16'b1010100000100110, 1'b0);
		prog_cycle_task(16'b0001100000100110, 1'b1);
		prog_cycle_task(16'b1001100000100110, 1'b0);
		prog_cycle_task(16'b0101100000100110, 1'b0);
		prog_cycle_task(16'b1101100000100110, 1'b1);
		prog_cycle_task(16'b0011100000100110, 1'b0);
		prog_cycle_task(16'b1011100000100110, 1'b0);
		prog_cycle_task(16'b0000010000100110, 1'b1);
		prog_cycle_task(16'b1000010000100110, 1'b0);
		prog_cycle_task(16'b0100010000100110, 1'b0);
		prog_cycle_task(16'b1100010000100110, 1'b1);
		prog_cycle_task(16'b0010010000100110, 1'b0);
		prog_cycle_task(16'b1010010000100110, 1'b0);
		prog_cycle_task(16'b0001010000100110, 1'b1);
		prog_cycle_task(16'b1001010000100110, 1'b0);
		prog_cycle_task(16'b0101010000100110, 1'b0);
		prog_cycle_task(16'b1101010000100110, 1'b1);
		prog_cycle_task(16'b0011010000100110, 1'b0);
		prog_cycle_task(16'b1011010000100110, 1'b0);
		prog_cycle_task(16'b0000110000100110, 1'b1);
		prog_cycle_task(16'b1000110000100110, 1'b1);
		prog_cycle_task(16'b0001110000100110, 1'b1);
		prog_cycle_task(16'b1001110000100110, 1'b1);
		prog_cycle_task(16'b0000001000100110, 1'b1);
		prog_cycle_task(16'b1000001000100110, 1'b1);
		prog_cycle_task(16'b0001001000100110, 1'b1);
		prog_cycle_task(16'b1001001000100110, 1'b1);
		prog_cycle_task(16'b0000101000100110, 1'b1);
		prog_cycle_task(16'b1000101000100110, 1'b1);
		prog_cycle_task(16'b0001101000100110, 1'b1);
		prog_cycle_task(16'b1001101000100110, 1'b1);
		prog_cycle_task(16'b0000011000100110, 1'b1);
		prog_cycle_task(16'b1000011000100110, 1'b1);
		prog_cycle_task(16'b0001011000100110, 1'b1);
		prog_cycle_task(16'b1001011000100110, 1'b1);
		prog_cycle_task(16'b0000111000100110, 1'b1);
		prog_cycle_task(16'b1000111000100110, 1'b1);
		prog_cycle_task(16'b0000000000010110, 1'b1);
		prog_cycle_task(16'b1000000000010110, 1'b0);
		prog_cycle_task(16'b0100000000010110, 1'b0);
		prog_cycle_task(16'b1100000000010110, 1'b1);
		prog_cycle_task(16'b0010000000010110, 1'b0);
		prog_cycle_task(16'b1010000000010110, 1'b0);
		prog_cycle_task(16'b0001000000010110, 1'b1);
		prog_cycle_task(16'b1001000000010110, 1'b1);
		prog_cycle_task(16'b0000100000010110, 1'b1);
		prog_cycle_task(16'b1000100000010110, 1'b0);
		prog_cycle_task(16'b0100100000010110, 1'b0);
		prog_cycle_task(16'b1100100000010110, 1'b1);
		prog_cycle_task(16'b0010100000010110, 1'b0);
		prog_cycle_task(16'b1010100000010110, 1'b0);
		prog_cycle_task(16'b0001100000010110, 1'b1);
		prog_cycle_task(16'b1001100000010110, 1'b0);
		prog_cycle_task(16'b0101100000010110, 1'b0);
		prog_cycle_task(16'b1101100000010110, 1'b0);
		prog_cycle_task(16'b0011100000010110, 1'b1);
		prog_cycle_task(16'b1011100000010110, 1'b0);
		prog_cycle_task(16'b0000010000010110, 1'b1);
		prog_cycle_task(16'b1000010000010110, 1'b1);
		prog_cycle_task(16'b0001010000010110, 1'b1);
		prog_cycle_task(16'b1001010000010110, 1'b1);
		prog_cycle_task(16'b0000000000110110, 1'b1);
		prog_cycle_task(16'b1000000000110110, 1'b0);
		prog_cycle_task(16'b0100000000110110, 1'b0);
		prog_cycle_task(16'b1100000000110110, 1'b1);
		prog_cycle_task(16'b0010000000110110, 1'b0);
		prog_cycle_task(16'b1010000000110110, 1'b0);
		prog_cycle_task(16'b0001000000110110, 1'b1);
		prog_cycle_task(16'b1001000000110110, 1'b0);
		prog_cycle_task(16'b0101000000110110, 1'b0);
		prog_cycle_task(16'b1101000000110110, 1'b1);
		prog_cycle_task(16'b0011000000110110, 1'b0);
		prog_cycle_task(16'b1011000000110110, 1'b0);
		prog_cycle_task(16'b0000100000110110, 1'b0);
		prog_cycle_task(16'b1000100000110110, 1'b1);
		prog_cycle_task(16'b0100100000110110, 1'b0);
		prog_cycle_task(16'b1100100000110110, 1'b1);
		prog_cycle_task(16'b0010100000110110, 1'b0);
		prog_cycle_task(16'b1010100000110110, 1'b0);
		prog_cycle_task(16'b0001100000110110, 1'b1);
		prog_cycle_task(16'b1001100000110110, 1'b0);
		prog_cycle_task(16'b0101100000110110, 1'b0);
		prog_cycle_task(16'b1101100000110110, 1'b1);
		prog_cycle_task(16'b0011100000110110, 1'b0);
		prog_cycle_task(16'b1011100000110110, 1'b0);
		prog_cycle_task(16'b0000010000110110, 1'b0);
		prog_cycle_task(16'b1000010000110110, 1'b1);
		prog_cycle_task(16'b0100010000110110, 1'b0);
		prog_cycle_task(16'b1100010000110110, 1'b1);
		prog_cycle_task(16'b0010010000110110, 1'b0);
		prog_cycle_task(16'b1010010000110110, 1'b0);
		prog_cycle_task(16'b0001010000110110, 1'b1);
		prog_cycle_task(16'b1001010000110110, 1'b0);
		prog_cycle_task(16'b0101010000110110, 1'b0);
		prog_cycle_task(16'b1101010000110110, 1'b1);
		prog_cycle_task(16'b0011010000110110, 1'b0);
		prog_cycle_task(16'b1011010000110110, 1'b0);
		prog_cycle_task(16'b0000110000110110, 1'b0);
		prog_cycle_task(16'b1000110000110110, 1'b1);
		prog_cycle_task(16'b0100110000110110, 1'b0);
		prog_cycle_task(16'b1100110000110110, 1'b1);
		prog_cycle_task(16'b0010110000110110, 1'b0);
		prog_cycle_task(16'b1010110000110110, 1'b0);
		prog_cycle_task(16'b0001110000110110, 1'b1);
		prog_cycle_task(16'b1001110000110110, 1'b0);
		prog_cycle_task(16'b0101110000110110, 1'b0);
		prog_cycle_task(16'b1101110000110110, 1'b1);
		prog_cycle_task(16'b0011110000110110, 1'b0);
		prog_cycle_task(16'b1011110000110110, 1'b0);
		prog_cycle_task(16'b0000001000110110, 1'b0);
		prog_cycle_task(16'b1000001000110110, 1'b1);
		prog_cycle_task(16'b0100001000110110, 1'b0);
		prog_cycle_task(16'b1100001000110110, 1'b1);
		prog_cycle_task(16'b0010001000110110, 1'b0);
		prog_cycle_task(16'b1010001000110110, 1'b0);
		prog_cycle_task(16'b0001001000110110, 1'b1);
		prog_cycle_task(16'b1001001000110110, 1'b1);
		prog_cycle_task(16'b0000101000110110, 1'b0);
		prog_cycle_task(16'b1000101000110110, 1'b1);
		prog_cycle_task(16'b0000000000001110, 1'b0);
		prog_cycle_task(16'b1000000000001110, 1'b0);
		prog_cycle_task(16'b0100000000001110, 1'b0);
		prog_cycle_task(16'b1100000000001110, 1'b0);
		prog_cycle_task(16'b0010000000001110, 1'b0);
		prog_cycle_task(16'b1010000000001110, 1'b0);
		prog_cycle_task(16'b0110000000001110, 1'b0);
		prog_cycle_task(16'b1110000000001110, 1'b0);
		prog_cycle_task(16'b0001000000001110, 1'b0);
		prog_cycle_task(16'b1001000000001110, 1'b0);
		prog_cycle_task(16'b0101000000001110, 1'b0);
		prog_cycle_task(16'b1101000000001110, 1'b0);
		prog_cycle_task(16'b0011000000001110, 1'b0);
		prog_cycle_task(16'b1011000000001110, 1'b0);
		prog_cycle_task(16'b0111000000001110, 1'b0);
		prog_cycle_task(16'b1111000000001110, 1'b0);
		prog_cycle_task(16'b0000100000001110, 1'b0);
		prog_cycle_task(16'b1000100000001110, 1'b0);
		prog_cycle_task(16'b0100100000001110, 1'b1);
		prog_cycle_task(16'b0000010000001110, 1'b0);
		prog_cycle_task(16'b1000010000001110, 1'b0);
		prog_cycle_task(16'b0100010000001110, 1'b0);
		prog_cycle_task(16'b1100010000001110, 1'b0);
		prog_cycle_task(16'b0010010000001110, 1'b0);
		prog_cycle_task(16'b1010010000001110, 1'b0);
		prog_cycle_task(16'b0110010000001110, 1'b0);
		prog_cycle_task(16'b1110010000001110, 1'b0);
		prog_cycle_task(16'b0001010000001110, 1'b0);
		prog_cycle_task(16'b1001010000001110, 1'b0);
		prog_cycle_task(16'b0101010000001110, 1'b0);
		prog_cycle_task(16'b1101010000001110, 1'b0);
		prog_cycle_task(16'b0011010000001110, 1'b0);
		prog_cycle_task(16'b1011010000001110, 1'b0);
		prog_cycle_task(16'b0111010000001110, 1'b0);
		prog_cycle_task(16'b1111010000001110, 1'b0);
		prog_cycle_task(16'b0000110000001110, 1'b0);
		prog_cycle_task(16'b1000110000001110, 1'b0);
		prog_cycle_task(16'b0100110000001110, 1'b1);
		prog_cycle_task(16'b0000001000001110, 1'b0);
		prog_cycle_task(16'b1000001000001110, 1'b0);
		prog_cycle_task(16'b0100001000001110, 1'b0);
		prog_cycle_task(16'b1100001000001110, 1'b0);
		prog_cycle_task(16'b0010001000001110, 1'b0);
		prog_cycle_task(16'b1010001000001110, 1'b0);
		prog_cycle_task(16'b0110001000001110, 1'b0);
		prog_cycle_task(16'b1110001000001110, 1'b0);
		prog_cycle_task(16'b0001001000001110, 1'b0);
		prog_cycle_task(16'b1001001000001110, 1'b0);
		prog_cycle_task(16'b0101001000001110, 1'b0);
		prog_cycle_task(16'b1101001000001110, 1'b0);
		prog_cycle_task(16'b0011001000001110, 1'b0);
		prog_cycle_task(16'b1011001000001110, 1'b0);
		prog_cycle_task(16'b0111001000001110, 1'b0);
		prog_cycle_task(16'b1111001000001110, 1'b0);
		prog_cycle_task(16'b0000101000001110, 1'b0);
		prog_cycle_task(16'b1000101000001110, 1'b0);
		prog_cycle_task(16'b0100101000001110, 1'b1);
		prog_cycle_task(16'b0000011000001110, 1'b0);
		prog_cycle_task(16'b1000011000001110, 1'b0);
		prog_cycle_task(16'b0100011000001110, 1'b0);
		prog_cycle_task(16'b1100011000001110, 1'b0);
		prog_cycle_task(16'b0010011000001110, 1'b0);
		prog_cycle_task(16'b1010011000001110, 1'b0);
		prog_cycle_task(16'b0110011000001110, 1'b0);
		prog_cycle_task(16'b1110011000001110, 1'b0);
		prog_cycle_task(16'b0001011000001110, 1'b0);
		prog_cycle_task(16'b1001011000001110, 1'b0);
		prog_cycle_task(16'b0101011000001110, 1'b0);
		prog_cycle_task(16'b1101011000001110, 1'b0);
		prog_cycle_task(16'b0011011000001110, 1'b0);
		prog_cycle_task(16'b1011011000001110, 1'b0);
		prog_cycle_task(16'b0111011000001110, 1'b0);
		prog_cycle_task(16'b1111011000001110, 1'b0);
		prog_cycle_task(16'b0000111000001110, 1'b0);
		prog_cycle_task(16'b1000111000001110, 1'b0);
		prog_cycle_task(16'b0100111000001110, 1'b1);
		prog_cycle_task(16'b0000000100001110, 1'b0);
		prog_cycle_task(16'b1000000100001110, 1'b0);
		prog_cycle_task(16'b0100000100001110, 1'b1);
		prog_cycle_task(16'b1100000100001110, 1'b0);
		prog_cycle_task(16'b0010000100001110, 1'b0);
		prog_cycle_task(16'b1010000100001110, 1'b0);
		prog_cycle_task(16'b0110000100001110, 1'b0);
		prog_cycle_task(16'b1110000100001110, 1'b1);
		prog_cycle_task(16'b0000010100001110, 1'b0);
		prog_cycle_task(16'b1000010100001110, 1'b0);
		prog_cycle_task(16'b0100010100001110, 1'b1);
		prog_cycle_task(16'b1100010100001110, 1'b0);
		prog_cycle_task(16'b0010010100001110, 1'b0);
		prog_cycle_task(16'b1010010100001110, 1'b0);
		prog_cycle_task(16'b0110010100001110, 1'b0);
		prog_cycle_task(16'b1110010100001110, 1'b1);
		prog_cycle_task(16'b0000001100001110, 1'b0);
		prog_cycle_task(16'b1000001100001110, 1'b0);
		prog_cycle_task(16'b0100001100001110, 1'b1);
		prog_cycle_task(16'b1100001100001110, 1'b0);
		prog_cycle_task(16'b0010001100001110, 1'b0);
		prog_cycle_task(16'b1010001100001110, 1'b0);
		prog_cycle_task(16'b0110001100001110, 1'b0);
		prog_cycle_task(16'b1110001100001110, 1'b1);
		prog_cycle_task(16'b0000011100001110, 1'b0);
		prog_cycle_task(16'b1000011100001110, 1'b0);
		prog_cycle_task(16'b0100011100001110, 1'b1);
		prog_cycle_task(16'b1100011100001110, 1'b0);
		prog_cycle_task(16'b0010011100001110, 1'b0);
		prog_cycle_task(16'b1010011100001110, 1'b0);
		prog_cycle_task(16'b0110011100001110, 1'b0);
		prog_cycle_task(16'b1110011100001110, 1'b1);
		prog_cycle_task(16'b0000000010001110, 1'b0);
		prog_cycle_task(16'b1000000010001110, 1'b0);
		prog_cycle_task(16'b0100000010001110, 1'b1);
		prog_cycle_task(16'b1100000010001110, 1'b0);
		prog_cycle_task(16'b0010000010001110, 1'b0);
		prog_cycle_task(16'b1010000010001110, 1'b0);
		prog_cycle_task(16'b0110000010001110, 1'b0);
		prog_cycle_task(16'b1110000010001110, 1'b1);
		prog_cycle_task(16'b0000010010001110, 1'b0);
		prog_cycle_task(16'b1000010010001110, 1'b0);
		prog_cycle_task(16'b0100010010001110, 1'b1);
		prog_cycle_task(16'b1100010010001110, 1'b0);
		prog_cycle_task(16'b0010010010001110, 1'b0);
		prog_cycle_task(16'b1010010010001110, 1'b0);
		prog_cycle_task(16'b0110010010001110, 1'b0);
		prog_cycle_task(16'b1110010010001110, 1'b1);
		prog_cycle_task(16'b0000001010001110, 1'b0);
		prog_cycle_task(16'b1000001010001110, 1'b0);
		prog_cycle_task(16'b0100001010001110, 1'b1);
		prog_cycle_task(16'b1100001010001110, 1'b0);
		prog_cycle_task(16'b0010001010001110, 1'b0);
		prog_cycle_task(16'b1010001010001110, 1'b0);
		prog_cycle_task(16'b0110001010001110, 1'b0);
		prog_cycle_task(16'b1110001010001110, 1'b1);
		prog_cycle_task(16'b0000011010001110, 1'b0);
		prog_cycle_task(16'b1000011010001110, 1'b0);
		prog_cycle_task(16'b0100011010001110, 1'b1);
		prog_cycle_task(16'b1100011010001110, 1'b0);
		prog_cycle_task(16'b0010011010001110, 1'b0);
		prog_cycle_task(16'b1010011010001110, 1'b0);
		prog_cycle_task(16'b0110011010001110, 1'b0);
		prog_cycle_task(16'b1110011010001110, 1'b1);
		prog_cycle_task(16'b0000000110001110, 1'b0);
		prog_cycle_task(16'b1000000110001110, 1'b0);
		prog_cycle_task(16'b0100000110001110, 1'b1);
		prog_cycle_task(16'b1100000110001110, 1'b0);
		prog_cycle_task(16'b0010000110001110, 1'b0);
		prog_cycle_task(16'b1010000110001110, 1'b0);
		prog_cycle_task(16'b0110000110001110, 1'b0);
		prog_cycle_task(16'b1110000110001110, 1'b1);
		prog_cycle_task(16'b0000010110001110, 1'b0);
		prog_cycle_task(16'b1000010110001110, 1'b0);
		prog_cycle_task(16'b0100010110001110, 1'b1);
		prog_cycle_task(16'b1100010110001110, 1'b0);
		prog_cycle_task(16'b0010010110001110, 1'b0);
		prog_cycle_task(16'b1010010110001110, 1'b0);
		prog_cycle_task(16'b0110010110001110, 1'b0);
		prog_cycle_task(16'b1110010110001110, 1'b1);
		prog_cycle_task(16'b0000001110001110, 1'b0);
		prog_cycle_task(16'b1000001110001110, 1'b0);
		prog_cycle_task(16'b0100001110001110, 1'b1);
		prog_cycle_task(16'b1100001110001110, 1'b0);
		prog_cycle_task(16'b0010001110001110, 1'b0);
		prog_cycle_task(16'b1010001110001110, 1'b0);
		prog_cycle_task(16'b0110001110001110, 1'b0);
		prog_cycle_task(16'b1110001110001110, 1'b1);
		prog_cycle_task(16'b0000011110001110, 1'b0);
		prog_cycle_task(16'b1000011110001110, 1'b0);
		prog_cycle_task(16'b0100011110001110, 1'b1);
		prog_cycle_task(16'b1100011110001110, 1'b0);
		prog_cycle_task(16'b0010011110001110, 1'b0);
		prog_cycle_task(16'b1010011110001110, 1'b0);
		prog_cycle_task(16'b0110011110001110, 1'b0);
		prog_cycle_task(16'b1110011110001110, 1'b1);
		prog_cycle_task(16'b0000000001001110, 1'b0);
		prog_cycle_task(16'b1000000001001110, 1'b0);
		prog_cycle_task(16'b0100000001001110, 1'b1);
		prog_cycle_task(16'b1100000001001110, 1'b0);
		prog_cycle_task(16'b0010000001001110, 1'b0);
		prog_cycle_task(16'b1010000001001110, 1'b0);
		prog_cycle_task(16'b0110000001001110, 1'b0);
		prog_cycle_task(16'b1110000001001110, 1'b1);
		prog_cycle_task(16'b0000010001001110, 1'b0);
		prog_cycle_task(16'b1000010001001110, 1'b0);
		prog_cycle_task(16'b0100010001001110, 1'b1);
		prog_cycle_task(16'b1100010001001110, 1'b0);
		prog_cycle_task(16'b0010010001001110, 1'b0);
		prog_cycle_task(16'b1010010001001110, 1'b0);
		prog_cycle_task(16'b0110010001001110, 1'b0);
		prog_cycle_task(16'b1110010001001110, 1'b1);
		prog_cycle_task(16'b0000001001001110, 1'b0);
		prog_cycle_task(16'b1000001001001110, 1'b0);
		prog_cycle_task(16'b0100001001001110, 1'b1);
		prog_cycle_task(16'b1100001001001110, 1'b0);
		prog_cycle_task(16'b0010001001001110, 1'b0);
		prog_cycle_task(16'b1010001001001110, 1'b0);
		prog_cycle_task(16'b0110001001001110, 1'b0);
		prog_cycle_task(16'b1110001001001110, 1'b1);
		prog_cycle_task(16'b0000011001001110, 1'b0);
		prog_cycle_task(16'b1000011001001110, 1'b0);
		prog_cycle_task(16'b0100011001001110, 1'b1);
		prog_cycle_task(16'b1100011001001110, 1'b0);
		prog_cycle_task(16'b0010011001001110, 1'b0);
		prog_cycle_task(16'b1010011001001110, 1'b0);
		prog_cycle_task(16'b0110011001001110, 1'b0);
		prog_cycle_task(16'b1110011001001110, 1'b1);
		prog_cycle_task(16'b0000000000101110, 1'b1);
		prog_cycle_task(16'b1000000000101110, 1'b0);
		prog_cycle_task(16'b0100000000101110, 1'b0);
		prog_cycle_task(16'b1100000000101110, 1'b0);
		prog_cycle_task(16'b0010000000101110, 1'b1);
		prog_cycle_task(16'b1010000000101110, 1'b0);
		prog_cycle_task(16'b0110000000101110, 1'b0);
		prog_cycle_task(16'b1110000000101110, 1'b0);
		prog_cycle_task(16'b0001000000101110, 1'b1);
		prog_cycle_task(16'b1001000000101110, 1'b0);
		prog_cycle_task(16'b0101000000101110, 1'b0);
		prog_cycle_task(16'b1101000000101110, 1'b0);
		prog_cycle_task(16'b0011000000101110, 1'b1);
		prog_cycle_task(16'b1011000000101110, 1'b0);
		prog_cycle_task(16'b0111000000101110, 1'b0);
		prog_cycle_task(16'b1111000000101110, 1'b0);
		prog_cycle_task(16'b0000100000101110, 1'b1);
		prog_cycle_task(16'b1000100000101110, 1'b0);
		prog_cycle_task(16'b0100100000101110, 1'b0);
		prog_cycle_task(16'b1100100000101110, 1'b1);
		prog_cycle_task(16'b0010100000101110, 1'b0);
		prog_cycle_task(16'b1010100000101110, 1'b0);
		prog_cycle_task(16'b0001100000101110, 1'b1);
		prog_cycle_task(16'b1001100000101110, 1'b0);
		prog_cycle_task(16'b0101100000101110, 1'b0);
		prog_cycle_task(16'b1101100000101110, 1'b0);
		prog_cycle_task(16'b0011100000101110, 1'b1);
		prog_cycle_task(16'b1011100000101110, 1'b0);
		prog_cycle_task(16'b0111100000101110, 1'b0);
		prog_cycle_task(16'b1111100000101110, 1'b0);
		prog_cycle_task(16'b0000010000101110, 1'b1);
		prog_cycle_task(16'b1000010000101110, 1'b0);
		prog_cycle_task(16'b0100010000101110, 1'b0);
		prog_cycle_task(16'b1100010000101110, 1'b0);
		prog_cycle_task(16'b0010010000101110, 1'b1);
		prog_cycle_task(16'b1010010000101110, 1'b0);
		prog_cycle_task(16'b0110010000101110, 1'b0);
		prog_cycle_task(16'b1110010000101110, 1'b0);
		prog_cycle_task(16'b0001010000101110, 1'b1);
		prog_cycle_task(16'b1001010000101110, 1'b0);
		prog_cycle_task(16'b0101010000101110, 1'b0);
		prog_cycle_task(16'b1101010000101110, 1'b1);
		prog_cycle_task(16'b0011010000101110, 1'b0);
		prog_cycle_task(16'b1011010000101110, 1'b0);
		prog_cycle_task(16'b0000110000101110, 1'b0);
		prog_cycle_task(16'b1000110000101110, 1'b0);
		prog_cycle_task(16'b0100110000101110, 1'b1);
		prog_cycle_task(16'b1100110000101110, 1'b0);
		prog_cycle_task(16'b0010110000101110, 1'b1);
		prog_cycle_task(16'b1010110000101110, 1'b0);
		prog_cycle_task(16'b0110110000101110, 1'b0);
		prog_cycle_task(16'b1110110000101110, 1'b0);
		prog_cycle_task(16'b0001110000101110, 1'b1);
		prog_cycle_task(16'b1001110000101110, 1'b0);
		prog_cycle_task(16'b0101110000101110, 1'b0);
		prog_cycle_task(16'b1101110000101110, 1'b0);
		prog_cycle_task(16'b0011110000101110, 1'b1);
		prog_cycle_task(16'b1011110000101110, 1'b0);
		prog_cycle_task(16'b0111110000101110, 1'b0);
		prog_cycle_task(16'b1111110000101110, 1'b0);
		prog_cycle_task(16'b0000001000101110, 1'b1);
		prog_cycle_task(16'b1000001000101110, 1'b0);
		prog_cycle_task(16'b0100001000101110, 1'b0);
		prog_cycle_task(16'b1100001000101110, 1'b1);
		prog_cycle_task(16'b0010001000101110, 1'b0);
		prog_cycle_task(16'b1010001000101110, 1'b0);
		prog_cycle_task(16'b0001001000101110, 1'b1);
		prog_cycle_task(16'b1001001000101110, 1'b0);
		prog_cycle_task(16'b0101001000101110, 1'b0);
		prog_cycle_task(16'b1101001000101110, 1'b0);
		prog_cycle_task(16'b0011001000101110, 1'b1);
		prog_cycle_task(16'b1011001000101110, 1'b0);
		prog_cycle_task(16'b0111001000101110, 1'b0);
		prog_cycle_task(16'b1111001000101110, 1'b0);
		prog_cycle_task(16'b0000101000101110, 1'b1);
		prog_cycle_task(16'b1000101000101110, 1'b0);
		prog_cycle_task(16'b0100101000101110, 1'b0);
		prog_cycle_task(16'b1100101000101110, 1'b0);
		prog_cycle_task(16'b0010101000101110, 1'b1);
		prog_cycle_task(16'b1010101000101110, 1'b0);
		prog_cycle_task(16'b0110101000101110, 1'b0);
		prog_cycle_task(16'b1110101000101110, 1'b0);
		prog_cycle_task(16'b0001101000101110, 1'b1);
		prog_cycle_task(16'b1001101000101110, 1'b0);
		prog_cycle_task(16'b0101101000101110, 1'b0);
		prog_cycle_task(16'b1101101000101110, 1'b1);
		prog_cycle_task(16'b0011101000101110, 1'b0);
		prog_cycle_task(16'b1011101000101110, 1'b0);
		prog_cycle_task(16'b0000000000011110, 1'b1);
		prog_cycle_task(16'b1000000000011110, 1'b0);
		prog_cycle_task(16'b0100000000011110, 1'b0);
		prog_cycle_task(16'b1100000000011110, 1'b1);
		prog_cycle_task(16'b0010000000011110, 1'b0);
		prog_cycle_task(16'b1010000000011110, 1'b0);
		prog_cycle_task(16'b0001000000011110, 1'b1);
		prog_cycle_task(16'b1001000000011110, 1'b1);
		prog_cycle_task(16'b0000100000011110, 1'b1);
		prog_cycle_task(16'b1000100000011110, 1'b0);
		prog_cycle_task(16'b0100100000011110, 1'b0);
		prog_cycle_task(16'b1100100000011110, 1'b1);
		prog_cycle_task(16'b0010100000011110, 1'b0);
		prog_cycle_task(16'b1010100000011110, 1'b0);
		prog_cycle_task(16'b0001100000011110, 1'b1);
		prog_cycle_task(16'b1001100000011110, 1'b0);
		prog_cycle_task(16'b0101100000011110, 1'b0);
		prog_cycle_task(16'b1101100000011110, 1'b1);
		prog_cycle_task(16'b0011100000011110, 1'b0);
		prog_cycle_task(16'b1011100000011110, 1'b0);
		prog_cycle_task(16'b0000010000011110, 1'b1);
		prog_cycle_task(16'b1000010000011110, 1'b1);
		prog_cycle_task(16'b0001010000011110, 1'b1);
		prog_cycle_task(16'b1001010000011110, 1'b1);
		prog_cycle_task(16'b0000000000111110, 1'b1);
		prog_cycle_task(16'b1000000000111110, 1'b0);
		prog_cycle_task(16'b0100000000111110, 1'b0);
		prog_cycle_task(16'b1100000000111110, 1'b1);
		prog_cycle_task(16'b0010000000111110, 1'b0);
		prog_cycle_task(16'b1010000000111110, 1'b0);
		prog_cycle_task(16'b0001000000111110, 1'b1);
		prog_cycle_task(16'b1001000000111110, 1'b1);
		prog_cycle_task(16'b0000100000111110, 1'b1);
		prog_cycle_task(16'b1000100000111110, 1'b0);
		prog_cycle_task(16'b0100100000111110, 1'b0);
		prog_cycle_task(16'b1100100000111110, 1'b1);
		prog_cycle_task(16'b0010100000111110, 1'b0);
		prog_cycle_task(16'b1010100000111110, 1'b0);
		prog_cycle_task(16'b0001100000111110, 1'b1);
		prog_cycle_task(16'b1001100000111110, 1'b1);
		prog_cycle_task(16'b0000010000111110, 1'b1);
		prog_cycle_task(16'b1000010000111110, 1'b1);
		prog_cycle_task(16'b0000000000000001, 1'b0);
		prog_cycle_task(16'b1000000000000001, 1'b0);
		prog_cycle_task(16'b0100000000000001, 1'b0);
		prog_cycle_task(16'b1100000000000001, 1'b0);
		prog_cycle_task(16'b0010000000000001, 1'b0);
		prog_cycle_task(16'b1010000000000001, 1'b0);
		prog_cycle_task(16'b0110000000000001, 1'b0);
		prog_cycle_task(16'b1110000000000001, 1'b0);
		prog_cycle_task(16'b0001000000000001, 1'b0);
		prog_cycle_task(16'b1001000000000001, 1'b0);
		prog_cycle_task(16'b0101000000000001, 1'b0);
		prog_cycle_task(16'b1101000000000001, 1'b0);
		prog_cycle_task(16'b0011000000000001, 1'b0);
		prog_cycle_task(16'b1011000000000001, 1'b0);
		prog_cycle_task(16'b0111000000000001, 1'b0);
		prog_cycle_task(16'b1111000000000001, 1'b0);
		prog_cycle_task(16'b0000100000000001, 1'b0);
		prog_cycle_task(16'b1000100000000001, 1'b0);
		prog_cycle_task(16'b0100100000000001, 1'b1);
		prog_cycle_task(16'b0000010000000001, 1'b0);
		prog_cycle_task(16'b1000010000000001, 1'b0);
		prog_cycle_task(16'b0100010000000001, 1'b0);
		prog_cycle_task(16'b1100010000000001, 1'b0);
		prog_cycle_task(16'b0010010000000001, 1'b0);
		prog_cycle_task(16'b1010010000000001, 1'b0);
		prog_cycle_task(16'b0110010000000001, 1'b0);
		prog_cycle_task(16'b1110010000000001, 1'b0);
		prog_cycle_task(16'b0001010000000001, 1'b0);
		prog_cycle_task(16'b1001010000000001, 1'b0);
		prog_cycle_task(16'b0101010000000001, 1'b0);
		prog_cycle_task(16'b1101010000000001, 1'b0);
		prog_cycle_task(16'b0011010000000001, 1'b0);
		prog_cycle_task(16'b1011010000000001, 1'b0);
		prog_cycle_task(16'b0111010000000001, 1'b0);
		prog_cycle_task(16'b1111010000000001, 1'b0);
		prog_cycle_task(16'b0000110000000001, 1'b0);
		prog_cycle_task(16'b1000110000000001, 1'b0);
		prog_cycle_task(16'b0100110000000001, 1'b1);
		prog_cycle_task(16'b0000001000000001, 1'b0);
		prog_cycle_task(16'b1000001000000001, 1'b0);
		prog_cycle_task(16'b0100001000000001, 1'b0);
		prog_cycle_task(16'b1100001000000001, 1'b0);
		prog_cycle_task(16'b0010001000000001, 1'b0);
		prog_cycle_task(16'b1010001000000001, 1'b0);
		prog_cycle_task(16'b0110001000000001, 1'b0);
		prog_cycle_task(16'b1110001000000001, 1'b0);
		prog_cycle_task(16'b0001001000000001, 1'b0);
		prog_cycle_task(16'b1001001000000001, 1'b0);
		prog_cycle_task(16'b0101001000000001, 1'b0);
		prog_cycle_task(16'b1101001000000001, 1'b0);
		prog_cycle_task(16'b0011001000000001, 1'b0);
		prog_cycle_task(16'b1011001000000001, 1'b0);
		prog_cycle_task(16'b0111001000000001, 1'b0);
		prog_cycle_task(16'b1111001000000001, 1'b0);
		prog_cycle_task(16'b0000101000000001, 1'b0);
		prog_cycle_task(16'b1000101000000001, 1'b0);
		prog_cycle_task(16'b0100101000000001, 1'b1);
		prog_cycle_task(16'b0000011000000001, 1'b0);
		prog_cycle_task(16'b1000011000000001, 1'b0);
		prog_cycle_task(16'b0100011000000001, 1'b0);
		prog_cycle_task(16'b1100011000000001, 1'b0);
		prog_cycle_task(16'b0010011000000001, 1'b0);
		prog_cycle_task(16'b1010011000000001, 1'b0);
		prog_cycle_task(16'b0110011000000001, 1'b0);
		prog_cycle_task(16'b1110011000000001, 1'b0);
		prog_cycle_task(16'b0001011000000001, 1'b0);
		prog_cycle_task(16'b1001011000000001, 1'b0);
		prog_cycle_task(16'b0101011000000001, 1'b0);
		prog_cycle_task(16'b1101011000000001, 1'b0);
		prog_cycle_task(16'b0011011000000001, 1'b0);
		prog_cycle_task(16'b1011011000000001, 1'b0);
		prog_cycle_task(16'b0111011000000001, 1'b0);
		prog_cycle_task(16'b1111011000000001, 1'b0);
		prog_cycle_task(16'b0000111000000001, 1'b0);
		prog_cycle_task(16'b1000111000000001, 1'b0);
		prog_cycle_task(16'b0100111000000001, 1'b1);
		prog_cycle_task(16'b0000000100000001, 1'b0);
		prog_cycle_task(16'b1000000100000001, 1'b0);
		prog_cycle_task(16'b0100000100000001, 1'b1);
		prog_cycle_task(16'b1100000100000001, 1'b0);
		prog_cycle_task(16'b0010000100000001, 1'b0);
		prog_cycle_task(16'b1010000100000001, 1'b0);
		prog_cycle_task(16'b0110000100000001, 1'b0);
		prog_cycle_task(16'b1110000100000001, 1'b1);
		prog_cycle_task(16'b0000010100000001, 1'b0);
		prog_cycle_task(16'b1000010100000001, 1'b0);
		prog_cycle_task(16'b0100010100000001, 1'b1);
		prog_cycle_task(16'b1100010100000001, 1'b0);
		prog_cycle_task(16'b0010010100000001, 1'b0);
		prog_cycle_task(16'b1010010100000001, 1'b0);
		prog_cycle_task(16'b0110010100000001, 1'b0);
		prog_cycle_task(16'b1110010100000001, 1'b1);
		prog_cycle_task(16'b0000001100000001, 1'b0);
		prog_cycle_task(16'b1000001100000001, 1'b0);
		prog_cycle_task(16'b0100001100000001, 1'b1);
		prog_cycle_task(16'b1100001100000001, 1'b0);
		prog_cycle_task(16'b0010001100000001, 1'b0);
		prog_cycle_task(16'b1010001100000001, 1'b0);
		prog_cycle_task(16'b0110001100000001, 1'b0);
		prog_cycle_task(16'b1110001100000001, 1'b1);
		prog_cycle_task(16'b0000011100000001, 1'b0);
		prog_cycle_task(16'b1000011100000001, 1'b0);
		prog_cycle_task(16'b0100011100000001, 1'b1);
		prog_cycle_task(16'b1100011100000001, 1'b0);
		prog_cycle_task(16'b0010011100000001, 1'b0);
		prog_cycle_task(16'b1010011100000001, 1'b0);
		prog_cycle_task(16'b0110011100000001, 1'b0);
		prog_cycle_task(16'b1110011100000001, 1'b1);
		prog_cycle_task(16'b0000000010000001, 1'b0);
		prog_cycle_task(16'b1000000010000001, 1'b0);
		prog_cycle_task(16'b0100000010000001, 1'b1);
		prog_cycle_task(16'b1100000010000001, 1'b0);
		prog_cycle_task(16'b0010000010000001, 1'b0);
		prog_cycle_task(16'b1010000010000001, 1'b0);
		prog_cycle_task(16'b0110000010000001, 1'b0);
		prog_cycle_task(16'b1110000010000001, 1'b1);
		prog_cycle_task(16'b0000010010000001, 1'b0);
		prog_cycle_task(16'b1000010010000001, 1'b0);
		prog_cycle_task(16'b0100010010000001, 1'b1);
		prog_cycle_task(16'b1100010010000001, 1'b0);
		prog_cycle_task(16'b0010010010000001, 1'b0);
		prog_cycle_task(16'b1010010010000001, 1'b0);
		prog_cycle_task(16'b0110010010000001, 1'b0);
		prog_cycle_task(16'b1110010010000001, 1'b1);
		prog_cycle_task(16'b0000001010000001, 1'b0);
		prog_cycle_task(16'b1000001010000001, 1'b0);
		prog_cycle_task(16'b0100001010000001, 1'b1);
		prog_cycle_task(16'b1100001010000001, 1'b0);
		prog_cycle_task(16'b0010001010000001, 1'b0);
		prog_cycle_task(16'b1010001010000001, 1'b0);
		prog_cycle_task(16'b0110001010000001, 1'b0);
		prog_cycle_task(16'b1110001010000001, 1'b1);
		prog_cycle_task(16'b0000011010000001, 1'b0);
		prog_cycle_task(16'b1000011010000001, 1'b0);
		prog_cycle_task(16'b0100011010000001, 1'b1);
		prog_cycle_task(16'b1100011010000001, 1'b0);
		prog_cycle_task(16'b0010011010000001, 1'b0);
		prog_cycle_task(16'b1010011010000001, 1'b0);
		prog_cycle_task(16'b0110011010000001, 1'b0);
		prog_cycle_task(16'b1110011010000001, 1'b1);
		prog_cycle_task(16'b0000000110000001, 1'b0);
		prog_cycle_task(16'b1000000110000001, 1'b0);
		prog_cycle_task(16'b0100000110000001, 1'b1);
		prog_cycle_task(16'b1100000110000001, 1'b0);
		prog_cycle_task(16'b0010000110000001, 1'b0);
		prog_cycle_task(16'b1010000110000001, 1'b0);
		prog_cycle_task(16'b0110000110000001, 1'b0);
		prog_cycle_task(16'b1110000110000001, 1'b1);
		prog_cycle_task(16'b0000010110000001, 1'b0);
		prog_cycle_task(16'b1000010110000001, 1'b0);
		prog_cycle_task(16'b0100010110000001, 1'b1);
		prog_cycle_task(16'b1100010110000001, 1'b0);
		prog_cycle_task(16'b0010010110000001, 1'b0);
		prog_cycle_task(16'b1010010110000001, 1'b0);
		prog_cycle_task(16'b0110010110000001, 1'b0);
		prog_cycle_task(16'b1110010110000001, 1'b1);
		prog_cycle_task(16'b0000001110000001, 1'b0);
		prog_cycle_task(16'b1000001110000001, 1'b0);
		prog_cycle_task(16'b0100001110000001, 1'b1);
		prog_cycle_task(16'b1100001110000001, 1'b0);
		prog_cycle_task(16'b0010001110000001, 1'b0);
		prog_cycle_task(16'b1010001110000001, 1'b0);
		prog_cycle_task(16'b0110001110000001, 1'b0);
		prog_cycle_task(16'b1110001110000001, 1'b1);
		prog_cycle_task(16'b0000011110000001, 1'b0);
		prog_cycle_task(16'b1000011110000001, 1'b0);
		prog_cycle_task(16'b0100011110000001, 1'b1);
		prog_cycle_task(16'b1100011110000001, 1'b0);
		prog_cycle_task(16'b0010011110000001, 1'b0);
		prog_cycle_task(16'b1010011110000001, 1'b0);
		prog_cycle_task(16'b0110011110000001, 1'b0);
		prog_cycle_task(16'b1110011110000001, 1'b1);
		prog_cycle_task(16'b0000000001000001, 1'b0);
		prog_cycle_task(16'b1000000001000001, 1'b0);
		prog_cycle_task(16'b0100000001000001, 1'b1);
		prog_cycle_task(16'b1100000001000001, 1'b0);
		prog_cycle_task(16'b0010000001000001, 1'b0);
		prog_cycle_task(16'b1010000001000001, 1'b0);
		prog_cycle_task(16'b0110000001000001, 1'b0);
		prog_cycle_task(16'b1110000001000001, 1'b1);
		prog_cycle_task(16'b0000010001000001, 1'b0);
		prog_cycle_task(16'b1000010001000001, 1'b0);
		prog_cycle_task(16'b0100010001000001, 1'b1);
		prog_cycle_task(16'b1100010001000001, 1'b0);
		prog_cycle_task(16'b0010010001000001, 1'b0);
		prog_cycle_task(16'b1010010001000001, 1'b0);
		prog_cycle_task(16'b0110010001000001, 1'b0);
		prog_cycle_task(16'b1110010001000001, 1'b1);
		prog_cycle_task(16'b0000001001000001, 1'b0);
		prog_cycle_task(16'b1000001001000001, 1'b0);
		prog_cycle_task(16'b0100001001000001, 1'b1);
		prog_cycle_task(16'b1100001001000001, 1'b0);
		prog_cycle_task(16'b0010001001000001, 1'b0);
		prog_cycle_task(16'b1010001001000001, 1'b0);
		prog_cycle_task(16'b0110001001000001, 1'b0);
		prog_cycle_task(16'b1110001001000001, 1'b1);
		prog_cycle_task(16'b0000011001000001, 1'b0);
		prog_cycle_task(16'b1000011001000001, 1'b0);
		prog_cycle_task(16'b0100011001000001, 1'b1);
		prog_cycle_task(16'b1100011001000001, 1'b0);
		prog_cycle_task(16'b0010011001000001, 1'b0);
		prog_cycle_task(16'b1010011001000001, 1'b0);
		prog_cycle_task(16'b0110011001000001, 1'b0);
		prog_cycle_task(16'b1110011001000001, 1'b1);
		prog_cycle_task(16'b0000000000000000, 1'b0);

// Port assign configuration
		`uvm_do_with(req,{req.address == 16'b0000000000000000; req.data_in == 1'b0; req.IE == 64'hFFFFFFFFFFFDFFFF;})


endtask;

`endif
