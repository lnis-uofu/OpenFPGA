// Benchmark "top" written by ABC on Thu Feb 21 17:22:32 2019

module elliptic ( clk, 
    tin_psv39_8_8_, tin_psv39_0_0_, tin_psv13_5_5_, tin_psv2_13_13_,
    tin_psv2_8_8_, pinp_2_2_, tin_psv38_2_2_, tin_psv33_5_5_,
    tin_psv26_6_6_, tin_psv2_9_9_, pinp_3_3_, tin_psv18_2_2_,
    tin_psv39_9_9_, tin_psv39_1_1_, tin_psv13_6_6_, tin_psv2_6_6_,
    pinp_0_0_, tin_psv38_3_3_, tin_psv33_6_6_, tin_psv26_13_13_,
    tin_psv26_12_12_, tin_psv26_7_7_, tin_psv2_7_7_, pinp_1_1_,
    preset_0_0_, tin_psv18_3_3_, tin_psv39_2_2_, tin_psv33_12_12_,
    tin_psv33_11_11_, tin_psv33_10_10_, tin_psv13_7_7_, tin_psv2_10_10_,
    tin_psv38_4_4_, tin_psv39_10_10_, tin_psv33_7_7_, tin_psv26_15_15_,
    tin_psv26_14_14_, tin_psv26_8_8_, tin_psv26_0_0_, tin_psv13_12_12_,
    tin_psv13_11_11_, tin_psv18_4_4_, tin_psv39_3_3_, tin_psv13_8_8_,
    tin_psv13_0_0_, pinp_15_15_, pinp_12_12_, tin_psv38_5_5_,
    tin_psv33_8_8_, tin_psv33_0_0_, tin_psv26_9_9_, tin_psv26_1_1_,
    tin_psv13_10_10_, tin_psv18_5_5_, tin_psv39_4_4_, tin_psv13_9_9_,
    tin_psv13_1_1_, tin_psv2_15_15_, tin_psv2_11_11_, tin_psv2_0_0_,
    tin_psv38_14_14_, tin_psv38_12_12_, tin_psv38_10_10_, tin_psv38_6_6_,
    tin_psv18_15_15_, tin_psv18_13_13_, tin_psv18_11_11_, tin_psv33_9_9_,
    tin_psv33_1_1_, tin_psv26_2_2_, tin_psv2_1_1_, pclk, tin_psv38_15_15_,
    tin_psv38_11_11_, tin_psv18_12_12_, tin_psv18_6_6_, tin_psv39_5_5_,
    tin_psv13_2_2_, pinp_14_14_, pinp_11_11_, pinp_8_8_, tin_psv38_7_7_,
    tin_psv39_12_12_, tin_psv39_11_11_, tin_psv33_2_2_, tin_psv26_3_3_,
    tin_psv13_14_14_, tin_psv13_13_13_, pinp_9_9_, tin_psv18_10_10_,
    tin_psv18_7_7_, tin_psv39_6_6_, tin_psv33_15_15_, tin_psv33_14_14_,
    tin_psv33_13_13_, tin_psv13_3_3_, tin_psv2_14_14_, tin_psv2_12_12_,
    tin_psv2_4_4_, pinp_6_6_, tin_psv38_8_8_, tin_psv38_0_0_,
    tin_psv39_14_14_, tin_psv39_13_13_, tin_psv33_3_3_, tin_psv26_11_11_,
    tin_psv26_10_10_, tin_psv26_4_4_, tin_psv13_15_15_, tin_psv2_5_5_,
    pinp_7_7_, tin_psv18_8_8_, tin_psv18_0_0_, tin_psv39_7_7_,
    tin_psv13_4_4_, tin_psv2_2_2_, pinp_13_13_, pinp_10_10_, pinp_4_4_,
    tin_psv38_9_9_, tin_psv38_1_1_, preset, tin_psv39_15_15_,
    tin_psv33_4_4_, tin_psv26_5_5_, tin_psv2_3_3_, pinp_5_5_,
    tin_psv38_13_13_, tin_psv18_14_14_, tin_psv18_9_9_, tin_psv18_1_1_,
    psv39_8_8_, psv39_0_0_, psv13_5_5_, psv2_13_13_, psv2_8_8_, psv38_2_2_,
    psv33_5_5_, psv26_6_6_, psv2_9_9_, psv18_2_2_, psv39_9_9_, psv39_1_1_,
    psv13_6_6_, psv2_6_6_, psv38_3_3_, psv33_6_6_, psv26_13_13_,
    psv26_12_12_, psv26_7_7_, psv2_7_7_, psv18_3_3_, psv39_2_2_,
    psv33_12_12_, psv33_11_11_, psv33_10_10_, psv13_7_7_, psv2_10_10_,
    psv38_4_4_, psv39_10_10_, psv33_7_7_, psv26_15_15_, psv26_14_14_,
    psv26_8_8_, psv26_0_0_, psv13_12_12_, psv13_11_11_, psv18_4_4_,
    psv39_3_3_, psv13_8_8_, psv13_0_0_, psv38_5_5_, psv33_8_8_, psv33_0_0_,
    psv26_9_9_, psv26_1_1_, psv13_10_10_, psv18_5_5_, psv39_4_4_,
    psv13_9_9_, psv13_1_1_, psv2_15_15_, psv2_11_11_, psv2_0_0_,
    psv38_14_14_, psv38_12_12_, psv38_10_10_, psv38_6_6_, psv18_15_15_,
    psv18_13_13_, psv18_11_11_, psv33_9_9_, psv33_1_1_, psv26_2_2_,
    psv2_1_1_, psv38_15_15_, psv38_11_11_, psv18_12_12_, psv18_6_6_,
    psv39_5_5_, psv13_2_2_, pover_0_0_, psv38_7_7_, psv39_12_12_,
    psv39_11_11_, psv33_2_2_, psv26_3_3_, psv13_14_14_, psv13_13_13_,
    psv18_10_10_, psv18_7_7_, psv39_6_6_, psv33_15_15_, psv33_14_14_,
    psv33_13_13_, psv13_3_3_, psv2_14_14_, psv2_12_12_, psv2_4_4_,
    psv38_8_8_, psv38_0_0_, pdn, psv39_14_14_, psv39_13_13_, psv33_3_3_,
    psv26_11_11_, psv26_10_10_, psv26_4_4_, psv13_15_15_, psv2_5_5_,
    psv18_8_8_, psv18_0_0_, psv39_7_7_, psv13_4_4_, psv2_2_2_, psv38_9_9_,
    psv38_1_1_, psv39_15_15_, psv33_4_4_, psv26_5_5_, psv2_3_3_,
    psv38_13_13_, psv18_14_14_, psv18_9_9_, psv18_1_1_  );
  input clk, tin_psv39_8_8_, tin_psv39_0_0_, tin_psv13_5_5_, tin_psv2_13_13_,
    tin_psv2_8_8_, pinp_2_2_, tin_psv38_2_2_, tin_psv33_5_5_,
    tin_psv26_6_6_, tin_psv2_9_9_, pinp_3_3_, tin_psv18_2_2_,
    tin_psv39_9_9_, tin_psv39_1_1_, tin_psv13_6_6_, tin_psv2_6_6_,
    pinp_0_0_, tin_psv38_3_3_, tin_psv33_6_6_, tin_psv26_13_13_,
    tin_psv26_12_12_, tin_psv26_7_7_, tin_psv2_7_7_, pinp_1_1_,
    preset_0_0_, tin_psv18_3_3_, tin_psv39_2_2_, tin_psv33_12_12_,
    tin_psv33_11_11_, tin_psv33_10_10_, tin_psv13_7_7_, tin_psv2_10_10_,
    tin_psv38_4_4_, tin_psv39_10_10_, tin_psv33_7_7_, tin_psv26_15_15_,
    tin_psv26_14_14_, tin_psv26_8_8_, tin_psv26_0_0_, tin_psv13_12_12_,
    tin_psv13_11_11_, tin_psv18_4_4_, tin_psv39_3_3_, tin_psv13_8_8_,
    tin_psv13_0_0_, pinp_15_15_, pinp_12_12_, tin_psv38_5_5_,
    tin_psv33_8_8_, tin_psv33_0_0_, tin_psv26_9_9_, tin_psv26_1_1_,
    tin_psv13_10_10_, tin_psv18_5_5_, tin_psv39_4_4_, tin_psv13_9_9_,
    tin_psv13_1_1_, tin_psv2_15_15_, tin_psv2_11_11_, tin_psv2_0_0_,
    tin_psv38_14_14_, tin_psv38_12_12_, tin_psv38_10_10_, tin_psv38_6_6_,
    tin_psv18_15_15_, tin_psv18_13_13_, tin_psv18_11_11_, tin_psv33_9_9_,
    tin_psv33_1_1_, tin_psv26_2_2_, tin_psv2_1_1_, pclk, tin_psv38_15_15_,
    tin_psv38_11_11_, tin_psv18_12_12_, tin_psv18_6_6_, tin_psv39_5_5_,
    tin_psv13_2_2_, pinp_14_14_, pinp_11_11_, pinp_8_8_, tin_psv38_7_7_,
    tin_psv39_12_12_, tin_psv39_11_11_, tin_psv33_2_2_, tin_psv26_3_3_,
    tin_psv13_14_14_, tin_psv13_13_13_, pinp_9_9_, tin_psv18_10_10_,
    tin_psv18_7_7_, tin_psv39_6_6_, tin_psv33_15_15_, tin_psv33_14_14_,
    tin_psv33_13_13_, tin_psv13_3_3_, tin_psv2_14_14_, tin_psv2_12_12_,
    tin_psv2_4_4_, pinp_6_6_, tin_psv38_8_8_, tin_psv38_0_0_,
    tin_psv39_14_14_, tin_psv39_13_13_, tin_psv33_3_3_, tin_psv26_11_11_,
    tin_psv26_10_10_, tin_psv26_4_4_, tin_psv13_15_15_, tin_psv2_5_5_,
    pinp_7_7_, tin_psv18_8_8_, tin_psv18_0_0_, tin_psv39_7_7_,
    tin_psv13_4_4_, tin_psv2_2_2_, pinp_13_13_, pinp_10_10_, pinp_4_4_,
    tin_psv38_9_9_, tin_psv38_1_1_, preset, tin_psv39_15_15_,
    tin_psv33_4_4_, tin_psv26_5_5_, tin_psv2_3_3_, pinp_5_5_,
    tin_psv38_13_13_, tin_psv18_14_14_, tin_psv18_9_9_, tin_psv18_1_1_;
  output psv39_8_8_, psv39_0_0_, psv13_5_5_, psv2_13_13_, psv2_8_8_,
    psv38_2_2_, psv33_5_5_, psv26_6_6_, psv2_9_9_, psv18_2_2_, psv39_9_9_,
    psv39_1_1_, psv13_6_6_, psv2_6_6_, psv38_3_3_, psv33_6_6_,
    psv26_13_13_, psv26_12_12_, psv26_7_7_, psv2_7_7_, psv18_3_3_,
    psv39_2_2_, psv33_12_12_, psv33_11_11_, psv33_10_10_, psv13_7_7_,
    psv2_10_10_, psv38_4_4_, psv39_10_10_, psv33_7_7_, psv26_15_15_,
    psv26_14_14_, psv26_8_8_, psv26_0_0_, psv13_12_12_, psv13_11_11_,
    psv18_4_4_, psv39_3_3_, psv13_8_8_, psv13_0_0_, psv38_5_5_, psv33_8_8_,
    psv33_0_0_, psv26_9_9_, psv26_1_1_, psv13_10_10_, psv18_5_5_,
    psv39_4_4_, psv13_9_9_, psv13_1_1_, psv2_15_15_, psv2_11_11_,
    psv2_0_0_, psv38_14_14_, psv38_12_12_, psv38_10_10_, psv38_6_6_,
    psv18_15_15_, psv18_13_13_, psv18_11_11_, psv33_9_9_, psv33_1_1_,
    psv26_2_2_, psv2_1_1_, psv38_15_15_, psv38_11_11_, psv18_12_12_,
    psv18_6_6_, psv39_5_5_, psv13_2_2_, pover_0_0_, psv38_7_7_,
    psv39_12_12_, psv39_11_11_, psv33_2_2_, psv26_3_3_, psv13_14_14_,
    psv13_13_13_, psv18_10_10_, psv18_7_7_, psv39_6_6_, psv33_15_15_,
    psv33_14_14_, psv33_13_13_, psv13_3_3_, psv2_14_14_, psv2_12_12_,
    psv2_4_4_, psv38_8_8_, psv38_0_0_, pdn, psv39_14_14_, psv39_13_13_,
    psv33_3_3_, psv26_11_11_, psv26_10_10_, psv26_4_4_, psv13_15_15_,
    psv2_5_5_, psv18_8_8_, psv18_0_0_, psv39_7_7_, psv13_4_4_, psv2_2_2_,
    psv38_9_9_, psv38_1_1_, psv39_15_15_, psv33_4_4_, psv26_5_5_,
    psv2_3_3_, psv38_13_13_, psv18_14_14_, psv18_9_9_, psv18_1_1_;
  reg n_n9280, n_n9172, n_n9260, n_n7726, n_n8270, n_n8196, n_n9150,
    n_n9267, n_n7779, n_n9503, n_n8150, n_n9401, n_n7341, n_n9180, n_n8592,
    n_n8871, n_n7252, n_n7271, n_n6991, n_n8557, n_n7707, n_n7552, ndn3_23,
    n_n9548, n_n9467, n_n8002, n_n6950, n_n8930, n_n7244, n_n7819, n_n8883,
    n_n7709, n_n9580, n_n9130, n_n9486, n_n9235, n_n7522, n_n7373, n_n9085,
    n_n9638, n_n7452, n_n8775, n_n7654, n_n8410, n_n8208, n_n8377, n_n7558,
    n_n7599, n_n8225, n_n8202, n_n7670, n_n7888, n_n7889, n_n8597, n_n8152,
    n_n8394, n_n7812, n_n7816, n_n9141, n_n7332, n_n8758, n_n7765, n_n7877,
    n_n7814, n_n9008, n_n7581, n_n7376, n_n7970, pover_0_0_, n_n8599,
    n_n8227, n_n9442, n_n9485, n_n7148, n_n9311, n_n9273, ndn3_9, n_n8613,
    n_n8533, n_n8699, n_n8609, n_n8308, n_n8655, n_n8981, n_n7583, n_n9198,
    n_n9602, n_n8786, n_n9598, n_n7738, n_n8573, n_n9473, n_n9000, n_n8001,
    n_n9554, n_n8508, n_n9635, n_n7190, n_n8702, n_n9106, n_n7409, n_n9437,
    n_n9052, n_n8647, n_n9265, n_n7179, ndn3_13, ndn3_17, ndn3_25, ndn3_29,
    n_n9539, n_n7953, n_n8488, nen3_22, n_n9438, n_n8132, n_n8661, n_n7759,
    n_n8333, n_n9399, n_n7798, n_n9434, n_n7910, n_n9528, n_n7850, n_n8251,
    n_n7937, n_n8482, n_n9290, n_n8007, n_n7556, n_n9064, n_n9398, n_n9412,
    n_n9361, n_n9304, n_n7651, n_n7712, n_n7735, n_n7934, n_n7811, n_n8053,
    n_n9015, n_n8066, n_n9518, n_n8091, n_n9257, n_n8175, n_n8491, n_n8114,
    n_n7951, n_n8913, n_n8035, n_n8631, n_n8243, n_n7857, ngfdn_3, n_n7791,
    n_n9175, n_n9588, n_n9049, n_n9483, n_n9410, n_n7691, n_n7740, n_n7602,
    n_n7783, n_n7948, n_n7054, n_n9343, n_n9400, nsr1_2, n_n9127, n_n8531,
    n_n9335, n_n7324, n_n9611, n_n8112, n_n9406, n_n9618, n_n9613, n_n9242,
    n_n7384, n_n8884, n_n7462, n_n7908, n_n8765, n_n7909, n_n7898, n_n9135,
    n_n8862, n_n8037, ndn3_18, ndn3_22, n_n8974, n_n7286, n_n9223, n_n7306,
    n_n9169, n_n9125, nen3_39, n_n8278, n_n9557, n_n7758, n_n9391, n_n8110,
    n_n9597, n_n8568, n_n7428, n_n7931, n_n7742, n_n7236, n_n8219, n_n9568,
    n_n9200, n_n8545, n_n7823, n_n8005, n_n8736, n_n9339, n_n8499, n_n8086,
    n_n7803, n_n7640, n_n9098, n_n7160, n_n7713, n_n9566, n_n7955, n_n8414,
    n_n8006, n_n9560, n_n8742, n_n7174, n_n8882, n_n7546, n_n8282, n_n8998,
    n_n7656, n_n9465, n_n9601, n_n8875, n_n7954, n_n8959, n_n8957, n_n8247,
    n_n8258, n_n7641, n_n8843, n_n9321, n_n7702, nsr3_23, n_n8199, n_n7983,
    n_n7217, n_n7821, n_n9489, n_n8348, n_n9408, n_n8445, n_n9501, n_n7831,
    n_n7757, n_n9174, n_n9432, n_n8678, n_n8024, n_n7806, n_n8996, n_n7918,
    n_n8260, n_n9341, n_n9189, n_n9096, ndn3_30, n_n7775, n_n7693, nen3_16,
    n_n7643, n_n8941, n_n8042, n_n8681, n_n8659, n_n9110, n_n9573, n_n8951,
    n_n9589, n_n9387, n_n8279, n_n7790, n_n8406, n_n8582, n_n7911, n_n7474,
    n_n8466, n_n6984, n_n7760, n_n7847, n_n9559, n_n7362, n_n9300, n_n9550,
    n_n9492, n_n8777, n_n7764, n_n7826, n_n7777, n_n7824, n_n8173, n_n7498,
    n_n9148, n_n8753, n_n8772, n_n8049, n_n9362, ndn1_4, n_n9561, n_n9004,
    n_n8203, n_n8153, n_n9263, n_n8369, n_n9331, n_n7454, ndn3_7, n_n7527,
    n_n9036, n_n7875, n_n8697, n_n9497, n_n7291, nsr3_13, nsr3_38, n_n8240,
    n_n7703, n_n9282, n_n8237, n_n8935, n_n9244, n_n8648, n_n8235, n_n8611,
    n_n9045, n_n9334, n_n8572, n_n9491, n_n9134, n_n9555, n_n9336, n_n7050,
    n_n9346, n_n7140, n_n7681, n_n6948, n_n8549, ndn3_19, ndn3_28, n_n7102,
    n_n8093, n_n9041, n_n8381, n_n8810, nen3_36, n_n9047, n_n9333, n_n7736,
    n_n7820, n_n8986, n_n8891, n_n8000, n_n7968, n_n8750, n_n9558, n_n9368,
    n_n8519, n_n6956, n_n8298, n_n9397, n_n7017, n_n8638, n_n9552, n_n8964,
    n_n8016, n_n7603, n_n7696, n_n8589, n_n9337, n_n9132, n_n8652, n_n8707,
    n_n9407, n_n9044, n_n8808, nsr3_30, n_n8274, n_n8615, n_n8238, n_n7854,
    n_n8649, n_n8236, n_n8269, n_n9592, n_n8022, n_n8744, n_n8529, n_n7967,
    n_n9487, n_n8685, n_n9531, n_n9510, n_n7771, n_n8480, n_n8543, n_n7789,
    ndn3_11, ndn3_15, ndn3_21, n_n7584, n_n8354, n_n6952, n_n8864, n_n7930,
    n_n7962, n_n7929, n_n9316, n_n9102, n_n7308, n_n7657, n_n9264, n_n8760,
    n_n6912, n_n7887, n_n8911, n_n7952, n_n8704, n_n7876, n_n9596, n_n8430,
    n_n9019, n_n7699, n_n7375, n_n7936, n_n8340, n_n8809, n_n6961, n_n9429,
    n_n7743, n_n8980, n_n7582, n_n8968, n_n9371, n_n8741, n_n9502, n_n9373,
    n_n9248, n_n7822, n_n9054, n_n8273, n_n6937, n_n9342, n_n9325, n_n9609,
    n_n9623, n_n9470, n_n7570, n_n9310, n_n9366, n_n7181, n_n8739, n_n8939,
    n_n7256, n_n8983, n_n7487, n_n9268, n_n8906, n_n7988, n_n9181, n_n8725,
    n_n8626, ndn3_27, n_n8210, n_n7415, n_n8900, nen3_19, n_n8762, n_n8512,
    n_n8095, n_n8982, n_n7387, n_n9494, n_n7689, n_n7835, n_n9157, n_n8552,
    n_n7381, n_n9446, n_n8633, n_n7684, n_n7310, n_n8402, n_n9315, n_n7950,
    n_n8504, n_n8456, n_n7514, n_n7315, n_n9476, n_n8276, n_n8833, n_n7923,
    n_n9395, n_n9512, n_n9319, nsr3_35, n_n7154, n_n9495, n_n9137, n_n8854,
    n_n9183, n_n9323, n_n9349, n_n7896, n_n8073, n_n8970, n_n9314, n_n8486,
    n_n7246, n_n7866, n_n9599, n_n7635, n_n8984, n_n7360, n_n8794, n_n9108,
    n_n9286, ndn3_12, ndn3_16, n_n7708, n_n7807, n_n7650, n_n7947, n_n9500,
    n_n7734, n_n8464, n_n7659, n_n7630, n_n7756, n_n8691, n_n9176, n_n9327,
    n_n7995, n_n7395, n_n7878, n_n7507, n_n7959, n_n7825, n_n8009, n_n8281,
    n_n7685, n_n8106, n_n7687, n_n7766, n_n7880, n_n8961, n_n8014, n_n9278,
    n_n9087, n_n9182, n_n7852, n_n9324, nak3_13, n_n9416, nsr3_14, n_n8603,
    n_n7026, n_n8856, n_n8272, n_n9312, n_n7985, n_n8312, n_n7231, n_n9396,
    n_n8801, n_n8683, ndn3_39, n_n8245, n_n9458, n_n9302, n_n7392, n_n6963,
    n_n7808, n_n7225, n_n7817, n_n8201, n_n7793, n_n8177, n_n8389, n_n9440,
    n_n7683, n_n7761, n_n7667, n_n7980, n_n7509, n_n7813, n_n8396, n_n9535,
    n_n7209, n_n7003, n_n7695, n_n7624, n_n8791, n_n7374, n_n7429, n_n7944,
    n_n9266, n_n8100, n_n6988, n_n6986, n_n8933, n_n7117, n_n9043, n_n8241,
    n_n9219, n_n8198, n_n8081, n_n8575, n_n8710, n_n7622, n_n7966, n_n7885,
    n_n7033, ndn3_34, n_n9186, ndn3_50, n_n7879, n_n7019, n_n9171, n_n7261,
    n_n8223, n_n8989, n_n7993, n_n7845, n_n8253, n_n8889, n_n7809, n_n8918,
    n_n8515, n_n7933, n_n8075, n_n7338, n_n8104, n_n8171, n_n9059, n_n9023,
    n_n7692, n_n9441, n_n6920, n_n8831, n_n8441, n_n9576, n_n9252, n_n9363,
    ndn3_4, n_n9247, n_n7561, n_n8923, n_n7978, n_n8978, n_n9499, n_n8713,
    n_n8944, n_n8239, n_n7652, n_n9042, n_n8530, n_n9271, n_n9318, n_n7706,
    n_n7964, n_n8222, n_n8898, n_n7976, n_n7649, n_n7604, n_n7961, n_n7424,
    n_n7476, n_n9259, n_n9309, n_n9161, n_n8436, n_n9121, n_n8061, n_n8004,
    n_n9360, n_n9205, n_n8392, n_n9034, n_n8375, n_n8328, n_n9298, n_n7598,
    n_n8506, pdn, n_n7737, n_n7420, n_n9291, n_n7946, n_n8584, n_n9308,
    n_n9403, n_n7284, n_n9270, n_n7390, n_n9351, n_n6968, n_n8668, n_n9605,
    n_n7013, n_n9626, n_n8200, n_n9028, n_n8803, n_n9570, n_n8366, n_n9050,
    n_n8650, n_n8574, n_n7276, n_n9212, n_n8384, ndn3_35, n_n8449, ndn3_46,
    n_n7554, n_n8743, n_n8277, n_n9359, n_n8425, n_n9104, n_n9221, n_n9448,
    n_n9537, n_n8003, n_n7467, n_n8233, n_n7932, n_n8064, n_n9162, n_n7971,
    n_n8055, n_n7711, n_n8256, n_n7925, n_n7762, n_n7668, n_n7914, n_n7873,
    n_n7849, n_n9421, n_n7626, n_n7848, n_n8263, n_n9100, n_n9393, n_n9591,
    n_n7588, n_n9123, n_n9159, n_n9128, n_n8045, n_n7728, n_n8929, n_n7739,
    n_n9355, n_n9394, n_n8470, n_n8571, n_n8796, ndn3_36, n_n7990, n_n8781,
    n_n8817, n_n9160, n_n9092, n_n8513, n_n8213, n_n8581, n_n9284, n_n7837,
    n_n8224, n_n9203, n_n7655, n_n8946, n_n7052, n_n9615, n_n8473, n_n7741,
    n_n9460, n_n7912, n_n7606, n_n9021, n_n7781, n_n7810, n_n7108, n_n7697,
    n_n7642, n_n9595, n_n7694, n_n8221, n_n7600, n_n7935, n_n9230, n_n7701,
    n_n7510, n_n7627, n_n8502, n_n8516, n_n7913, n_n9320, n_n7411, n_n9129,
    n_n9053, n_n7069, n_n8617, n_n7242, n_n8230, n_n9294, n_n8249, n_n8972,
    n_n7074, n_n7493, n_n8290, n_n8821, n_n7769, n_n7491, n_n9600, n_n9317,
    n_n8047, n_n9629, n_n9126, n_n9508, n_n9155, n_n8528, ndn3_37, ndn3_42,
    n_n9358, n_n8185, nen3_28, n_n8839, n_n7903, n_n9139, n_n9075, n_n9439,
    n_n9353, n_n7665, n_n8798, n_n7146, n_n7890, n_n7176, n_n8477, n_n8514,
    n_n8636, n_n7183, n_n8657, n_n9493, n_n7969, n_n9255, n_n8535, n_n8619,
    n_n8909, n_n7744, n_n9119, n_n7827, n_n8916, n_n8729, n_n9011, n_n8779,
    n_n6980, n_n7715, n_n9067, n_n9164, n_n7402, n_n8938, n_n9046, n_n8789,
    n_n9390, n_n7768, n_n9136, n_n8670, n_n8644, n_n9178, n_n8188, n_n7083,
    n_n9344, n_n7366, n_n8361, n_n9228, n_n9402, n_n8510, n_n8881, n_n9404,
    n_n9424, n_n9031, nsr3_37, n_n8197, n_n8468, n_n7121, n_n7511, ndn3_44,
    n_n9322, n_n7682, n_n9603, nlc1_2, n_n8408, n_n8577, n_n7079, n_n8828,
    n_n9340, n_n8586, n_n7901, n_n8628, n_n8869, n_n7710, n_n8993, n_n9586,
    n_n8852, n_n8583, n_n8011, n_n7717, n_n8326, n_n9163, n_n8344, n_n8296,
    n_n8116, n_n8267, n_n7686, n_n9061, n_n9338, n_n7688, n_n9081, n_n6910,
    n_n8727, n_n7674, n_n7330, n_n8966, n_n7843, n_n8847, n_n9376, n_n7553,
    n_n9292, n_n7464, n_n8146, n_n8439, n_n9498, n_n8118, n_n9452, n_n9239,
    n_n9237, n_n9488, ndn3_2, n_n9522, n_n9313, n_n7435, n_n8665, n_n9593,
    n_n8303, n_n7022, n_n9173, n_n9261, n_n7150, n_n9455, n_n8371, nsr3_20,
    n_n8271, n_n9542, n_n7444, ndn3_40, n_n7130, n_n9347, n_n8102, n_n9225,
    n_n8462, n_n8088, n_n9026, n_n9289, n_n7661, n_n8108, n_n8921, n_n7859,
    n_n7732, n_n7956, n_n9520, n_n7666, n_n7678, n_n7846, n_n8280, n_n8841,
    n_n7336, n_n8226, n_n8151, n_n7644, n_n8770, n_n8423, n_n7763, n_n9525,
    n_n8033, n_n7881, n_n7815, n_n9232, n_n7792, n_n9563, n_n8672, n_n7346,
    n_n7949, n_n8756, n_n8641, n_n8192, n_n8058, n_n8561, n_n9306, n_n9165,
    n_n8850, n_n9210, ndn2_2, n_n7342, n_n8051, n_n7136, n_n9348, n_n9006,
    n_n7653, n_n7905, n_n9166, n_n7065, n_n9490, n_n7024, n_n7586, n_n8416,
    n_n8937, n_n8141, n_n7853, n_n8121, n_n9604, n_n9496, n_n8195, n_n9516,
    n_n9077, n_n9436, n_n9051, n_n7664, n_n8419, n_n7874, n_n9133, n_n9392,
    n_n7770, ndn3_32, n_n7601, n_n8206, n_n7927, n_n9606, n_n7111, n_n9269,
    ndn3_38, n_n7886, n_n9179, n_n9357, n_n9594, n_n7628, n_n8454, ndn3_20,
    n_n9505, nen3_34, n_n9632, n_n7076, n_n9262, n_n9048, n_n9578, n_n8135,
    ndn3_26, n_n7500, n_n6974, n_n8605, n_n9296, n_n7156, n_n7920, n_n8895,
    n_n8991, n_n8139, n_n9275, n_n7203, n_n9590, n_n7344, n_n6976, n_n7629,
    ndn3_14, n_n7862, n_n9013, n_n7288, n_n8078, n_n7334, n_n7704, n_n7788,
    n_n8526, n_n9556, n_n9345, n_n8447, n_n7485, n_n8570, n_n7453, n_n7928,
    n_n8646, n_n9405, n_n8948, n_n9131, n_n8216, n_n9177, n_n7844, n_n8811,
    n_n9145, n_n8428, n_n8858, n_n8580;
  wire n4845, n4846, n4847, n4848, n4849_1, n4850, n4851, n4852, n4853,
    n4854_1, n4855, n4856, n4857, n4858, n4859_1, n4860, n4861, n4862,
    n4863, n4864_1, n4865, n4866, n4867, n4868, n4869_1, n4870, n4871,
    n4872, n4873, n4874_1, n4875, n4876, n4877, n4878, n4879_1, n4880,
    n4881, n4882, n4883, n4884_1, n4885, n4886, n4887, n4888, n4889_1,
    n4890, n4891, n4892, n4893, n4894_1, n4895, n4896, n4897, n4898,
    n4899_1, n4900, n4901, n4902, n4903, n4904_1, n4905, n4906, n4907,
    n4908, n4909_1, n4910, n4911, n4912, n4913, n4914_1, n4915, n4916,
    n4917, n4918, n4919_1, n4920, n4921, n4922, n4923, n4924_1, n4925,
    n4926, n4927, n4928, n4929_1, n4930, n4931, n4932, n4933, n4934_1,
    n4935, n4936, n4937, n4938, n4939_1, n4940, n4941, n4942, n4943,
    n4944_1, n4945, n4946, n4947, n4948, n4949_1, n4950, n4951, n4952,
    n4953, n4954_1, n4955, n4956, n4957, n4958, n4959_1, n4960, n4961,
    n4962, n4963, n4964_1, n4965, n4966, n4967, n4968, n4969_1, n4970,
    n4971, n4972, n4973, n4974_1, n4975, n4976, n4977, n4978, n4979_1,
    n4980, n4981, n4982, n4983, n4984_1, n4985, n4986, n4987, n4988,
    n4989_1, n4990, n4991, n4992, n4993, n4994_1, n4995, n4996, n4997,
    n4998, n4999_1, n5000, n5001, n5002, n5003, n5004_1, n5005, n5006,
    n5007, n5008, n5009_1, n5010, n5011, n5012, n5013, n5014_1, n5015,
    n5016, n5017, n5018, n5019_1, n5020, n5021, n5022, n5023, n5024_1,
    n5025, n5026, n5027, n5028, n5029_1, n5030, n5031, n5032, n5033,
    n5034_1, n5035, n5036, n5037, n5038, n5039_1, n5040, n5041, n5042,
    n5043, n5044_1, n5045, n5046, n5047, n5048, n5049_1, n5050, n5051,
    n5052, n5053, n5054_1, n5055, n5056, n5057, n5058, n5059_1, n5060,
    n5061, n5062, n5063, n5064_1, n5065, n5066, n5067, n5068, n5069_1,
    n5070, n5071, n5072, n5073, n5074_1, n5075, n5076, n5077, n5078,
    n5079_1, n5080, n5081, n5082, n5083, n5084_1, n5085, n5086, n5087,
    n5088, n5089_1, n5090, n5091, n5092, n5093, n5094_1, n5095, n5096,
    n5097, n5098, n5099_1, n5100, n5101, n5102, n5103, n5104_1, n5105,
    n5106, n5107, n5108, n5109_1, n5110, n5111, n5112, n5113, n5114_1,
    n5115, n5116, n5117, n5118, n5119_1, n5120, n5121, n5122, n5123,
    n5124_1, n5125, n5126, n5127, n5128, n5129_1, n5130, n5131, n5132,
    n5133, n5134_1, n5135, n5136, n5137, n5138, n5139_1, n5140, n5141,
    n5142, n5143, n5144_1, n5145, n5146, n5147, n5148, n5149_1, n5150,
    n5151, n5152, n5153, n5154_1, n5155, n5156, n5157, n5158, n5159_1,
    n5160, n5161, n5162, n5163, n5164_1, n5165, n5166, n5167, n5168,
    n5169_1, n5170, n5171, n5172, n5173, n5174_1, n5175, n5176, n5177,
    n5178, n5179_1, n5180, n5181, n5182, n5183, n5184_1, n5185, n5186,
    n5187, n5188, n5189_1, n5190, n5191, n5192, n5193, n5194_1, n5195,
    n5196, n5197, n5198, n5199_1, n5200, n5201, n5202, n5203, n5204_1,
    n5205, n5206, n5207, n5208, n5209_1, n5210, n5211, n5212, n5213,
    n5214_1, n5215, n5216, n5217, n5218, n5219_1, n5220, n5221, n5222,
    n5223, n5224_1, n5225, n5226, n5227, n5228, n5229_1, n5230, n5231,
    n5232, n5233, n5234_1, n5235, n5236, n5237, n5238, n5239_1, n5240,
    n5241, n5242, n5243, n5244_1, n5245, n5246, n5247, n5248, n5249_1,
    n5250, n5251, n5252, n5253, n5254_1, n5255, n5256, n5257, n5258,
    n5259_1, n5260, n5261, n5262, n5263, n5264_1, n5265, n5266, n5267,
    n5268, n5269_1, n5270, n5271, n5272, n5273, n5274_1, n5275, n5276,
    n5277, n5278, n5279_1, n5280, n5281, n5282, n5283, n5284_1, n5285,
    n5286, n5287, n5288, n5289_1, n5290, n5291, n5292, n5293, n5294_1,
    n5295, n5296, n5297, n5298, n5299_1, n5300, n5301, n5302, n5303,
    n5304_1, n5305, n5306, n5307, n5308, n5309_1, n5310, n5311, n5312,
    n5313, n5314_1, n5315, n5316, n5317, n5318, n5319_1, n5320, n5321,
    n5322, n5323, n5324_1, n5325, n5326, n5327, n5328, n5329_1, n5330,
    n5331, n5332, n5333, n5334_1, n5335, n5336, n5337, n5338, n5339_1,
    n5340, n5341, n5342, n5343, n5344_1, n5345, n5346, n5347, n5348,
    n5349_1, n5350, n5351, n5352, n5353, n5354_1, n5355, n5356, n5357,
    n5358, n5359_1, n5360, n5361, n5362, n5363, n5364_1, n5365, n5366,
    n5367, n5368, n5369_1, n5370, n5371, n5372, n5373, n5374_1, n5375,
    n5376, n5377, n5378, n5379_1, n5380, n5381, n5382, n5383, n5384_1,
    n5385, n5386, n5387, n5388, n5389_1, n5390, n5391, n5392, n5393,
    n5394_1, n5395, n5396, n5397, n5398, n5399_1, n5400, n5401, n5402,
    n5403, n5404_1, n5405, n5406, n5407, n5408, n5409_1, n5410, n5411,
    n5412, n5413, n5414_1, n5415, n5416, n5417, n5418, n5419_1, n5420,
    n5421, n5422, n5423, n5424_1, n5425, n5426, n5427, n5428, n5429_1,
    n5430, n5431, n5432, n5433, n5434_1, n5435, n5436, n5437, n5438,
    n5439_1, n5440, n5441, n5442, n5443, n5444_1, n5445, n5446, n5447,
    n5448, n5449_1, n5450, n5451, n5452, n5453, n5454_1, n5455, n5456,
    n5457, n5458, n5459_1, n5460, n5461, n5462, n5463, n5464_1, n5465,
    n5466, n5467, n5468, n5469_1, n5470, n5471, n5472, n5473, n5474_1,
    n5475, n5476, n5477, n5478, n5479_1, n5480, n5481, n5482, n5483,
    n5484_1, n5485, n5486, n5487, n5488, n5489_1, n5490, n5491, n5492,
    n5493, n5494_1, n5495, n5496, n5497, n5498, n5499_1, n5500, n5501,
    n5502, n5503, n5504_1, n5505, n5506, n5507, n5508, n5509_1, n5510,
    n5511, n5512, n5513, n5514_1, n5515, n5516, n5517, n5518, n5519_1,
    n5520, n5521, n5522, n5523, n5524_1, n5525, n5526, n5527, n5528,
    n5529_1, n5530, n5531, n5532, n5533, n5534_1, n5535, n5536, n5537,
    n5538, n5539_1, n5540, n5541, n5542, n5543, n5544_1, n5545, n5546,
    n5547, n5548, n5549_1, n5550, n5551, n5552, n5553, n5554_1, n5555,
    n5556, n5557, n5558, n5559_1, n5560, n5561, n5562, n5563, n5564_1,
    n5565, n5566, n5567, n5568, n5569_1, n5570, n5571, n5572, n5573,
    n5574_1, n5575, n5576, n5577, n5578, n5579_1, n5580, n5581, n5582,
    n5583, n5584_1, n5585, n5586, n5587, n5588, n5589_1, n5590, n5591,
    n5592, n5593, n5594_1, n5595, n5596, n5597, n5598, n5599_1, n5600,
    n5601, n5602, n5603, n5604_1, n5605, n5606, n5607, n5608, n5609_1,
    n5610, n5611, n5612, n5613, n5614_1, n5615, n5616, n5617, n5618,
    n5619_1, n5620, n5621, n5622, n5623, n5624_1, n5625, n5626, n5627,
    n5628, n5629_1, n5630, n5631, n5632, n5633, n5634_1, n5635, n5636,
    n5637, n5638, n5639_1, n5640, n5641, n5642, n5643, n5644_1, n5645,
    n5646, n5647, n5648, n5649_1, n5650, n5651, n5652, n5653, n5654_1,
    n5655, n5656, n5657, n5658, n5659_1, n5660, n5661, n5662, n5663,
    n5664_1, n5665, n5666, n5667, n5668, n5669_1, n5670, n5671, n5672,
    n5673, n5674_1, n5675, n5676, n5677, n5678, n5679_1, n5680, n5681,
    n5682, n5683, n5684_1, n5685, n5686, n5687, n5688, n5689_1, n5690,
    n5691, n5692, n5693, n5694_1, n5695, n5696, n5697, n5698, n5699_1,
    n5700, n5701, n5702, n5703, n5704_1, n5705, n5706, n5707, n5708,
    n5709_1, n5710, n5711, n5712, n5713, n5714_1, n5715, n5716, n5717,
    n5718, n5719_1, n5720, n5721, n5722, n5723, n5724_1, n5725, n5726,
    n5727, n5728, n5729_1, n5730, n5731, n5732, n5733, n5734_1, n5735,
    n5736, n5737, n5738, n5739_1, n5740, n5741, n5742, n5743, n5744_1,
    n5745, n5746, n5747, n5748, n5749_1, n5750, n5751, n5752, n5753,
    n5754_1, n5755, n5756, n5757, n5758, n5759_1, n5760, n5761, n5762,
    n5763, n5764_1, n5765, n5766, n5767, n5768, n5769_1, n5770, n5771,
    n5772, n5773, n5774_1, n5775, n5776, n5777, n5778, n5779_1, n5780,
    n5781, n5782, n5783, n5784_1, n5785, n5786, n5787, n5788, n5789_1,
    n5790, n5791, n5792, n5793, n5794_1, n5795, n5796, n5797, n5798,
    n5799_1, n5800, n5801, n5802, n5803, n5804_1, n5805, n5806, n5807,
    n5808, n5809_1, n5810, n5811, n5812, n5813, n5814_1, n5815, n5816,
    n5817, n5818, n5819_1, n5820, n5821, n5822, n5823, n5824_1, n5825,
    n5826, n5827, n5828, n5829_1, n5830, n5831, n5832, n5833, n5834_1,
    n5835, n5836, n5837, n5838, n5839_1, n5840, n5841, n5842, n5843,
    n5844_1, n5845, n5846, n5847, n5848, n5849_1, n5850, n5851, n5852,
    n5853, n5854_1, n5855, n5856, n5857, n5858, n5859_1, n5860, n5861,
    n5862, n5863, n5864_1, n5865, n5866, n5867, n5868, n5869_1, n5870,
    n5871, n5872, n5873, n5874_1, n5875, n5876, n5877, n5878, n5879_1,
    n5880, n5881, n5882, n5883, n5884_1, n5885, n5886, n5887, n5888,
    n5889_1, n5890, n5891, n5892, n5893, n5894_1, n5895, n5896, n5897,
    n5898, n5899_1, n5900, n5901, n5902, n5903, n5904_1, n5905, n5906,
    n5907, n5908, n5909_1, n5910, n5911, n5912, n5913, n5914_1, n5915,
    n5916, n5917, n5918, n5919_1, n5920, n5921, n5922, n5923, n5924_1,
    n5925, n5926, n5927, n5928, n5929_1, n5930, n5931, n5932, n5933,
    n5934_1, n5935, n5936, n5937, n5938, n5939_1, n5940, n5941, n5942,
    n5943, n5944_1, n5945, n5946, n5947, n5948, n5949_1, n5950, n5951,
    n5952, n5953, n5954_1, n5955, n5956, n5957, n5958, n5959_1, n5960,
    n5961, n5962, n5963, n5964_1, n5965, n5966, n5967, n5968, n5969_1,
    n5970, n5971, n5972, n5973, n5974_1, n5975, n5976, n5977, n5978,
    n5979_1, n5980, n5981, n5982, n5983, n5984_1, n5985, n5986, n5987,
    n5988, n5989_1, n5990, n5991, n5992, n5993, n5994_1, n5995, n5996,
    n5997, n5998, n5999_1, n6000, n6001, n6002, n6003, n6004_1, n6005,
    n6006, n6007, n6008, n6009_1, n6010, n6011, n6012, n6013, n6014_1,
    n6015, n6016, n6017, n6018, n6019_1, n6020, n6021, n6022, n6023,
    n6024_1, n6025, n6026, n6027, n6028, n6029_1, n6030, n6031, n6032,
    n6033, n6034_1, n6035, n6036, n6037, n6038, n6039_1, n6040, n6041,
    n6042, n6043, n6044_1, n6045, n6046, n6047, n6048, n6049_1, n6050,
    n6051, n6052, n6053, n6054_1, n6055, n6056, n6057, n6058, n6059_1,
    n6060, n6061, n6062, n6063, n6064_1, n6065, n6066, n6067, n6068,
    n6069_1, n6070, n6071, n6072, n6073, n6074_1, n6075, n6076, n6077,
    n6078, n6079_1, n6080, n6081, n6082, n6083, n6084_1, n6085, n6086,
    n6087, n6088, n6089_1, n6090, n6091, n6092, n6093, n6094_1, n6095,
    n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
    n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
    n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
    n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
    n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
    n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
    n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
    n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
    n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
    n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
    n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
    n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
    n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
    n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
    n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
    n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
    n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
    n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
    n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
    n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
    n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
    n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
    n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
    n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
    n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
    n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
    n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
    n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
    n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
    n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
    n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
    n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
    n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
    n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
    n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
    n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
    n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
    n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
    n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
    n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
    n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
    n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
    n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
    n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
    n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
    n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
    n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
    n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
    n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
    n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
    n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
    n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
    n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
    n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
    n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
    n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
    n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
    n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
    n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
    n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
    n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
    n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
    n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
    n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
    n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
    n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
    n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
    n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
    n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
    n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
    n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
    n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
    n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
    n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
    n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
    n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
    n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
    n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
    n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
    n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
    n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
    n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
    n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
    n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
    n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
    n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
    n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
    n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
    n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
    n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
    n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
    n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
    n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
    n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
    n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
    n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
    n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
    n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
    n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
    n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
    n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
    n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
    n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
    n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
    n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
    n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
    n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
    n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
    n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
    n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
    n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
    n7206, n7207, n7208, n7209, n7210, n7211, n7212, n491, n496, n501,
    n506, n511, n516, n521, n526, n531, n536, n541, n546, n551, n556, n561,
    n566, n571, n576, n581, n586, n591, n596, n601, n606, n611, n616, n621,
    n626, n631, n636, n641, n646, n651, n656, n661, n666, n671, n676, n681,
    n686, n691, n696, n701, n706, n711, n716, n721, n726, n731, n736, n741,
    n746, n751, n756, n761, n766, n771, n776, n781, n786, n791, n796, n801,
    n806, n811, n816, n821, n826, n831, n835, n840, n845, n850, n855, n860,
    n865, n870, n875, n880, n885, n890, n895, n900, n905, n910, n915, n920,
    n925, n930, n935, n940, n945, n950, n955, n960, n965, n970, n975, n980,
    n985, n990, n995, n1000, n1005, n1010, n1015, n1020, n1025, n1030,
    n1035, n1040, n1045, n1050, n1055, n1060, n1065, n1070, n1075, n1080,
    n1085, n1090, n1095, n1100, n1105, n1110, n1115, n1120, n1125, n1130,
    n1135, n1140, n1145, n1150, n1155, n1160, n1165, n1170, n1175, n1180,
    n1185, n1190, n1195, n1200, n1205, n1210, n1215, n1220, n1225, n1230,
    n1235, n1240, n1245, n1250, n1255, n1260, n1265, n1270, n1275, n1280,
    n1285, n1290, n1295, n1300, n1305, n1310, n1315, n1320, n1325, n1330,
    n1335, n1340, n1345, n1350, n1355, n1360, n1365, n1370, n1375, n1380,
    n1385, n1390, n1395, n1400, n1405, n1410, n1415, n1420, n1425, n1430,
    n1435, n1440, n1445, n1450, n1455, n1460, n1465, n1470, n1475, n1480,
    n1485, n1490, n1495, n1500, n1505, n1510, n1515, n1520, n1525, n1530,
    n1535, n1540, n1545, n1550, n1555, n1560, n1565, n1570, n1575, n1580,
    n1585, n1590, n1595, n1600, n1605, n1610, n1615, n1620, n1625, n1630,
    n1635, n1640, n1645, n1650, n1655, n1660, n1665, n1670, n1675, n1680,
    n1685, n1690, n1695, n1700, n1705, n1710, n1715, n1720, n1725, n1730,
    n1735, n1740, n1745, n1750, n1755, n1760, n1765, n1770, n1775, n1780,
    n1785, n1790, n1795, n1800, n1805, n1810, n1815, n1820, n1825, n1830,
    n1835, n1840, n1845, n1850, n1855, n1860, n1865, n1870, n1875, n1880,
    n1885, n1890, n1895, n1900, n1905, n1910, n1915, n1920, n1925, n1930,
    n1935, n1940, n1945, n1950, n1955, n1960, n1965, n1970, n1975, n1980,
    n1985, n1990, n1995, n2000, n2005, n2010, n2015, n2020, n2025, n2030,
    n2035, n2040, n2045, n2050, n2055, n2060, n2065, n2070, n2075, n2080,
    n2085, n2090, n2095, n2100, n2105, n2110, n2115, n2120, n2125, n2130,
    n2135, n2140, n2145, n2150, n2155, n2160, n2165, n2170, n2175, n2180,
    n2185, n2190, n2195, n2200, n2205, n2210, n2215, n2220, n2225, n2230,
    n2235, n2240, n2245, n2250, n2255, n2260, n2265, n2270, n2275, n2280,
    n2285, n2290, n2295, n2300, n2305, n2310, n2315, n2320, n2325, n2330,
    n2335, n2340, n2345, n2350, n2355, n2360, n2365, n2370, n2375, n2380,
    n2385, n2390, n2395, n2400, n2405, n2410, n2415, n2420, n2425, n2430,
    n2435, n2440, n2445, n2450, n2455, n2460, n2465, n2470, n2475, n2480,
    n2485, n2490, n2495, n2500, n2505, n2510, n2515, n2520, n2525, n2530,
    n2535, n2540, n2545, n2550, n2555, n2560, n2565, n2570, n2575, n2580,
    n2585, n2590, n2595, n2600, n2605, n2610, n2615, n2620, n2625, n2630,
    n2635, n2640, n2645, n2650, n2655, n2660, n2665, n2670, n2675, n2680,
    n2685, n2690, n2695, n2700, n2705, n2710, n2715, n2720, n2725, n2730,
    n2735, n2740, n2745, n2750, n2755, n2760, n2765, n2770, n2775, n2780,
    n2785, n2790, n2795, n2800, n2805, n2810, n2815, n2820, n2825, n2830,
    n2835, n2840, n2845, n2850, n2855, n2860, n2865, n2870, n2875, n2880,
    n2885, n2890, n2895, n2900, n2905, n2910, n2915, n2920, n2925, n2930,
    n2935, n2940, n2945, n2950, n2955, n2960, n2965, n2970, n2975, n2980,
    n2985, n2990, n2995, n3000, n3005, n3010, n3015, n3020, n3025, n3030,
    n3035, n3040, n3045, n3050, n3055, n3060, n3065, n3070, n3075, n3080,
    n3085, n3090, n3095, n3100, n3105, n3110, n3115, n3120, n3125, n3130,
    n3135, n3140, n3145, n3150, n3155, n3160, n3165, n3170, n3175, n3180,
    n3185, n3190, n3195, n3200, n3205, n3210, n3215, n3220, n3225, n3230,
    n3235, n3240, n3245, n3250, n3255, n3260, n3265, n3270, n3275, n3280,
    n3285, n3290, n3295, n3300, n3305, n3310, n3315, n3320, n3325, n3330,
    n3335, n3340, n3345, n3350, n3355, n3360, n3365, n3370, n3375, n3380,
    n3385, n3390, n3395, n3400, n3405, n3410, n3415, n3420, n3425, n3430,
    n3435, n3440, n3445, n3450, n3455, n3460, n3465, n3470, n3475, n3480,
    n3485, n3490, n3495, n3500, n3505, n3510, n3515, n3520, n3525, n3530,
    n3535, n3540, n3545, n3550, n3555, n3560, n3565, n3570, n3575, n3580,
    n3585, n3590, n3595, n3600, n3605, n3610, n3615, n3620, n3625, n3630,
    n3635, n3640, n3645, n3650, n3655, n3660, n3665, n3670, n3675, n3680,
    n3685, n3690, n3695, n3700, n3705, n3710, n3715, n3720, n3725, n3730,
    n3735, n3740, n3745, n3750, n3755, n3760, n3765, n3770, n3775, n3780,
    n3785, n3790, n3795, n3800, n3805, n3810, n3815, n3820, n3825, n3830,
    n3835, n3840, n3845, n3850, n3855, n3860, n3865, n3870, n3875, n3880,
    n3885, n3890, n3895, n3900, n3905, n3910, n3915, n3920, n3925, n3930,
    n3935, n3940, n3945, n3950, n3955, n3960, n3965, n3970, n3975, n3980,
    n3985, n3990, n3995, n4000, n4005, n4009, n4014, n4019, n4024, n4029,
    n4034, n4039, n4044, n4049, n4054, n4059, n4064, n4069, n4074, n4079,
    n4084, n4089, n4094, n4099, n4104, n4109, n4114, n4119, n4124, n4129,
    n4134, n4139, n4144, n4149, n4154, n4159, n4164, n4169, n4174, n4179,
    n4184, n4189, n4194, n4199, n4204, n4209, n4214, n4219, n4224, n4229,
    n4234, n4239, n4244, n4249, n4254, n4259, n4264, n4269, n4274, n4279,
    n4284, n4289, n4294, n4299, n4304, n4309, n4314, n4319, n4324, n4329,
    n4334, n4339, n4344, n4349, n4354, n4359, n4364, n4369, n4374, n4379,
    n4384, n4389, n4394, n4399, n4404, n4409, n4414, n4419, n4424, n4429,
    n4434, n4439, n4444, n4449, n4454, n4459, n4464, n4469, n4474, n4479,
    n4484, n4489, n4494, n4499, n4504, n4509, n4514, n4519, n4524, n4529,
    n4534, n4539, n4544, n4549, n4554, n4559, n4564, n4569, n4574, n4579,
    n4584, n4589, n4594, n4599, n4604, n4609, n4614, n4619, n4624, n4629,
    n4634, n4639, n4644, n4649, n4654, n4659, n4664, n4669, n4674, n4679,
    n4684, n4689, n4694, n4699, n4704, n4709, n4714, n4719, n4724, n4729,
    n4734, n4739, n4744, n4749, n4754, n4759, n4764, n4769, n4774, n4779,
    n4784, n4789, n4794, n4799, n4804, n4809, n4814, n4819, n4824, n4829,
    n4834, n4839, n4844, n4849, n4854, n4859, n4864, n4869, n4874, n4879,
    n4884, n4889, n4894, n4899, n4904, n4909, n4914, n4919, n4924, n4929,
    n4934, n4939, n4944, n4949, n4954, n4959, n4964, n4969, n4974, n4979,
    n4984, n4989, n4994, n4999, n5004, n5009, n5014, n5019, n5024, n5029,
    n5034, n5039, n5044, n5049, n5054, n5059, n5064, n5069, n5074, n5079,
    n5084, n5089, n5094, n5099, n5104, n5109, n5114, n5119, n5124, n5129,
    n5134, n5139, n5144, n5149, n5154, n5159, n5164, n5169, n5174, n5179,
    n5184, n5189, n5194, n5199, n5204, n5209, n5214, n5219, n5224, n5229,
    n5234, n5239, n5244, n5249, n5254, n5259, n5264, n5269, n5274, n5279,
    n5284, n5289, n5294, n5299, n5304, n5309, n5314, n5319, n5324, n5329,
    n5334, n5339, n5344, n5349, n5354, n5359, n5364, n5369, n5374, n5379,
    n5384, n5389, n5394, n5399, n5404, n5409, n5414, n5419, n5424, n5429,
    n5434, n5439, n5444, n5449, n5454, n5459, n5464, n5469, n5474, n5479,
    n5484, n5489, n5494, n5499, n5504, n5509, n5514, n5519, n5524, n5529,
    n5534, n5539, n5544, n5549, n5554, n5559, n5564, n5569, n5574, n5579,
    n5584, n5589, n5594, n5599, n5604, n5609, n5614, n5619, n5624, n5629,
    n5634, n5639, n5644, n5649, n5654, n5659, n5664, n5669, n5674, n5679,
    n5684, n5689, n5694, n5699, n5704, n5709, n5714, n5719, n5724, n5729,
    n5734, n5739, n5744, n5749, n5754, n5759, n5764, n5769, n5774, n5779,
    n5784, n5789, n5794, n5799, n5804, n5809, n5814, n5819, n5824, n5829,
    n5834, n5839, n5844, n5849, n5854, n5859, n5864, n5869, n5874, n5879,
    n5884, n5889, n5894, n5899, n5904, n5909, n5914, n5919, n5924, n5929,
    n5934, n5939, n5944, n5949, n5954, n5959, n5964, n5969, n5974, n5979,
    n5984, n5989, n5994, n5999, n6004, n6009, n6014, n6019, n6024, n6029,
    n6034, n6039, n6044, n6049, n6054, n6059, n6064, n6069, n6074, n6079,
    n6084, n6089, n6094;
  assign psv39_8_8_ = n_n7154 ? n_n9366 : tin_psv39_8_8_;
  assign psv39_0_0_ = n_n6986 ? n_n9424 : tin_psv39_0_0_;
  assign psv13_5_5_ = n_n7561 ? n_n9004 : tin_psv13_5_5_;
  assign psv2_13_13_ = n_n8245 ? n_n9169 : tin_psv2_13_13_;
  assign psv2_8_8_ = n_n8121 ? n_n8303 : tin_psv2_8_8_;
  assign psv38_2_2_ = n_n7146 ? n_n6910 : tin_psv38_2_2_;
  assign psv33_5_5_ = n_n7050 ? n_n9148 : tin_psv33_5_5_;
  assign psv26_6_6_ = n_n7622 ? n_n6980 : tin_psv26_6_6_;
  assign psv2_9_9_ = n_n8918 ? n_n7522 : tin_psv2_9_9_;
  assign psv18_2_2_ = n_n7905 ? n_n8801 : tin_psv18_2_2_;
  assign psv39_9_9_ = n_n7717 ? n_n7332 : tin_psv39_9_9_;
  assign psv39_1_1_ = n_n8946 ? n_n8430 : tin_psv39_1_1_;
  assign psv13_6_6_ = n_n8568 ? n_n7179 : tin_psv13_6_6_;
  assign psv2_6_6_ = n_n7150 ? n_n7022 : tin_psv2_6_6_;
  assign psv38_3_3_ = n_n7491 ? n_n7203 : tin_psv38_3_3_;
  assign psv33_6_6_ = n_n8243 ? n_n7344 : tin_psv33_6_6_;
  assign psv26_13_13_ = n_n7381 ? n_n7500 : tin_psv26_13_13_;
  assign psv26_12_12_ = n_n7798 ? n_n8488 : tin_psv26_12_12_;
  assign psv26_7_7_ = n_n7362 ? n_n8702 : tin_psv26_7_7_;
  assign psv2_7_7_ = n_n8392 ? n_n8061 : tin_psv2_7_7_;
  assign psv18_3_3_ = n_n7079 ? n_n7498 : tin_psv18_3_3_;
  assign psv39_2_2_ = n_n7978 ? n_n7726 : tin_psv39_2_2_;
  assign psv33_12_12_ = n_n7493 ? n_n8369 : tin_psv33_12_12_;
  assign psv33_11_11_ = n_n8665 ? n_n7923 : tin_psv33_11_11_;
  assign psv33_10_10_ = n_n9123 ? n_n9483 : tin_psv33_10_10_;
  assign psv13_7_7_ = n_n9228 ? n_n7546 : tin_psv13_7_7_;
  assign psv2_10_10_ = n_n7244 ? n_n8681 : tin_psv2_10_10_;
  assign psv38_4_4_ = n_n7052 ? n_n7674 : tin_psv38_4_4_;
  assign psv39_10_10_ = n_n7330 ? n_n8644 : tin_psv39_10_10_;
  assign psv33_7_7_ = n_n7140 ? n_n7843 : tin_psv33_7_7_;
  assign psv26_15_15_ = n_n8389 ? n_n9026 : tin_psv26_15_15_;
  assign psv26_14_14_ = n_n9200 ? n_n7392 : tin_psv26_14_14_;
  assign psv26_8_8_ = n_n6937 ? n_n7581 : tin_psv26_8_8_;
  assign psv26_0_0_ = n_n7246 ? n_n7017 : tin_psv26_0_0_;
  assign psv13_12_12_ = n_n8055 ? n_n8895 : tin_psv13_12_12_;
  assign psv13_11_11_ = n_n7336 ? n_n9548 : tin_psv13_11_11_;
  assign psv18_4_4_ = n_n9006 ? n_n9432 : tin_psv18_4_4_;
  assign psv39_3_3_ = n_n7507 ? n_n7108 : tin_psv39_3_3_;
  assign psv13_8_8_ = n_n7261 ? n_n7271 : tin_psv13_8_8_;
  assign psv13_0_0_ = n_n7176 ? n_n7775 : tin_psv13_0_0_;
  assign psv38_5_5_ = n_n8655 ? n_n7256 : tin_psv38_5_5_;
  assign psv33_8_8_ = n_n9306 ? n_n7288 : tin_psv33_8_8_;
  assign psv33_0_0_ = n_n8672 ? n_n8486 : tin_psv33_0_0_;
  assign psv26_9_9_ = n_n7310 ? n_n7360 : tin_psv26_9_9_;
  assign psv26_1_1_ = n_n7699 ? n_n7231 : tin_psv26_1_1_;
  assign psv13_10_10_ = n_n6956 ? n_n7976 : tin_psv13_10_10_;
  assign psv18_5_5_ = n_n7903 ? n_n7715 : tin_psv18_5_5_;
  assign psv39_4_4_ = n_n7117 ? n_n7121 : tin_psv39_4_4_;
  assign psv13_9_9_ = n_n7944 ? n_n9376 : tin_psv13_9_9_;
  assign psv13_1_1_ = n_n7013 ? n_n8589 : tin_psv13_1_1_;
  assign psv2_15_15_ = n_n6948 ? n_n8102 : tin_psv2_15_15_;
  assign psv2_11_11_ = n_n6952 ? n_n6963 : tin_psv2_11_11_;
  assign psv2_0_0_ = n_n7024 ? n_n8371 : tin_psv2_0_0_;
  assign psv38_14_14_ = n_n8454 ? n_n7174 : tin_psv38_14_14_;
  assign psv38_12_12_ = n_n8605 ? n_n7402 : tin_psv38_12_12_;
  assign psv38_10_10_ = n_n7181 ? n_n7284 : tin_psv38_10_10_;
  assign psv38_6_6_ = n_n7556 ? n_n7514 : tin_psv38_6_6_;
  assign psv18_15_15_ = n_n7019 ? n_n7074 : tin_psv18_15_15_;
  assign psv18_13_13_ = n_n7415 ? n_n7148 : tin_psv18_13_13_;
  assign psv18_11_11_ = n_n8195 ? n_n8439 : tin_psv18_11_11_;
  assign psv33_9_9_ = n_n8725 ? n_n9278 : tin_psv33_9_9_;
  assign psv33_1_1_ = n_n7635 ? n_n8091 : tin_psv33_1_1_;
  assign psv26_2_2_ = n_n7276 ? n_n7777 : tin_psv26_2_2_;
  assign psv2_1_1_ = n_n7467 ? n_n7678 : tin_psv2_1_1_;
  assign psv38_15_15_ = n_n8216 ? n_n8340 : tin_psv38_15_15_;
  assign psv38_11_11_ = n_n7033 ? n_n7857 : tin_psv38_11_11_;
  assign psv18_12_12_ = n_n8817 ? n_n9465 : tin_psv18_12_12_;
  assign psv18_6_6_ = n_n8230 ? n_n7156 : tin_psv18_6_6_;
  assign psv39_5_5_ = n_n8633 ? n_n8777 : tin_psv39_5_5_;
  assign psv13_2_2_ = n_n8251 ? n_n7130 : tin_psv13_2_2_;
  assign psv38_7_7_ = n_n8713 ? n_n8592 : tin_psv38_7_7_;
  assign psv39_12_12_ = n_n9476 ? n_n8100 : tin_psv39_12_12_;
  assign psv39_11_11_ = n_n7315 ? n_n7390 : tin_psv39_11_11_;
  assign psv33_2_2_ = n_n7209 ? n_n7111 : tin_psv33_2_2_;
  assign psv26_3_3_ = n_n7338 ? n_n8384 : tin_psv26_3_3_;
  assign psv13_14_14_ = n_n7959 ? n_n7252 : tin_psv13_14_14_;
  assign psv13_13_13_ = n_n8704 ? n_n6991 : tin_psv13_13_13_;
  assign psv18_10_10_ = n_n8974 ? n_n8146 : tin_psv18_10_10_;
  assign psv18_7_7_ = n_n7659 ? n_n8049 : tin_psv18_7_7_;
  assign psv39_6_6_ = n_n8047 ? n_n8073 : tin_psv39_6_6_;
  assign psv33_15_15_ = n_n7026 ? n_n8263 : tin_psv33_15_15_;
  assign psv33_14_14_ = n_n6988 ? n_n9429 : tin_psv33_14_14_;
  assign psv33_13_13_ = n_n8290 ? n_n7069 : tin_psv33_13_13_;
  assign psv13_3_3_ = n_n7586 ? n_n8850 : tin_psv13_3_3_;
  assign psv2_14_14_ = n_n8683 ? n_n7102 : tin_psv2_14_14_;
  assign psv2_12_12_ = n_n7286 ? n_n8132 : tin_psv2_12_12_;
  assign psv2_4_4_ = n_n7291 ? n_n8045 : tin_psv2_4_4_;
  assign psv38_8_8_ = n_n6984 ? n_n9421 : tin_psv38_8_8_;
  assign psv38_0_0_ = n_n8921 ? n_n8916 : tin_psv38_0_0_;
  assign psv39_14_14_ = n_n8441 ? n_n9371 : tin_psv39_14_14_;
  assign psv39_13_13_ = n_n8831 ? n_n7366 : tin_psv39_13_13_;
  assign psv33_3_3_ = n_n7409 ? n_n7420 : tin_psv33_3_3_;
  assign psv26_11_11_ = n_n7308 ? n_n8185 : tin_psv26_11_11_;
  assign psv26_10_10_ = n_n9580 ? n_n8781 : tin_psv26_10_10_;
  assign psv26_4_4_ = n_n8112 ? n_n8175 : tin_psv26_4_4_;
  assign psv13_15_15_ = n_n8406 ? n_n9145 : tin_psv13_15_15_;
  assign psv2_5_5_ = n_n9446 ? n_n7395 : tin_psv2_5_5_;
  assign psv18_8_8_ = n_n7242 ? n_n8678 : tin_psv18_8_8_;
  assign psv18_0_0_ = n_n7065 ? n_n7190 : tin_psv18_0_0_;
  assign psv39_7_7_ = n_n7183 ? n_n7160 : tin_psv39_7_7_;
  assign psv13_4_4_ = n_n9085 ? n_n9096 : tin_psv13_4_4_;
  assign psv2_2_2_ = n_n8510 ? n_n7054 : tin_psv2_2_2_;
  assign psv38_9_9_ = n_n8944 ? n_n8428 : tin_psv38_9_9_;
  assign psv38_1_1_ = n_n9373 ? n_n7964 : tin_psv38_1_1_;
  assign psv39_15_15_ = n_n7411 ? n_n8361 : tin_psv39_15_15_;
  assign psv33_4_4_ = n_n7003 ? n_n7462 : tin_psv33_4_4_;
  assign psv26_5_5_ = n_n8423 ? n_n7076 : tin_psv26_5_5_;
  assign psv2_3_3_ = n_n6912 ? n_n8750 : tin_psv2_3_3_;
  assign psv38_13_13_ = n_n9531 ? n_n6920 : tin_psv38_13_13_;
  assign psv18_14_14_ = n_n8762 ? n_n7435 : tin_psv18_14_14_;
  assign psv18_9_9_ = n_n6950 ? n_n6961 : tin_psv18_9_9_;
  assign psv18_1_1_ = n_n7387 ? n_n9535 : tin_psv18_1_1_;
  assign n491 = ~n4956 & ~preset & n_n9280;
  assign n496 = n6728 | (n_n9434 & n4845 & n4967);
  assign n501 = n6727 | (n_n9537 & n4845 & n4967);
  assign n506 = n6725 | n6726;
  assign n511 = ~n4956 & ~preset & n_n8270;
  assign n516 = ~n4956 & ~preset & n_n8196;
  assign n521 = ~n4956 & ~preset & n_n9150;
  assign n526 = n6479 | n6480;
  assign n531 = n6356 | (n1270 & n4848);
  assign n536 = n6354 | n6355;
  assign n541 = n6320 | n6321;
  assign n546 = n6319 | (ndn3_11 & ~ndn3_12 & n4850);
  assign n551 = ~preset & (n4851 ? n4930 : n_n7341);
  assign n556 = ~preset & (n4852 ? n4868 : n_n9180);
  assign n561 = n6317 | n6318;
  assign n566 = n6316 | (nen3_39 & ~ndn3_39 & n4855);
  assign n571 = n6314 | n6315;
  assign n576 = n6312 | n6313;
  assign n581 = n6310 | n6311;
  assign n586 = n6197 | (n4858 & n7122) | (~n4858 & n7121);
  assign n591 = n6196 | (n_n8354 & n4845 & n4967);
  assign n596 = ~preset & (n4859_1 ? n4903 : n_n7552);
  assign n601 = ~preset & ~nsr3_23;
  assign n606 = n6194 | n6195;
  assign n611 = n6192 | n6193;
  assign n616 = n6190 | n6191;
  assign n621 = ~preset & (n_n6950 | (ndn3_42 & ~ndn3_44));
  assign n626 = ~n4862 & (n_n8930 | (n4967 & n7089));
  assign n631 = ~preset & (n_n7244 | (~ndn3_42 & ndn3_40));
  assign n636 = n6189 | (n_n9512 & n4864_1 & n4967);
  assign n641 = ~preset & (n4865 ? n4868 : n_n8883);
  assign n646 = n6187 | n6188;
  assign n651 = ~preset & (n_n9580 | (nen3_22 & ~ndn3_22));
  assign n656 = n6186 | (n_n9353 & n4867 & n4967);
  assign n661 = n6185 | (n4863 & n4868);
  assign n666 = n6184 | (n4853 & (n4969_1 ^ n4970));
  assign n671 = n6182 | n6183;
  assign n676 = ~preset & (n4869_1 ? n4903 : n_n7373);
  assign n681 = ~preset & (n_n9085 | (~ngfdn_3 & ndn3_46));
  assign n686 = n6178 | n6179 | n6180 | n6181;
  assign n691 = n6177 | (~ndn3_29 & ndn3_28 & n4873);
  assign n696 = n6145 | n6146;
  assign n701 = ~preset & (n4875 ? n4930 : n_n7654);
  assign n706 = ~preset & (n4876 ? n4887 : n_n8410);
  assign n711 = n6082 | (ndn3_17 & ~ndn3_18 & n4878);
  assign n716 = n6081 | (~ndn3_7 & ndn3_4 & n4873);
  assign n721 = n6079_1 | n6080;
  assign n726 = n6078 | (n_n9512 & n4845 & n4967);
  assign n731 = n6077 | (~ndn3_19 & nen3_19 & n4855);
  assign n736 = ~preset & (n4865 ? n4848 : n_n8202);
  assign n741 = ~preset & (n4880 ? n4930 : n_n7670);
  assign n746 = n6075 | n6076;
  assign n751 = n6073 | n6074_1;
  assign n756 = n6071 | n6072;
  assign n761 = n6069_1 | n6070;
  assign n766 = n6068 | (n_n8449 & n4883 & n4967);
  assign n771 = n6067 | (n_n8419 & n4883 & n4967);
  assign n776 = n6065 | n6066;
  assign n781 = ~preset & (n4849_1 ? n4903 : n_n9141);
  assign n786 = n6063 | n6064_1;
  assign n791 = n6061 | n6062;
  assign n796 = n6059_1 | n6060;
  assign n801 = n6058 | (ndn3_11 & ~ndn3_12 & n4873);
  assign n806 = n6056 | n6057;
  assign n811 = n6054_1 | n6055;
  assign n816 = n6052 | n6053;
  assign n821 = ~preset & (n4854_1 ? n4903 : n_n7376);
  assign n826 = n6051 | (ndn3_9 & ~ndn3_11 & n4878);
  assign n831 = (n4005 & n4884_1) | (~preset & pover_0_0_ & ~n4884_1);
  assign n835 = ~preset & (n4877 ? n4887 : n_n8599);
  assign n840 = n6050 | (ndn3_11 & ~ndn3_12 & n4855);
  assign n845 = ~n4956 & ~preset & n_n9442;
  assign n850 = ~preset & (n4860 ? n4868 : n_n9485);
  assign n855 = n6048 | n6049_1;
  assign n860 = n6047 | (n_n9284 & n4864_1 & n4967);
  assign n865 = n6046 | (ndn3_19 & ~ndn3_21 & n4873);
  assign n870 = ~preset & ~ngfdn_3 & (ndn3_9 | ndn3_7);
  assign n875 = ~n4956 & ~preset & n_n8613;
  assign n880 = n6045 | (n_n8707 & n4867 & n4967);
  assign n885 = n6044_1 | (n_n9512 & n4886 & n4967);
  assign n890 = n6042 | n6043;
  assign n895 = n6041 | (n4853 & n4887);
  assign n900 = ~preset & (n_n8655 | (~ndn3_46 & ndn3_44));
  assign n905 = n6040 | (~ndn3_29 & ndn3_28 & n4888);
  assign n910 = ~n4956 & ~preset & n_n7583;
  assign n915 = n7174 | (n_n9248 & (~n_n9247 | ~n4902));
  assign n920 = n6038 | n6039_1;
  assign n925 = n6037 | (~ndn3_7 & ndn3_4 & n4888);
  assign n930 = n6035 | n6036;
  assign n935 = ~preset & (n4889_1 ? n4903 : n_n7738);
  assign n940 = ~n4956 & ~preset & n_n8573;
  assign n945 = ~preset & (n4880 ? n4868 : n_n9473);
  assign n950 = n6034_1 | (~ndn3_25 & ndn3_22 & n4873);
  assign n955 = n6033 | (n_n8557 & n4890 & n4967);
  assign n960 = ~n4956 & ~preset & n_n9554;
  assign n965 = ~n4956 & ~preset & n_n8508;
  assign n970 = n6031 | n6032;
  assign n975 = n6029_1 | n6030;
  assign n980 = n6027 | n6028;
  assign n985 = n6025 | n6026;
  assign n990 = ~preset & (n_n7409 | (ngfdn_3 & ~ndn3_50));
  assign n995 = ~n4956 & ~preset & n_n9437;
  assign n1000 = n6023 | n6024_1;
  assign n1005 = ~n4956 & ~preset & n_n8647;
  assign n1010 = n6021 | n6022;
  assign n1015 = n6019_1 | n6020;
  assign n1020 = ~preset & ~nsr3_13;
  assign n1025 = ~preset & ~ngfdn_3 & (ndn3_17 | ndn3_16);
  assign n1030 = ~preset & ~ngfdn_3 & (ndn3_25 | ndn3_22);
  assign n1035 = ~preset & ~ngfdn_3 & (ndn3_29 | ndn3_28);
  assign n1040 = ~n4956 & ~preset & n_n9539;
  assign n1045 = n6018 | (n_n8821 & n4883 & n4967);
  assign n1050 = n6016 | n6017;
  assign n1055 = ~preset & ~ngfdn_3 & (nen3_22 | ~nsr3_23);
  assign n1060 = ~n4956 & ~preset & n_n9438;
  assign n1065 = n6014_1 | n6015;
  assign n1070 = n6013 | (n_n9416 & n4891 & n4967);
  assign n1075 = n6011 | n6012;
  assign n1080 = n6009_1 | n6010;
  assign n1085 = n6008 | (n_n9353 & n4886 & n4967);
  assign n1090 = ~preset & (n_n7798 | (nen3_22 & ~ndn3_22));
  assign n1095 = n6004_1 | n6005 | n6006 | n6007;
  assign n1100 = ~preset & (n4859_1 ? n4904_1 : n_n7910);
  assign n1105 = ~preset & (n4881 ? n4903 : n_n9528);
  assign n1110 = n6002 | n6003;
  assign n1115 = ~preset & (n_n8251 | (~ngfdn_3 & ndn3_46));
  assign n1120 = n6000 | n6001;
  assign n1125 = n5998 | n5999_1;
  assign n1130 = ~n4956 & ~preset & n_n9290;
  assign n1135 = n5996 | n5997;
  assign n1140 = ~preset & (n_n7556 | (~ndn3_46 & ndn3_44));
  assign n1145 = n5995 | (n_n8449 & n4886 & n4967);
  assign n1150 = n5993 | n5994_1;
  assign n1155 = n5992 | (ndn3_19 & ~ndn3_21 & n4855);
  assign n1160 = ~n4956 & ~preset & n_n9361;
  assign n1165 = ~preset & (n4885 ? n4848 : n_n9304);
  assign n1170 = n5991 | (n_n8652 & n4896 & n4967);
  assign n1175 = ~preset & (n4877 ? n4848 : n_n7712);
  assign n1180 = n5990 | (n_n8707 & n4896 & n4967);
  assign n1185 = n5989_1 | (n_n8549 & n4883 & n4967);
  assign n1190 = n5988 | (~nsr3_13 & ~ndn3_15 & n4855);
  assign n1195 = n5986 | n5987;
  assign n1200 = ~preset & (n4849_1 ? n4930 : n_n9015);
  assign n1205 = n5985 | (n_n8354 & n4891 & n4967);
  assign n1210 = ~preset & (n4880 ? n4887 : n_n9518);
  assign n1215 = n5983 | n5984_1;
  assign n1220 = n5982 | (n_n9448 & n4883 & n4967);
  assign n1225 = n5980 | n5981;
  assign n1230 = n5978 | n5979_1;
  assign n1235 = n5976 | n5977;
  assign n1240 = ~preset & (n4849_1 ? n4887 : n_n7951);
  assign n1245 = n5974_1 | n5973 | (n_n8913 & n4898);
  assign n1250 = ~preset & (n4877 ? n4903 : n_n8035);
  assign n1255 = n5972 | n5971 | (n_n8631 & n4898);
  assign n1260 = ~preset & (n_n8243 | (ngfdn_3 & ~ndn3_50));
  assign n1265 = n5969_1 | n5970;
  assign n1270 = ndn3_46 & ~preset & ~ngfdn_3;
  assign n1275 = n5968 | (ndn3_9 & ~ndn3_11 & n4855);
  assign n1280 = ~preset & (n4859_1 ? n4868 : n_n9175);
  assign n1285 = n5966 | n5967;
  assign n1290 = n5965 | (n_n9284 & n4891 & n4967);
  assign n1295 = n5963 | n5964_1;
  assign n1300 = ~n4956 & ~preset & n_n9410;
  assign n1305 = n5962 | (n4861 & n4887);
  assign n1310 = n5961 | (n_n8707 & n4886 & n4967);
  assign n1315 = n5960 | (n_n9512 & n4867 & n4967);
  assign n1320 = n5958 | n5959_1;
  assign n1325 = n5957 | (n4863 & n4887);
  assign n1330 = n5955 | n5956;
  assign n1335 = n5954_1 | (~nsr3_13 & ~ndn3_15 & n4888);
  assign n1340 = n5953 | (nen3_16 & ~ndn3_16 & n4850);
  assign n1345 = n5952 | preset | pdn;
  assign n1350 = n5951 | (n_n9353 & n4845 & n4967);
  assign n1355 = ~n4956 & ~preset & n_n8531;
  assign n1360 = n5950 | (n_n9638 & n4845 & n4967);
  assign n1365 = n5949_1 | (n1270 & (n4985 ^ n4986));
  assign n1370 = n5948 | (nen3_39 & ~ndn3_39 & n4878);
  assign n1375 = ~preset & (n_n8112 | (nen3_22 & ~ndn3_22));
  assign n1380 = n5946 | n5947;
  assign n1385 = ~preset & (n4889_1 ? n4887 : n_n9618);
  assign n1390 = n5944_1 | n5945;
  assign n1395 = ~n4956 & ~preset & n_n9242;
  assign n1400 = n5943 | (n4848 & n4853);
  assign n1405 = ~preset & (n4882 ? n4868 : n_n8884);
  assign n1410 = n5941 | n5942;
  assign n1415 = n5940 | (n_n8549 & n4845 & n4967);
  assign n1420 = n5939_1 | (n4853 & (n4976 ^ n4977));
  assign n1425 = ~preset & (n4876 ? n4904_1 : n_n7909);
  assign n1430 = n5938 | (n4861 & (n4976 ^ n4977));
  assign n1435 = n5937 | (~ndn3_4 & ndn3_2 & n4850);
  assign n1440 = ~preset & (n4860 ? n4930 : n_n8862);
  assign n1445 = ~n4956 & ~preset & n_n8037;
  assign n1450 = ~preset & ~ngfdn_3 & (ndn3_17 | ndn3_18);
  assign n1455 = ~preset & ~ngfdn_3 & (nen3_22 | ndn3_22);
  assign n1460 = ~preset & (n_n8974 | (ndn3_42 & ~ndn3_44));
  assign n1465 = ~preset & (n_n7286 | (~ndn3_42 & ndn3_40));
  assign n1470 = n5935 | n5936;
  assign n1475 = ~preset & n4902;
  assign n1480 = n5933 | n5934_1;
  assign n1485 = n5931 | n5932;
  assign n1490 = ~preset & ~ngfdn_3 & (nen3_39 | ~nsr3_38);
  assign n1495 = n5929_1 | n5930;
  assign n1500 = ~n4956 & ~preset & n_n9557;
  assign n1505 = n5928 | (n_n8354 & n4896 & n4967);
  assign n1510 = n5926 | n5927;
  assign n1515 = n5924_1 | n5925;
  assign n1520 = n5923 | (n_n9537 & n4886 & n4967);
  assign n1525 = ~preset & (n_n8568 | (~ngfdn_3 & ndn3_46));
  assign n1530 = n5921 | n5922;
  assign n1535 = ~preset & (n4889_1 ? n4904_1 : n_n7931);
  assign n1540 = ~preset & (n4879_1 ? n4903 : n_n7742);
  assign n1545 = n5920 | (ndn3_19 & ~ndn3_21 & n4878);
  assign n1550 = n5919_1 | (n_n8549 & n4886 & n4967);
  assign n1555 = ~preset & (n4874_1 ? n4904_1 : n_n9568);
  assign n1560 = ~preset & (n_n9200 | (nen3_22 & ~ndn3_22));
  assign n1565 = n5917 | n5918;
  assign n1570 = n5915 | n5916;
  assign n1575 = n5914_1 | (nen3_16 & ~ndn3_16 & n4878);
  assign n1580 = n5912 | n5913;
  assign n1585 = n5910 | n5911;
  assign n1590 = ~preset & (n4880 ? n4903 : n_n8499);
  assign n1595 = n5908 | n5909_1;
  assign n1600 = n5906 | n5907;
  assign n1605 = n5905 | (ndn3_29 & ~ndn3_32 & n4873);
  assign n1610 = n5903 | n5904_1;
  assign n1615 = n5901 | n5902;
  assign n1620 = ~preset & (n4852 ? n4848 : n_n7713);
  assign n1625 = ~preset & (n4852 ? n4930 : n_n9566);
  assign n1630 = n5899_1 | n5900;
  assign n1635 = n5897 | n5898;
  assign n1640 = n5896 | (~ndn3_7 & ndn3_4 & n4878);
  assign n1645 = ~n4956 & ~preset & n_n9560;
  assign n1650 = n5894_1 | n5895;
  assign n1655 = n5892 | n5893;
  assign n1660 = ~preset & (n4851 ? n4868 : n_n8882);
  assign n1665 = n5890 | n5891;
  assign n1670 = n5888 | n5889_1;
  assign n1675 = n5887 | (ndn3_25 & ~ndn3_26 & n4888);
  assign n1680 = n5885 | n5886;
  assign n1685 = n5883 | n5884_1;
  assign n1690 = n5882 | (n_n9537 & n4883 & n4967);
  assign n1695 = ~n4956 & ~preset & n_n8875;
  assign n1700 = n5880 | n5881;
  assign n1705 = n5878 | n5879_1;
  assign n1710 = n5877 | (n4846 & n4887);
  assign n1715 = n5876 | (n4863 & n4903);
  assign n1720 = n5875 | (n4853 & (n4971 ^ n4972));
  assign n1725 = n5874_1 | (n_n9416 & n4867 & n4967);
  assign n1730 = n5873 | (n_n8821 & n4886 & n4967);
  assign n1735 = n5871 | n5872;
  assign n1740 = ~n4956 & ~preset & n_n7702;
  assign n1745 = n7177 | (nsr3_23 & ~ndn3_19);
  assign n1750 = ~n4956 & ~preset & n_n8199;
  assign n1755 = ~n4956 & ~preset & n_n7983;
  assign n1760 = n5870 | (n1270 & n4904_1);
  assign n1765 = n5868 | n5869_1;
  assign n1770 = n5867 | (n_n9434 & n4896 & n4967);
  assign n1775 = ~n4956 & ~preset & n_n8348;
  assign n1780 = n5865 | n5866;
  assign n1785 = n5864_1 | (n_n8549 & n4890 & n4967);
  assign n1790 = n5862 | n5863;
  assign n1795 = n5861 | (n_n9638 & n4896 & n4967);
  assign n1800 = n5860 | (n4848 & n4863);
  assign n1805 = n5858 | n5859_1;
  assign n1810 = n5856 | n5857;
  assign n1815 = n5854_1 | n5855;
  assign n1820 = n5853 | (n4863 & (n4976 ^ n4977));
  assign n1825 = n5852 | (n_n8419 & n4890 & n4967);
  assign n1830 = n5851 | (n4846 & (n4976 ^ n4977));
  assign n1835 = n5850 | (n_n8354 & n4890 & n4967);
  assign n1840 = n5849_1 | (n_n8652 & n4883 & n4967);
  assign n1845 = n5848 | (ndn3_17 & ~ndn3_18 & n4888);
  assign n1850 = n5847 | (n_n8707 & n4883 & n4967);
  assign n1855 = n5845 | n5846;
  assign n1860 = ~preset & ~nsr3_30;
  assign n1865 = n5843 | n5844_1;
  assign n1870 = ~preset & (n4859_1 ? n4887 : n_n7693);
  assign n1875 = ~preset & ~ngfdn_3 & (nen3_16 | ~nsr3_14);
  assign n1880 = n5841 | n5842;
  assign n1885 = n5840 | (~ndn3_29 & ndn3_28 & n4878);
  assign n1890 = n5839_1 | (n_n9512 & n4891 & n4967);
  assign n1895 = n5837 | n5838;
  assign n1900 = n5836 | (n_n8821 & n4891 & n4967);
  assign n1905 = ~preset & (n4880 ? n4848 : n_n9110);
  assign n1910 = n5834_1 | n5835;
  assign n1915 = n5833 | (n4853 & n4868);
  assign n1920 = n5832 | (n4863 & (n4969_1 ^ n4970));
  assign n1925 = n5830 | n5831;
  assign n1930 = n5828 | n5829_1;
  assign n1935 = n5827 | (~ndn3_27 & ndn3_26 & n4855);
  assign n1940 = ~preset & (n_n8406 | (~ngfdn_3 & ndn3_46));
  assign n1945 = n5826 | (~ndn3_19 & nen3_19 & n4878);
  assign n1950 = n5825 | (n_n8549 & n4867 & n4967);
  assign n1955 = ~preset & (n4869_1 ? n4887 : n_n7474);
  assign n1960 = n5824_1 | (n1270 & (n4954_1 ^ n4955));
  assign n1965 = ~preset & (n_n6984 | (~ndn3_46 & ndn3_44));
  assign n1970 = n5823 | (n4848 & n4866);
  assign n1975 = n5821 | n5822;
  assign n1980 = ~n4956 & ~preset & n_n9559;
  assign n1985 = ~preset & (n_n7362 | (nen3_22 & ~ndn3_22));
  assign n1990 = n5819_1 | n5820;
  assign n1995 = ~n4956 & ~preset & n_n9550;
  assign n2000 = ~preset & (n4889_1 ? n4868 : n_n9492);
  assign n2005 = n5817 | n5818;
  assign n2010 = ~preset & (n4879_1 ? n4848 : n_n7764);
  assign n2015 = n5815 | n5816;
  assign n2020 = n5813 | n5814_1;
  assign n2025 = n5811 | n5812;
  assign n2030 = ~n4956 & ~preset & n_n8173;
  assign n2035 = n5809_1 | n5810;
  assign n2040 = n5807 | n5808;
  assign n2045 = ~preset & (n4882 ? n4887 : n_n8753);
  assign n2050 = ~preset & (n4852 ? n4904_1 : n_n8772);
  assign n2055 = n5805 | n5806;
  assign n2060 = ~n4956 & ~preset & n_n9362;
  assign n2065 = ndn1_4 & ~preset & ~pdn;
  assign n2070 = ~n4956 & ~preset & n_n9561;
  assign n2075 = n5803 | n5804_1;
  assign n2080 = ~preset & (n4849_1 ? n4848 : n_n8203);
  assign n2085 = n5801 | n5802;
  assign n2090 = n5799_1 | n5800;
  assign n2095 = n5797 | n5798;
  assign n2100 = ~n4956 & ~preset & n_n9331;
  assign n2105 = n5796 | (~ndn3_19 & nen3_19 & n4873);
  assign n2110 = ~preset & ~ngfdn_3 & (ndn3_7 | ndn3_4);
  assign n2115 = n5795 | (n4853 & n4903);
  assign n2120 = n5794_1 | (n4863 & (n4971 ^ n4972));
  assign n2125 = n5793 | (n_n9416 & n4886 & n4967);
  assign n2130 = n5792 | (n_n8821 & n4867 & n4967);
  assign n2135 = ~preset & (n4881 ? n4868 : n_n9497);
  assign n2140 = ~preset & (n_n7291 | (~ndn3_42 & ndn3_40));
  assign n2145 = n7178 | (nsr3_13 & ~ndn3_12);
  assign n2150 = n7179 | (nsr3_38 & ~nen3_36);
  assign n2155 = ~n4956 & ~preset & n_n8240;
  assign n2160 = ~n4956 & ~preset & n_n7703;
  assign n2165 = n5791 | (n1270 & n4887);
  assign n2170 = ~n4956 & ~preset & n_n8237;
  assign n2175 = ~n4956 & ~preset & n_n8935;
  assign n2180 = ~n4956 & ~preset & n_n9244;
  assign n2185 = ~n4956 & ~preset & n_n8648;
  assign n2190 = ~n4956 & ~preset & n_n8235;
  assign n2195 = ~preset & (n4854_1 ? n4904_1 : n_n8611);
  assign n2200 = n5789_1 | n5790;
  assign n2205 = n5788 | (ndn3_29 & ~ndn3_32 & n4888);
  assign n2210 = ~n4956 & ~preset & n_n8572;
  assign n2215 = n5786 | n5787;
  assign n2220 = n5785 | (~ndn3_9 & ndn3_7 & n4850);
  assign n2225 = ~n4956 & ~preset & n_n9555;
  assign n2230 = n5783 | n5784_1;
  assign n2235 = ~preset & (n_n7050 | (ngfdn_3 & ~ndn3_50));
  assign n2240 = n5782 | (~ndn3_9 & ndn3_7 & n4888);
  assign n2245 = ~preset & (n_n7140 | (ngfdn_3 & ~ndn3_50));
  assign n2250 = n5781 | (n_n9448 & n4890 & n4967);
  assign n2255 = ~preset & (n_n6948 | (~ndn3_42 & ndn3_40));
  assign n2260 = n5777 | n5778 | n5779_1 | n5780;
  assign n2265 = ~preset & ~ngfdn_3 & (ndn3_19 | nen3_19);
  assign n2270 = ~preset & ~ngfdn_3 & (ndn3_28 | nen3_28);
  assign n2275 = n5775 | n5776;
  assign n2280 = n5773 | n5774_1;
  assign n2285 = n5772 | (n4861 & (n4954_1 ^ n4955));
  assign n2290 = n5771 | (n_n8707 & n4891 & n4967);
  assign n2295 = n5770 | (~ndn3_19 & nen3_19 & n4850);
  assign n2300 = ~preset & ~ngfdn_3 & (nen3_36 | ~nsr3_37);
  assign n2305 = n5769_1 | (n_n9284 & n4867 & n4967);
  assign n2310 = n5767 | n5768;
  assign n2315 = ~preset & (n4892 ? n4903 : n_n7736);
  assign n2320 = n5765 | n5766;
  assign n2325 = n5763 | n5764_1;
  assign n2330 = ~preset & (n4892 ? n4887 : n_n8891);
  assign n2335 = n5761 | n5762;
  assign n2340 = n5760 | (n_n8557 & n4867 & n4967);
  assign n2345 = n5758 | n5759_1;
  assign n2350 = ~n4956 & ~preset & n_n9558;
  assign n2355 = n5757 | (n4866 & (n4954_1 ^ n4955));
  assign n2360 = n5756 | (~nsr3_13 & ~ndn3_15 & n4878);
  assign n2365 = ~preset & (n_n6956 | (~ngfdn_3 & ndn3_46));
  assign n2370 = ~preset & (n4847 ? n4903 : n_n8298);
  assign n2375 = n5755 | (~ndn3_25 & ndn3_22 & n4850);
  assign n2380 = n5753 | n5754_1;
  assign n2385 = n5751 | n5752;
  assign n2390 = ~n4956 & ~preset & n_n9552;
  assign n2395 = n5750 | n5749_1 | (n_n8964 & n4898);
  assign n2400 = ~n4956 & ~preset & n_n8016;
  assign n2405 = n5747 | n5748;
  assign n2410 = ~preset & (n4874_1 ? n4887 : n_n7696);
  assign n2415 = n5745 | n5746;
  assign n2420 = n5744_1 | (~ndn3_27 & ndn3_26 & n4888);
  assign n2425 = n5743 | (n_n9353 & n4891 & n4967);
  assign n2430 = n7181 | (~preset & n_n8652 & ~n5001);
  assign n2435 = n7184 | (~preset & n_n8707 & ~n5001);
  assign n2440 = n5741 | n5742;
  assign n2445 = n5739_1 | n5740;
  assign n2450 = n5738 | (~ndn3_29 & ndn3_28 & n4850);
  assign n2455 = n7185 | (nsr3_30 & ~nak3_13);
  assign n2460 = ~n4956 & ~preset & n_n8274;
  assign n2465 = ~n4956 & ~preset & n_n8615;
  assign n2470 = ~n4956 & ~preset & n_n8238;
  assign n2475 = ~n4956 & ~preset & n_n7854;
  assign n2480 = ~n4956 & ~preset & n_n8649;
  assign n2485 = ~n4956 & ~preset & n_n8236;
  assign n2490 = ~n4956 & ~preset & n_n8269;
  assign n2495 = n5737 | (n_n9537 & n4896 & n4967);
  assign n2500 = n5735 | n5736;
  assign n2505 = n5733 | n5734_1;
  assign n2510 = ~n4956 & ~preset & n_n8529;
  assign n2515 = n5732 | (nen3_36 & ~ndn3_36 & n4878);
  assign n2520 = n5731 | (n_n9434 & n4890 & n4967);
  assign n2525 = ~n4956 & ~preset & n_n8685;
  assign n2530 = ~preset & (n_n9531 | (~ndn3_46 & ndn3_44));
  assign n2535 = ~n4956 & ~preset & n_n9510;
  assign n2540 = ~n4956 & ~preset & n_n7771;
  assign n2545 = n5730 | (n_n8449 & n4845 & n4967);
  assign n2550 = n5728 | n5729_1;
  assign n2555 = n5727 | (nen3_36 & ~ndn3_36 & n4855);
  assign n2560 = ~preset & ~ngfdn_3 & (ndn3_9 | ndn3_11);
  assign n2565 = ~preset & ~ngfdn_3 & (~nsr3_13 | ndn3_15);
  assign n2570 = ~preset & ~ngfdn_3 & (ndn3_19 | ndn3_21);
  assign n2575 = ~n4956 & ~preset & n_n7584;
  assign n2580 = n5723 | n5724_1 | n5725 | n5726;
  assign n2585 = ~preset & (n_n6952 | (~ndn3_42 & ndn3_40));
  assign n2590 = n5722 | (ndn3_29 & ~ndn3_32 & n4878);
  assign n2595 = n5720 | n5721;
  assign n2600 = n5718 | n5719_1;
  assign n2605 = n5717 | (n_n8549 & n4896 & n4967);
  assign n2610 = n5716 | (n_n9284 & n4886 & n4967);
  assign n2615 = n5714_1 | n5715;
  assign n2620 = ~preset & (n_n7308 | (nen3_22 & ~ndn3_22));
  assign n2625 = n5712 | n5713;
  assign n2630 = n5711 | (n_n9537 & n4867 & n4967);
  assign n2635 = n5709_1 | n5710;
  assign n2640 = ~preset & (n_n6912 | (~ndn3_42 & ndn3_40));
  assign n2645 = n5707 | n5708;
  assign n2650 = n5706 | n5705 | (n_n8911 & n4898);
  assign n2655 = ~preset & (n4881 ? n4887 : n_n7952);
  assign n2660 = ~preset & (n_n8704 | (~ngfdn_3 & ndn3_46));
  assign n2665 = n5704_1 | (nen3_16 & ~ndn3_16 & n4873);
  assign n2670 = n5703 | (n4866 & (n4969_1 ^ n4970));
  assign n2675 = n5701 | n5702;
  assign n2680 = ~preset & (n4882 ? n4848 : n_n9019);
  assign n2685 = ~preset & (n_n7699 | (nen3_22 & ~ndn3_22));
  assign n2690 = ~preset & (n4882 ? n4903 : n_n7375);
  assign n2695 = n5699_1 | n5700;
  assign n2700 = n5697 | n5698;
  assign n2705 = n5696 | (ndn3_25 & ~ndn3_26 & n4850);
  assign n2710 = n5694_1 | n5695;
  assign n2715 = n5692 | n5693;
  assign n2720 = n5690 | n5691;
  assign n2725 = n5689_1 | (~ndn3_34 & nen3_34 & n4888);
  assign n2730 = ~n4956 & ~preset & n_n7582;
  assign n2735 = ~n4956 & ~preset & n_n8968;
  assign n2740 = n5687 | n5688;
  assign n2745 = n5685 | n5686;
  assign n2750 = n5683 | n5684_1;
  assign n2755 = ~preset & (n_n9373 | (~ndn3_46 & ndn3_44));
  assign n2760 = n4862 | (n_n9248 & (~n_n9247 | ~n4902));
  assign n2765 = n5682 | (n4866 & (n4971 ^ n4972));
  assign n2770 = n5680 | n5681;
  assign n2775 = ~n4956 & ~preset & n_n8273;
  assign n2780 = ~preset & (n_n6937 | (nen3_22 & ~ndn3_22));
  assign n2785 = n5679_1 | (nen3_16 & ~ndn3_16 & n4888);
  assign n2790 = n5677 | n5678;
  assign n2795 = n5676 | (n4846 & n4904_1);
  assign n2800 = n5675 | (n4863 & (n4985 ^ n4986));
  assign n2805 = n5673 | n5674_1;
  assign n2810 = n5671 | n5672;
  assign n2815 = n5670 | (n_n9284 & n4890 & n4967);
  assign n2820 = n5668 | n5669_1;
  assign n2825 = ~preset & (n_n7181 | (~ndn3_46 & ndn3_44));
  assign n2830 = n5666 | n5667;
  assign n2835 = n5664_1 | n5665;
  assign n2840 = n5662 | n5663;
  assign n2845 = n5661 | (~ndn3_17 & ndn3_16 & n4888);
  assign n2850 = ~preset & (n4851 ? n4903 : n_n7487);
  assign n2855 = n5659_1 | n5660;
  assign n2860 = n5657 | n5658;
  assign n2865 = n5656 | (n_n8449 & n4864_1 & n4967);
  assign n2870 = ~preset & (n4874_1 ? n4868 : n_n9181);
  assign n2875 = ~preset & (n_n8725 | (ngfdn_3 & ~ndn3_50));
  assign n2880 = n5654_1 | n5655;
  assign n2885 = ~preset & ~ngfdn_3 & (ndn3_27 | ndn3_26);
  assign n2890 = n5653 | (n_n8652 & n4891 & n4967);
  assign n2895 = ~preset & (n_n7415 | (ndn3_42 & ~ndn3_44));
  assign n2900 = n5652 | (n_n8557 & n4896 & n4967);
  assign n2905 = ~preset & ~ngfdn_3 & (nen3_19 | ~nsr3_20);
  assign n2910 = ~preset & (n_n8762 | (ndn3_42 & ~ndn3_44));
  assign n2915 = ~preset & (n4880 ? n4904_1 : n_n8512);
  assign n2920 = n5651 | (n_n8821 & n4864_1 & n4967);
  assign n2925 = n5650 | (~ndn3_19 & nen3_19 & n4888);
  assign n2930 = ~preset & (n_n7387 | (ndn3_42 & ~ndn3_44));
  assign n2935 = n5649_1 | (n_n9434 & n4886 & n4967);
  assign n2940 = n5647 | n5648;
  assign n2945 = n5645 | n5646;
  assign n2950 = ~preset & (n4892 ? n4848 : n_n9157);
  assign n2955 = n5644_1 | (nen3_36 & ~ndn3_36 & n4873);
  assign n2960 = ~preset & (n_n7381 | (nen3_22 & ~ndn3_22));
  assign n2965 = ~preset & (n_n9446 | (~ndn3_42 & ndn3_40));
  assign n2970 = ~preset & (n_n8633 | (ndn3_39 & ~ndn3_40));
  assign n2975 = n5643 | (n4866 & (n4976 ^ n4977));
  assign n2980 = ~preset & (n_n7310 | (nen3_22 & ~ndn3_22));
  assign n2985 = n5642 | (ndn3_17 & ~ndn3_18 & n4855);
  assign n2990 = n5640 | n5641;
  assign n2995 = n5639_1 | (n_n8821 & n4896 & n4967);
  assign n3000 = n5637 | n5638;
  assign n3005 = n5635 | n5636;
  assign n3010 = n5633 | n5634_1;
  assign n3015 = ~preset & (n_n7315 | (ndn3_39 & ~ndn3_40));
  assign n3020 = ~preset & (n_n9476 | (ndn3_39 & ~ndn3_40));
  assign n3025 = n5631 | n5632;
  assign n3030 = n5630 | (n_n9638 & n4883 & n4967);
  assign n3035 = n5628 | n5629_1;
  assign n3040 = n5627 | (~ndn3_28 & nen3_28 & n4850);
  assign n3045 = n7190 | (~n4894_1 & (n7188 | n7189));
  assign n3050 = n5624_1 | n5625;
  assign n3055 = n7191 | (~ndn3_29 & nsr3_35);
  assign n3060 = ~preset & (n_n7154 | (ndn3_39 & ~ndn3_40));
  assign n3065 = ~preset & (n4875 ? n4868 : n_n9495);
  assign n3070 = n5622 | n5623;
  assign n3075 = n5621 | (n4866 & n4887);
  assign n3080 = n5619_1 | n5620;
  assign n3085 = n5617 | n5618;
  assign n3090 = n5615 | n5616;
  assign n3095 = n5614_1 | (n4853 & (n4985 ^ n4986));
  assign n3100 = n5612 | n5613;
  assign n3105 = ~n4956 & ~preset & n_n8970;
  assign n3110 = n5610 | n5611;
  assign n3115 = n5608 | n5609_1;
  assign n3120 = ~preset & (n_n7246 | (nen3_22 & ~ndn3_22));
  assign n3125 = n5606 | n5607;
  assign n3130 = n5604_1 | n5605;
  assign n3135 = ~preset & (n_n7635 | (ngfdn_3 & ~ndn3_50));
  assign n3140 = n5603 | (ndn3_11 & ~ndn3_12 & n4888);
  assign n3145 = n5601 | n5602;
  assign n3150 = n5600 | (nen3_39 & ~ndn3_39 & n4850);
  assign n3155 = ~preset & (n4860 ? n4904_1 : n_n9108);
  assign n3160 = ~preset & (n4851 ? n4887 : n_n9286);
  assign n3165 = ~preset & ~ngfdn_3 & (ndn3_11 | ndn3_12);
  assign n3170 = ~preset & ~ngfdn_3 & (nen3_16 | ndn3_16);
  assign n3175 = ~preset & (n4876 ? n4848 : n_n7708);
  assign n3180 = n5599_1 | (n_n8419 & n4864_1 & n4967);
  assign n3185 = n5598 | (n_n8652 & n4864_1 & n4967);
  assign n3190 = ~preset & (n4860 ? n4887 : n_n7947);
  assign n3195 = n5596 | n5597;
  assign n3200 = n5595 | (n_n8707 & n4864_1 & n4967);
  assign n3205 = n5594_1 | (ndn3_19 & ~ndn3_21 & n4850);
  assign n3210 = ~preset & (n_n7659 | (ndn3_42 & ~ndn3_44));
  assign n3215 = ~n4956 & ~preset & n_n7630;
  assign n3220 = n5593 | (ndn3_19 & ~ndn3_21 & n4888);
  assign n3225 = ~n4956 & ~preset & n_n8691;
  assign n3230 = n5592 | (n_n9434 & n4867 & n4967);
  assign n3235 = n5591 | (~ndn3_28 & nen3_28 & n4873);
  assign n3240 = ~preset & (n4876 ? n4930 : n_n7995);
  assign n3245 = n5589_1 | n5590;
  assign n3250 = n5588 | (~nsr3_13 & ~ndn3_15 & n4873);
  assign n3255 = ~preset & (n_n7507 | (ndn3_39 & ~ndn3_40));
  assign n3260 = ~preset & (n_n7959 | (~ngfdn_3 & ndn3_46));
  assign n3265 = n5586 | n5587;
  assign n3270 = n5584_1 | n5585;
  assign n3275 = n5582 | n5583;
  assign n3280 = n5581 | (n_n9448 & n4886 & n4967);
  assign n3285 = ~preset & (n4881 ? n4904_1 : n_n8106);
  assign n3290 = n5579_1 | n5580;
  assign n3295 = n5577 | n5578;
  assign n3300 = n5575 | n5576;
  assign n3305 = n5574_1 | (~ndn3_9 & ndn3_7 & n4873);
  assign n3310 = n5573 | (~ndn3_9 & ndn3_7 & n4878);
  assign n3315 = n5571 | n5572;
  assign n3320 = ~preset & (n4885 ? n4930 : n_n9087);
  assign n3325 = n5569_1 | n5570;
  assign n3330 = ~n4956 & ~preset & n_n7852;
  assign n3335 = n5567 | n5568;
  assign n3340 = ~preset & (~n_n9198 | (~n4967 & n4974_1));
  assign n3345 = n5563 | n5564_1 | n5565 | n5566;
  assign n3350 = n7193 | preset | (nsr3_13 & nsr3_14);
  assign n3355 = n7197 | n5561 | n5562;
  assign n3360 = ~preset & (n_n7026 | (ngfdn_3 & ~ndn3_50));
  assign n3365 = n5559_1 | n5560;
  assign n3370 = ~n4956 & ~preset & n_n8272;
  assign n3375 = n5558 | (n_n9284 & n4896 & n4967);
  assign n3380 = ~n4956 & ~preset & n_n7985;
  assign n3385 = ~n4956 & ~preset & n_n8312;
  assign n3390 = n5556 | n5557;
  assign n3395 = n5554_1 | n5555;
  assign n3400 = n5552 | n5553;
  assign n3405 = ~preset & (n_n8683 | (~ndn3_42 & ndn3_40));
  assign n3410 = ~preset & ~ngfdn_3 & (nen3_39 | ndn3_39);
  assign n3415 = ~preset & (n_n8245 | (~ndn3_42 & ndn3_40));
  assign n3420 = n5551 | (~ndn3_34 & nen3_34 & n4873);
  assign n3425 = n5549_1 | n5550;
  assign n3430 = n5547 | n5548;
  assign n3435 = n5545 | n5546;
  assign n3440 = n5544_1 | (n_n8419 & n4896 & n4967);
  assign n3445 = n5543 | (n_n9638 & n4886 & n4967);
  assign n3450 = n5541 | n5542;
  assign n3455 = ~preset & (n4869_1 ? n4848 : n_n8201);
  assign n3460 = n5540 | (~ndn3_4 & ndn3_2 & n4855);
  assign n3465 = n5538 | n5539_1;
  assign n3470 = ~preset & (n_n8389 | (nen3_22 & ~ndn3_22));
  assign n3475 = ~n4956 & ~preset & n_n9440;
  assign n3480 = n5536 | n5537;
  assign n3485 = n5535 | (n_n8354 & n4886 & n4967);
  assign n3490 = n5534_1 | (n_n9448 & n4867 & n4967);
  assign n3495 = n5533 | (n_n9416 & n4896 & n4967);
  assign n3500 = n5531 | n5532;
  assign n3505 = n5530 | (~ndn3_7 & ndn3_4 & n4855);
  assign n3510 = n5529_1 | (n_n8354 & n4883 & n4967);
  assign n3515 = n5527 | n5528;
  assign n3520 = ~preset & (n_n7209 | (ngfdn_3 & ~ndn3_50));
  assign n3525 = ~preset & (n_n7003 | (ngfdn_3 & ~ndn3_50));
  assign n3530 = ~preset & (n4852 ? n4887 : n_n7695);
  assign n3535 = n5526 | (nen3_39 & ~ndn3_39 & n4873);
  assign n3540 = n5524_1 | n5525;
  assign n3545 = ~preset & (n4865 ? n4903 : n_n7374);
  assign n3550 = n5522 | n5523;
  assign n3555 = ~preset & (n_n7944 | (~ngfdn_3 & ndn3_46));
  assign n3560 = n5521 | (n_n9537 & n4891 & n4967);
  assign n3565 = n5519_1 | n5520;
  assign n3570 = ~preset & (n_n6988 | (ngfdn_3 & ~ndn3_50));
  assign n3575 = ~preset & (n_n6986 | (ndn3_39 & ~ndn3_40));
  assign n3580 = n5518 | n5517 | (n_n8933 & n4898);
  assign n3585 = ~preset & (n_n7117 | (ndn3_39 & ~ndn3_40));
  assign n3590 = n5516 | (n_n9284 & n4845 & n4967);
  assign n3595 = ~n4956 & ~preset & n_n8241;
  assign n3600 = n5515 | (n1270 & (n4971 ^ n4972));
  assign n3605 = ~n4956 & ~preset & n_n8198;
  assign n3610 = n5513 | n5514_1;
  assign n3615 = ~n4956 & ~preset & n_n8575;
  assign n3620 = ~n4956 & ~preset & n_n8710;
  assign n3625 = ~preset & (n_n7622 | (nen3_22 & ~ndn3_22));
  assign n3630 = n5512 | (n_n8557 & n4845 & n4967);
  assign n3635 = n5511 | (n_n8449 & n4890 & n4967);
  assign n3640 = ~preset & (n_n7033 | (~ndn3_46 & ndn3_44));
  assign n3645 = ~preset & ~ngfdn_3 & (ndn3_34 | nen3_34);
  assign n3650 = n5510 | (n_n9512 & n4883 & n4967);
  assign n3655 = ndn3_50 & ~preset & ~ngfdn_3;
  assign n3660 = n5509_1 | (n_n9416 & n4883 & n4967);
  assign n3665 = ~preset & (n_n7019 | (ndn3_42 & ~ndn3_44));
  assign n3670 = n5508 | (n4861 & n4868);
  assign n3675 = ~preset & (n_n7261 | (~ngfdn_3 & ndn3_46));
  assign n3680 = n5507 | (ndn3_29 & ~ndn3_32 & n4855);
  assign n3685 = n5505 | n5506;
  assign n3690 = ~preset & (n4876 ? n4903 : n_n7993);
  assign n3695 = n5503 | n5504_1;
  assign n3700 = n5501 | n5502;
  assign n3705 = n5499_1 | n5500;
  assign n3710 = n5497 | n5498;
  assign n3715 = ~preset & (n_n8918 | (~ndn3_42 & ndn3_40));
  assign n3720 = ~preset & (n4882 ? n4904_1 : n_n8515);
  assign n3725 = ~preset & (n4875 ? n4904_1 : n_n7933);
  assign n3730 = ~preset & (n4847 ? n4930 : n_n8075);
  assign n3735 = ~preset & (n_n7338 | (nen3_22 & ~ndn3_22));
  assign n3740 = ~preset & (n4882 ? n4930 : n_n8104);
  assign n3745 = ~n4956 & ~preset & n_n8171;
  assign n3750 = n5496 | (n_n8707 & n4890 & n4967);
  assign n3755 = n5494_1 | n5495;
  assign n3760 = n5492 | n5493;
  assign n3765 = ~n4956 & ~preset & n_n9441;
  assign n3770 = n5490 | n5491;
  assign n3775 = ~preset & (n_n8831 | (ndn3_39 & ~ndn3_40));
  assign n3780 = ~preset & (n_n8441 | (ndn3_39 & ~ndn3_40));
  assign n3785 = n5489_1 | (n4846 & n4903);
  assign n3790 = n5487 | n5488;
  assign n3795 = ~n4956 & ~preset & n_n9363;
  assign n3800 = ~preset & ~ngfdn_3 & (ndn3_4 | ndn3_2);
  assign n3805 = n5485 | n5486;
  assign n3810 = ~preset & (n_n7561 | (~ngfdn_3 & ndn3_46));
  assign n3815 = n5484_1 | n5483 | (n_n8923 & n4898);
  assign n3820 = ~preset & (n_n7978 | (ndn3_39 & ~ndn3_40));
  assign n3825 = n5482 | n5481 | (n_n8978 & n4898);
  assign n3830 = ~preset & (n4879_1 ? n4868 : n_n9499);
  assign n3835 = ~preset & (n_n8713 | (~ndn3_46 & ndn3_44));
  assign n3840 = ~preset & (n_n8944 | (~ndn3_46 & ndn3_44));
  assign n3845 = ~n4956 & ~preset & n_n8239;
  assign n3850 = ~preset & (n4889_1 ? n4930 : n_n7652);
  assign n3855 = n5479_1 | n5480;
  assign n3860 = ~n4956 & ~preset & n_n8530;
  assign n3865 = n5477 | n5478;
  assign n3870 = n5475 | n5476;
  assign n3875 = n5474_1 | (n4848 & n4861);
  assign n3880 = n5472 | n5473;
  assign n3885 = n5471 | (~ndn3_34 & nen3_34 & n4855);
  assign n3890 = n5469_1 | n5470;
  assign n3895 = n5467 | n5468;
  assign n3900 = n5466 | (~ndn3_27 & ndn3_26 & n4873);
  assign n3905 = n5464_1 | n5465;
  assign n3910 = ~n4956 & ~preset & n_n7961;
  assign n3915 = n5462 | n5463;
  assign n3920 = n5460 | n5461;
  assign n3925 = n5459_1 | (n4861 & (n4969_1 ^ n4970));
  assign n3930 = n5458 | (n4863 & (n4954_1 ^ n4955));
  assign n3935 = ~preset & (n_n9161 | n4956);
  assign n3940 = n5456 | n5457;
  assign n3945 = n5454_1 | n5455;
  assign n3950 = n5452 | n5453;
  assign n3955 = n5450 | n5451;
  assign n3960 = ~n4956 & ~preset & n_n9360;
  assign n3965 = n5449_1 | (ndn3_25 & ~ndn3_26 & n4855);
  assign n3970 = ~preset & (n_n8392 | (~ndn3_42 & ndn3_40));
  assign n3975 = n5448 | n5447 | (n_n9034 & n4898);
  assign n3980 = ~preset & (n4879_1 ? n4887 : n_n8375);
  assign n3985 = n5446 | (n_n9416 & n4845 & n4967);
  assign n3990 = ~n4956 & ~preset & n_n9298;
  assign n3995 = n5444_1 | n5445;
  assign n4000 = n5442 | n5443;
  assign n4005 = ~nsr1_2 & ~preset & ~pdn;
  assign n4009 = n5440 | n5441;
  assign n4014 = n5438 | n5439_1;
  assign n4019 = ~n4956 & ~preset & n_n9291;
  assign n4024 = n5436 | n5437;
  assign n4029 = n5435 | (ndn3_11 & ~ndn3_12 & n4878);
  assign n4034 = n5433 | n5434_1;
  assign n4039 = n5432 | (n_n9353 & n4883 & n4967);
  assign n4044 = n5430 | n5431;
  assign n4049 = n5428 | n5429_1;
  assign n4054 = n5426 | n5427;
  assign n4059 = ~preset & (n4885 ? n4887 : n_n9351);
  assign n4064 = n5425 | (n_n9638 & n4864_1 & n4967);
  assign n4069 = n_n8668 & ~n4862;
  assign n4074 = n5423 | n5424_1;
  assign n4079 = ~preset & (n_n7013 | (~ngfdn_3 & ndn3_46));
  assign n4084 = n5422 | (n1270 & n4930);
  assign n4089 = ~n4956 & ~preset & n_n8200;
  assign n4094 = n5421 | (n1270 & n4903);
  assign n4099 = ~n4956 & ~preset & n_n8803;
  assign n4104 = n5419_1 | n5420;
  assign n4109 = ~n4956 & ~preset & n_n8366;
  assign n4114 = n5417 | n5418;
  assign n4119 = ~n4956 & ~preset & n_n8650;
  assign n4124 = ~n4956 & ~preset & n_n8574;
  assign n4129 = ~preset & (n_n7276 | (nen3_22 & ~ndn3_22));
  assign n4134 = n5415 | n5416;
  assign n4139 = n5413 | n5414_1;
  assign n4144 = ~preset & ~nsr3_35;
  assign n4149 = n5409_1 | n5410 | n5411 | n5412;
  assign n4154 = ~preset & ~ngfdn_3 & (ndn3_46 | ndn3_44);
  assign n4159 = n5407 | n5408;
  assign n4164 = n5405 | n5406;
  assign n4169 = n5403 | n5404_1;
  assign n4174 = ~n4956 & ~preset & n_n9359;
  assign n4179 = ~preset & (n4892 ? n4904_1 : n_n8425);
  assign n4184 = n5402 | (n4846 & (n4969_1 ^ n4970));
  assign n4189 = n5401 | (n4853 & (n4954_1 ^ n4955));
  assign n4194 = n5397 | n5398 | n5399_1 | n5400;
  assign n4199 = n5393 | n5394_1 | n5395 | n5396;
  assign n4204 = n5392 | (~ndn3_25 & ndn3_22 & n4878);
  assign n4209 = ~preset & (n_n7467 | (~ndn3_42 & ndn3_40));
  assign n4214 = n5390 | n5391;
  assign n4219 = n5389_1 | (n4866 & n4904_1);
  assign n4224 = n5388 | (n_n8557 & n4886 & n4967);
  assign n4229 = ~preset & (n_n9162 | n4956);
  assign n4234 = n5387 | (~ndn3_4 & ndn3_2 & n4878);
  assign n4239 = ~preset & (n_n8055 | (~ngfdn_3 & ndn3_46));
  assign n4244 = n5386 | (n_n8354 & n4867 & n4967);
  assign n4249 = n5385 | (n1270 & (n4969_1 ^ n4970));
  assign n4254 = n5384_1 | (n_n9512 & n4896 & n4967);
  assign n4259 = ~preset & (n4875 ? n4848 : n_n7762);
  assign n4264 = n5382 | n5383;
  assign n4269 = n5380 | n5381;
  assign n4274 = n5379_1 | (n_n9416 & n4890 & n4967);
  assign n4279 = n5377 | n5378;
  assign n4284 = n5375 | n5376;
  assign n4289 = n5373 | n5374_1;
  assign n4294 = n5371 | n5372;
  assign n4299 = n5369_1 | n5370;
  assign n4304 = ~preset & (n4885 ? n4903 : n_n9100);
  assign n4309 = n5368 | (n_n9353 & n4864_1 & n4967);
  assign n4314 = n5367 | (n_n9537 & n4864_1 & n4967);
  assign n4319 = ~preset & (n4865 ? n4887 : n_n7588);
  assign n4324 = ~preset & (n_n9123 | (ngfdn_3 & ~ndn3_50));
  assign n4329 = n5366 | (~ndn3_28 & nen3_28 & n4888);
  assign n4334 = n5365 | (nen3_36 & ~ndn3_36 & n4850);
  assign n4339 = n5363 | n5364_1;
  assign n4344 = n5362 | (n4866 & n4930);
  assign n4349 = n5360 | n5361;
  assign n4354 = n5359_1 | (n4866 & n4903);
  assign n4359 = n5357 | n5358;
  assign n4364 = n5356 | (n_n9353 & n4896 & n4967);
  assign n4369 = n5355 | (n4861 & (n4985 ^ n4986));
  assign n4374 = ~n4956 & ~preset & n_n8571;
  assign n4379 = ~n4956 & ~preset & n_n8796;
  assign n4384 = ~preset & ~ngfdn_3 & (nen3_36 | ndn3_36);
  assign n4389 = n5354_1 | (n_n8354 & n4864_1 & n4967);
  assign n4394 = n5352 | n5353;
  assign n4399 = ~preset & (n_n8817 | (ndn3_42 & ~ndn3_44));
  assign n4404 = ~preset & (n_n9160 | n4956);
  assign n4409 = n5351 | (n_n8449 & n4896 & n4967);
  assign n4414 = ~preset & (n4869_1 ? n4904_1 : n_n8513);
  assign n4419 = n5349_1 | n5350;
  assign n4424 = n5348 | (ndn3_25 & ~ndn3_26 & n4878);
  assign n4429 = n7206 | (~preset & n_n9284 & ~n5001);
  assign n4434 = n5346 | n5347;
  assign n4439 = n5345 | (~ndn3_29 & ndn3_28 & n4855);
  assign n4444 = ~preset & (n4851 ? n4904_1 : n_n9203);
  assign n4449 = ~preset & (n4879_1 ? n4930 : n_n7655);
  assign n4454 = ~preset & (n_n8946 | (ndn3_39 & ~ndn3_40));
  assign n4459 = ~preset & (n_n7052 | (~ndn3_46 & ndn3_44));
  assign n4464 = ~preset & (n4851 ? n4848 : n_n9615);
  assign n4469 = n5344_1 | (~ndn3_25 & ndn3_22 & n4855);
  assign n4474 = ~preset & (n4875 ? n4903 : n_n7741);
  assign n4479 = n5342 | n5343;
  assign n4484 = ~preset & (n4877 ? n4904_1 : n_n7912);
  assign n4489 = n5341 | (n1270 & n4868);
  assign n4494 = ~preset & (n4875 ? n4887 : n_n9021);
  assign n4499 = n5339_1 | n5340;
  assign n4504 = n5338 | (nen3_16 & ~ndn3_16 & n4855);
  assign n4509 = n5336 | n5337;
  assign n4514 = n5334_1 | n5335;
  assign n4519 = n5333 | (ndn3_9 & ~ndn3_11 & n4873);
  assign n4524 = n5331 | n5332;
  assign n4529 = ~preset & (n4847 ? n4887 : n_n7694);
  assign n4534 = n5330 | (n_n9448 & n4891 & n4967);
  assign n4539 = n5328 | n5329_1;
  assign n4544 = ~preset & (n4879_1 ? n4904_1 : n_n7935);
  assign n4549 = n5326 | n5327;
  assign n4554 = ~n4956 & ~preset & n_n7701;
  assign n4559 = ~preset & (n4877 ? n4930 : n_n7510);
  assign n4564 = ~n4956 & ~preset & n_n7627;
  assign n4569 = n5324_1 | n5325;
  assign n4574 = ~preset & (n4849_1 ? n4904_1 : n_n8516);
  assign n4579 = ~preset & (n4847 ? n4904_1 : n_n7913);
  assign n4584 = n5323 | (n_n9284 & n4883 & n4967);
  assign n4589 = ~preset & (n_n7411 | (ndn3_39 & ~ndn3_40));
  assign n4594 = n5322 | (~ndn3_27 & ndn3_26 & n4850);
  assign n4599 = n5320 | n5321;
  assign n4604 = n5318 | n5319_1;
  assign n4609 = n5316 | n5317;
  assign n4614 = ~preset & (n_n7242 | (ndn3_42 & ~ndn3_44));
  assign n4619 = ~preset & (n_n8230 | (ndn3_42 & ~ndn3_44));
  assign n4624 = ~n4956 & ~preset & n_n9294;
  assign n4629 = n5315 | (n4863 & n4930);
  assign n4634 = ~n4956 & ~preset & n_n8972;
  assign n4639 = n5313 | n5314_1;
  assign n4644 = ~preset & (n_n7493 | (ngfdn_3 & ~ndn3_50));
  assign n4649 = ~preset & (n_n8290 | (ngfdn_3 & ~ndn3_50));
  assign n4654 = n5309_1 | n5310 | n5311 | n5312;
  assign n4659 = ~n4956 & ~preset & n_n7769;
  assign n4664 = ~preset & (n_n7491 | (~ndn3_46 & ndn3_44));
  assign n4669 = n5307 | n5308;
  assign n4674 = n5305 | n5306;
  assign n4679 = ~preset & (n_n8047 | (ndn3_39 & ~ndn3_40));
  assign n4684 = n5303 | n5304_1;
  assign n4689 = n5302 | (ndn3_29 & ~ndn3_32 & n4850);
  assign n4694 = n5300 | n5301;
  assign n4699 = n5299_1 | (n4846 & n4848);
  assign n4704 = ~n4956 & ~preset & n_n8528;
  assign n4709 = ~preset & ~nsr3_37;
  assign n4714 = ~preset & ~ngfdn_3 & (ndn3_42 | ndn3_40);
  assign n4719 = ~n4956 & ~preset & n_n9358;
  assign n4724 = n5297 | n5298;
  assign n4729 = ~preset & ~ngfdn_3 & (~nsr3_30 | nen3_28);
  assign n4734 = n5296 | (~ndn3_28 & nen3_28 & n4878);
  assign n4739 = ~preset & (n_n7903 | (ndn3_42 & ~ndn3_44));
  assign n4744 = n5294_1 | n5295;
  assign n4749 = ~preset & (n4892 ? n4930 : n_n9075);
  assign n4754 = ~n4956 & ~preset & n_n9439;
  assign n4759 = n7209 | n5292 | n5293;
  assign n4764 = n5290 | n5291;
  assign n4769 = n5289_1 | n5288 | (n_n8798 & n4898);
  assign n4774 = ~preset & (n_n7146 | (~ndn3_46 & ndn3_44));
  assign n4779 = n5286 | n5287;
  assign n4784 = ~preset & (n_n7176 | (~ngfdn_3 & ndn3_46));
  assign n4789 = n5285 | (n_n8652 & n4845 & n4967);
  assign n4794 = ~preset & (n4865 ? n4904_1 : n_n8514);
  assign n4799 = n5284_1 | (n_n8707 & n4845 & n4967);
  assign n4804 = ~preset & (n_n7183 | (ndn3_39 & ~ndn3_40));
  assign n4809 = n5283 | (n_n8419 & n4886 & n4967);
  assign n4814 = n5282 | (n4866 & n4868);
  assign n4819 = n5281 | (n_n8557 & n4891 & n4967);
  assign n4824 = n5279_1 | n5280;
  assign n4829 = n5278 | (n_n8549 & n4891 & n4967);
  assign n4834 = n5276 | n5277;
  assign n4839 = n5275 | (n_n8449 & n4891 & n4967);
  assign n4844 = n5273 | n5274_1;
  assign n4849 = n5271 | n5272;
  assign n4854 = n5269_1 | n5270;
  assign n4859 = n5267 | n5268;
  assign n4864 = n5265 | n5266;
  assign n4869 = n5264_1 | n5263 | (n_n9011 & n4898);
  assign n4874 = n5261 | n5262;
  assign n4879 = n5259_1 | n5260;
  assign n4884 = n5257 | n5258;
  assign n4889 = n5255 | n5256;
  assign n4894 = ~preset & (n_n9164 | n4956);
  assign n4899 = n5253 | n5254_1;
  assign n4904 = n5251 | n5252;
  assign n4909 = n5249_1 | n5250;
  assign n4914 = n5248 | (~ndn3_4 & ndn3_2 & n4873);
  assign n4919 = n5247 | (~ndn3_34 & nen3_34 & n4850);
  assign n4924 = ~n4956 & ~preset & n_n7768;
  assign n4929 = n5245 | n5246;
  assign n4934 = n5244_1 | (n4861 & n4930);
  assign n4939 = n5242 | n5243;
  assign n4944 = n5241 | (n_n9434 & n4891 & n4967);
  assign n4949 = n5239_1 | n5240;
  assign n4954 = n5238 | (n4853 & n4930);
  assign n4959 = n5237 | (n_n9638 & n4891 & n4967);
  assign n4964 = n5235 | n5236;
  assign n4969 = n5233 | n5234_1;
  assign n4974 = ~preset & (n_n9228 | (~ngfdn_3 & ndn3_46));
  assign n4979 = n5232 | (~nsr3_13 & ~ndn3_15 & n4850);
  assign n4984 = ~preset & (n_n8510 | (~ndn3_42 & ndn3_40));
  assign n4989 = ~preset & (n4869_1 ? n4868 : n_n8881);
  assign n4994 = n5231 | (~ndn3_7 & ndn3_4 & n4850);
  assign n4999 = n5229_1 | n5230;
  assign n5004 = n5228 | n5227 | (n_n9031 & n4898);
  assign n5009 = n7210 | (~nak3_13 & nsr3_37);
  assign n5014 = ~n4956 & ~preset & n_n8197;
  assign n5019 = n5225 | n5226;
  assign n5024 = n5223 | n5224_1;
  assign n5029 = n5221 | n5222;
  assign n5034 = ~preset & ~ngfdn_3 & (ndn3_42 | ndn3_44);
  assign n5039 = n5219_1 | n5220;
  assign n5044 = n5218 | (n_n9448 & n4864_1 & n4967);
  assign n5049 = n5216 | n5217;
  assign n5054 = ~preset & ~pdn & (nsr1_2 | nlc1_2);
  assign n5059 = n5214_1 | n5215;
  assign n5064 = ~n4956 & ~preset & n_n8577;
  assign n5069 = ~preset & (n_n7079 | (ndn3_42 & ~ndn3_44));
  assign n5074 = ~preset & (n4869_1 ? n4930 : n_n8828);
  assign n5079 = n5213 | (n_n9638 & n4867 & n4967);
  assign n5084 = n5211 | n5212;
  assign n5089 = ~preset & (n4874_1 ? n4848 : n_n7901);
  assign n5094 = n5209_1 | n5210;
  assign n5099 = n5208 | n5207 | (n_n8869 & n4898);
  assign n5104 = ~preset & (n4859_1 ? n4848 : n_n7710);
  assign n5109 = n5206 | n5205 | (n_n8993 & n4898);
  assign n5114 = ~preset & (n4885 ? n4904_1 : n_n9586);
  assign n5119 = ~preset & (n4889_1 ? n4848 : n_n8852);
  assign n5124 = n5204_1 | (~ndn3_17 & ndn3_16 & n4878);
  assign n5129 = n5202 | n5203;
  assign n5134 = ~preset & (n_n7717 | (ndn3_39 & ~ndn3_40));
  assign n5139 = n5201 | (n_n8821 & n4845 & n4967);
  assign n5144 = ~preset & (n_n9163 | n4956);
  assign n5149 = n5200 | (n_n8557 & n4883 & n4967);
  assign n5154 = n5198 | n5199_1;
  assign n5159 = n5196 | n5197;
  assign n5164 = n5194_1 | n5195;
  assign n5169 = n5192 | n5193;
  assign n5174 = n5191 | (n_n8652 & n4890 & n4967);
  assign n5179 = n5190 | (~ndn3_25 & ndn3_22 & n4888);
  assign n5184 = n5188 | n5189_1;
  assign n5189 = n5187 | (n_n9512 & n4890 & n4967);
  assign n5194 = n5185 | n5186;
  assign n5199 = n5184_1 | (~ndn3_17 & ndn3_16 & n4873);
  assign n5204 = n5182 | n5183;
  assign n5209 = ~preset & (n_n7330 | (ndn3_39 & ~ndn3_40));
  assign n5214 = n5180 | n5181;
  assign n5219 = n5178 | n5179_1;
  assign n5224 = n5177 | n5176 | (n_n8847 & n4898);
  assign n5229 = n5174_1 | n5175;
  assign n5234 = ~preset & (n4874_1 ? n4903 : n_n7553);
  assign n5239 = ~n4956 & ~preset & n_n9292;
  assign n5244 = ~preset & (n4854_1 ? n4887 : n_n7464);
  assign n5249 = n5172 | n5173;
  assign n5254 = n5170 | n5171;
  assign n5259 = n5169_1 | (n_n9434 & n4883 & n4967);
  assign n5264 = ~n4956 & ~preset & n_n8118;
  assign n5269 = n5168 | (n4846 & n4930);
  assign n5274 = n5167 | (n4861 & n4903);
  assign n5279 = n5166 | (n4861 & (n4971 ^ n4972));
  assign n5284 = n5165 | (n_n9434 & n4864_1 & n4967);
  assign n5289 = ~preset & ~ngfdn_3 & (ndn3_2 | n4949_1);
  assign n5294 = n5164_1 | (n_n8652 & n4867 & n4967);
  assign n5299 = n5162 | n5163;
  assign n5304 = n5160 | n5161;
  assign n5309 = ~preset & (n_n8665 | (ngfdn_3 & ~ndn3_50));
  assign n5314 = n5158 | n5159_1;
  assign n5319 = n5156 | n5157;
  assign n5324 = n5154_1 | n5155;
  assign n5329 = ~preset & (n4876 ? n4868 : n_n9173);
  assign n5334 = n5152 | n5153;
  assign n5339 = ~preset & (n_n7150 | (~ndn3_42 & ndn3_40));
  assign n5344 = n5151 | (nen3_36 & ~ndn3_36 & n4888);
  assign n5349 = n5149_1 | n5150;
  assign n5354 = n7211 | (~ndn3_17 & nsr3_20);
  assign n5359 = ~n4956 & ~preset & n_n8271;
  assign n5364 = n5147 | n5148;
  assign n5369 = n5146 | (n4853 & n4904_1);
  assign n5374 = ~preset & ~ngfdn_3 & (ndn3_39 | ndn3_40);
  assign n5379 = n5144_1 | n5145;
  assign n5384 = n5143 | (~ndn3_4 & ndn3_2 & n4888);
  assign n5389 = n5141 | n5142;
  assign n5394 = n5139_1 | n5140;
  assign n5399 = ~preset & (n4885 ? n4868 : n_n8462);
  assign n5404 = n5137 | n5138;
  assign n5409 = n5135 | n5136;
  assign n5414 = ~n4956 & ~preset & n_n9289;
  assign n5419 = ~preset & (n4881 ? n4930 : n_n7661);
  assign n5424 = n5133 | n5134_1;
  assign n5429 = ~preset & (n_n8921 | (~ndn3_46 & ndn3_44));
  assign n5434 = n5132 | (~ndn3_28 & nen3_28 & n4855);
  assign n5439 = n5131 | (n_n9448 & n4896 & n4967);
  assign n5444 = n5129_1 | n5130;
  assign n5449 = n5128 | (n4866 & (n4985 ^ n4986));
  assign n5454 = n5126 | n5127;
  assign n5459 = n5124_1 | n5125;
  assign n5464 = n5123 | (n_n8449 & n4867 & n4967);
  assign n5469 = n5121 | n5122;
  assign n5474 = n5120 | (n_n8419 & n4867 & n4967);
  assign n5479 = ~preset & (n_n7336 | (~ngfdn_3 & ndn3_46));
  assign n5484 = n5119_1 | (~ndn3_17 & ndn3_16 & n4855);
  assign n5489 = n5117 | n5118;
  assign n5494 = n5115 | n5116;
  assign n5499 = n5113 | n5114_1;
  assign n5504 = ~preset & (n_n8423 | (nen3_22 & ~ndn3_22));
  assign n5509 = ~preset & (n4881 ? n4848 : n_n7763);
  assign n5514 = n5112 | (n_n8419 & n4891 & n4967);
  assign n5519 = n5110 | n5111;
  assign n5524 = n5108 | n5109_1;
  assign n5529 = n5106 | n5107;
  assign n5534 = n5104_1 | n5105;
  assign n5539 = n5103 | (~ndn3_9 & ndn3_7 & n4855);
  assign n5544 = ~preset & (n4852 ? n4903 : n_n9563);
  assign n5549 = ~preset & (n_n8672 | (ngfdn_3 & ~ndn3_50));
  assign n5554 = ~preset & (n4854_1 ? n4930 : n_n7346);
  assign n5559 = n5102 | (n_n8821 & n4890 & n4967);
  assign n5564 = ~n4956 & ~preset & n_n8756;
  assign n5569 = ~preset & (n4874_1 ? n4930 : n_n8641);
  assign n5574 = n5100 | n5101;
  assign n5579 = n5099_1 | (ndn3_17 & ~ndn3_18 & n4873);
  assign n5584 = n5098 | n5097 | (n_n8561 & n4898);
  assign n5589 = ~preset & (n_n9306 | (ngfdn_3 & ~ndn3_50));
  assign n5594 = ~preset & (n_n9165 | n4956);
  assign n5599 = n5095 | n5096;
  assign n5604 = ~preset & (n4847 ? n4848 : n_n9210);
  assign n5609 = ~n4901 & ~preset & ndn2_2;
  assign n5614 = ~preset & (n4865 ? n4930 : n_n7342);
  assign n5619 = n5093 | n5094_1;
  assign n5624 = n5092 | (n4846 & (n4971 ^ n4972));
  assign n5629 = n5090 | n5091;
  assign n5634 = ~preset & (n_n9006 | (ndn3_42 & ~ndn3_44));
  assign n5639 = n5089_1 | (n_n8652 & n4886 & n4967);
  assign n5644 = ~preset & (n_n7905 | (ndn3_42 & ~ndn3_44));
  assign n5649 = ~preset & (n_n9166 | n4956);
  assign n5654 = ~preset & (n_n7065 | (ndn3_42 & ~ndn3_44));
  assign n5659 = ~preset & (n4892 ? n4868 : n_n9490);
  assign n5664 = ~preset & (n_n7024 | (~ndn3_42 & ndn3_40));
  assign n5669 = ~preset & (n_n7586 | (~ngfdn_3 & ndn3_46));
  assign n5674 = n5087 | n5088;
  assign n5679 = n5085 | n5086;
  assign n5684 = ~n4956 & ~preset & n_n8141;
  assign n5689 = ~n4956 & ~preset & n_n7853;
  assign n5694 = ~preset & (n_n8121 | (~ndn3_42 & ndn3_40));
  assign n5699 = n5083 | n5084_1;
  assign n5704 = ~preset & (n4849_1 ? n4868 : n_n9496);
  assign n5709 = ~preset & (n_n8195 | (ndn3_42 & ~ndn3_44));
  assign n5714 = ~preset & (n4860 ? n4848 : n_n9516);
  assign n5719 = n5082 | (~ndn3_27 & ndn3_26 & n4878);
  assign n5724 = ~n4956 & ~preset & n_n9436;
  assign n5729 = n5080 | n5081;
  assign n5734 = n5078 | n5079_1;
  assign n5739 = n5074_1 | n5075 | n5076 | n5077;
  assign n5744 = n5073 | (n_n9416 & n4864_1 & n4967);
  assign n5749 = n5072 | (ndn3_9 & ~ndn3_11 & n4850);
  assign n5754 = n5071 | (n_n9353 & n4890 & n4967);
  assign n5759 = ~n4956 & ~preset & n_n7770;
  assign n5764 = ~preset & ~ngfdn_3 & (ndn3_29 | ndn3_32);
  assign n5769 = n5069_1 | n5070;
  assign n5774 = n5068 | (n4846 & n4868);
  assign n5779 = n5067 | (n4863 & n4904_1);
  assign n5784 = n5065 | n5066;
  assign n5789 = n5063 | n5064_1;
  assign n5794 = n5061 | n5062;
  assign n5799 = ~preset & ~nsr3_38;
  assign n5804 = n5059_1 | n5060;
  assign n5809 = ~preset & (n4847 ? n4868 : n_n9179);
  assign n5814 = ~n4956 & ~preset & n_n9357;
  assign n5819 = n5057 | n5058;
  assign n5824 = ~n4956 & ~preset & n_n7628;
  assign n5829 = ~preset & (n_n8454 | (~ndn3_46 & ndn3_44));
  assign n5834 = ~preset & ~nsr3_20;
  assign n5839 = n5056 | (n_n9448 & n4845 & n4967);
  assign n5844 = ~preset & ~ngfdn_3 & (~nsr3_35 | nen3_34);
  assign n5849 = n5055 | (n4861 & n4904_1);
  assign n5854 = n5053 | n5054_1;
  assign n5859 = n5051 | n5052;
  assign n5864 = n5049_1 | n5050;
  assign n5869 = ~preset & (n_n9578 | n4956);
  assign n5874 = ~preset & (n4860 ? n4903 : n_n8135);
  assign n5879 = ~preset & ~ngfdn_3 & (ndn3_25 | ndn3_26);
  assign n5884 = n5047 | n5048;
  assign n5889 = n5046 | (n4846 & (n4985 ^ n4986));
  assign n5894 = ~preset & (n_n8605 | (~ndn3_46 & ndn3_44));
  assign n5899 = ~n4956 & ~preset & n_n9296;
  assign n5904 = n5044_1 | n5045;
  assign n5909 = n5043 | (n_n9638 & n4890 & n4967);
  assign n5914 = n5041 | n5042;
  assign n5919 = n5040 | (nen3_39 & ~ndn3_39 & n4888);
  assign n5924 = n5038 | n5039_1;
  assign n5929 = ~n4956 & ~preset & n_n9275;
  assign n5934 = n5036 | n5037;
  assign n5939 = n5035 | (n_n9537 & n4890 & n4967);
  assign n5944 = n5033 | n5034_1;
  assign n5949 = n5031 | n5032;
  assign n5954 = ~n4956 & ~preset & n_n7629;
  assign n5959 = ~preset & ~nsr3_14;
  assign n5964 = n5030 | (n4846 & (n4954_1 ^ n4955));
  assign n5969 = ~n4956 & ~preset & n_n9013;
  assign n5974 = n5028 | n5029_1;
  assign n5979 = n5027 | (n_n8557 & n4864_1 & n4967);
  assign n5984 = ~preset & (n4854_1 ? n4848 : n_n7334);
  assign n5989 = ~n4956 & ~preset & n_n7704;
  assign n5994 = n5026 | (n_n8419 & n4845 & n4967);
  assign n5999 = ~preset & (n4859_1 ? n4930 : n_n8526);
  assign n6004 = ~n4956 & ~preset & n_n9556;
  assign n6009 = n5025 | (ndn3_9 & ~ndn3_11 & n4888);
  assign n6014 = ~n4956 & ~preset & n_n8447;
  assign n6019 = n5023 | n5024_1;
  assign n6024 = ~n4956 & ~preset & n_n8570;
  assign n6029 = n5022 | (ndn3_25 & ~ndn3_26 & n4873);
  assign n6034 = n5021 | (n_n8549 & n4864_1 & n4967);
  assign n6039 = ~n4956 & ~preset & n_n8646;
  assign n6044 = n5019_1 | n5020;
  assign n6049 = n5018 | (n1270 & (n4976 ^ n4977));
  assign n6054 = n5017 | (ndn3_17 & ~ndn3_18 & n4850);
  assign n6059 = ~preset & (n_n8216 | (~ndn3_46 & ndn3_44));
  assign n6064 = ~preset & (n4877 ? n4868 : n_n9177);
  assign n6069 = n5015 | n5016;
  assign n6074 = n5014_1 | (~ndn3_17 & ndn3_16 & n4850);
  assign n6079 = n5012 | n5013;
  assign n6084 = n5010 | n5011;
  assign n6089 = ~preset & (n4854_1 ? n4868 : n_n8858);
  assign n6094 = n5009_1 | (~ndn3_34 & nen3_34 & n4878);
  assign n4845 = ~nsr3_37 & ~preset & ~ndn3_37;
  assign n4846 = ~ndn3_40 & ~preset & ndn3_39;
  assign n4847 = ndn3_9 & ~ndn3_11;
  assign n4848 = n5002 ? ((~n4988 & ~n4989_1) | (~n4976 & (~n4989_1 | (~n4988 & n4989_1)))) : ((n4988 & n4989_1) | (n4976 & (n4988 ^ n4989_1)));
  assign n4849_1 = ndn3_11 & ~ndn3_12;
  assign n4850 = ~preset & (n4996 ^ (n6545 | n6546));
  assign n4851 = ndn3_25 & ~ndn3_26;
  assign n4852 = ~ndn3_9 & ndn3_7;
  assign n4853 = ndn3_44 & ~preset & ~ndn3_46;
  assign n4854_1 = nen3_39 & ~ndn3_39;
  assign n4855 = ~preset & (n4980 ^ (n6352 | n6353));
  assign n4856 = n_n9247 & n_n9248 & ~preset & ~n_n7306;
  assign n4857 = n4856 & n5001;
  assign n4858 = n4998 ? ((n4905 & n4906) | (n_n8549 & (n4905 | n4906))) : ((~n4905 & ~n4906) | (~n_n8549 & (~n4905 | ~n4906)));
  assign n4859_1 = ~ndn3_27 & ndn3_26;
  assign n4860 = ~ndn3_34 & nen3_34;
  assign n4861 = ~ndn3_44 & ~preset & ndn3_42;
  assign n4862 = ~n_n9198 | preset | (~n4967 & n4974_1);
  assign n4863 = ndn3_40 & ~preset & ~ndn3_42;
  assign n4864_1 = ~ndn3_35 & ~preset & ~nsr3_35;
  assign n4865 = ~ndn3_19 & nen3_19;
  assign n4866 = ~ndn3_22 & ~preset & nen3_22;
  assign n4867 = ~nsr3_23 & ~preset & ~ndn3_23;
  assign n4868 = n4965 ? ((~n4978 & ~n4979_1) | (~n4972 & (~n4979_1 | (~n4978 & n4979_1)))) : ((n4978 & n4979_1) | (n4972 & (~n4978 ^ ~n4979_1)));
  assign n4869_1 = ~ndn3_29 & ndn3_28;
  assign n4870 = n6282 | n6283 | n6284 | n7095;
  assign n4871 = (n_n8821 & n4934_1) | ((n_n8821 | n4934_1) & (n7112 | n7113));
  assign n4872 = (n_n9638 & n4871) | ((n_n9638 | n4871) & (n7094 | n7095));
  assign n4873 = ~preset & (n5004_1 ^ (n6527 | n6528));
  assign n4874_1 = ~ndn3_4 & ndn3_2;
  assign n4875 = nen3_16 & ~ndn3_16;
  assign n4876 = nen3_36 & ~ndn3_36;
  assign n4877 = ndn3_17 & ~ndn3_18;
  assign n4878 = ~preset & (n4997 ^ (n6083 | n6084_1));
  assign n4879_1 = ~ndn3_7 & ndn3_4;
  assign n4880 = ndn3_29 & ~ndn3_32;
  assign n4881 = ~nsr3_13 & ~ndn3_15;
  assign n4882 = ~ndn3_17 & ndn3_16;
  assign n4883 = ~nsr3_13 & ~preset & ~ndn3_13;
  assign n4884_1 = pdn ? ~ndn1_4 : ~nsr1_2;
  assign n4885 = ndn3_19 & ~ndn3_21;
  assign n4886 = ~ndn3_20 & ~preset & ~nsr3_20;
  assign n4887 = n4966 ? ((~n5007 & ~n5008) | (~n4969_1 & (~n5008 | (~n5007 & n5008)))) : ((n5007 & n5008) | (n4969_1 & (~n5007 ^ ~n5008)));
  assign n4888 = ~preset & (n4987 ^ (n6433 | n6434));
  assign n4889_1 = ~ndn3_25 & ndn3_22;
  assign n4890 = ~ndn3_38 & ~preset & ~nsr3_38;
  assign n4891 = ~ndn3_14 & ~preset & ~nsr3_14;
  assign n4892 = ~ndn3_28 & nen3_28;
  assign n4893 = n6261 | n6262 | n6263 | n7097;
  assign n4894_1 = (n_n9512 & n4919_1) | ((n_n9512 | n4919_1) & (n7098 | n7099));
  assign n4895 = (n_n9434 & n4894_1) | ((n_n9434 | n4894_1) & (n7096 | n7097));
  assign n4896 = ~nsr3_30 & ~preset & ~ndn3_30;
  assign n4897 = n6857 | n6858;
  assign n4898 = ~preset & (n4975 ? n4967 : ~n5001);
  assign n4899_1 = ~n_n8631 ^ (n_n8561 | n4999_1);
  assign n4900 = n6859 | n6860;
  assign n4901 = ~nlc1_2 & preset_0_0_ & nsr1_2;
  assign n4902 = n7173 & n7172 & ~n4907 & ~n4940;
  assign n4903 = n4973 ? ((~n4981 & ~n4982) | (~n4955 & (~n4982 | (~n4981 & n4982)))) : ((n4981 & n4982) | (n4955 & (~n4981 ^ ~n4982)));
  assign n4904_1 = n4952 ? ((~n4994_1 & ~n4995) | (~n4986 & (~n4995 | (~n4994_1 & n4995)))) : ((n4994_1 & n4995) | (n4986 & (~n4994_1 ^ ~n4995)));
  assign n4905 = n6303 | n6304 | n6305 | n7091;
  assign n4906 = (n_n8449 & n4932) | ((n_n8449 | n4932) & (n7092 | n7093));
  assign n4907 = (~n_n8913 & ~n_n8964 & ~n4968) | (n_n8964 & (n_n8913 | n4968));
  assign n4908 = n6861 | n6862;
  assign n4909_1 = n_n8652 & (n7100 | n7101);
  assign n4910 = n6233 | n6234 | n6235 | n7101;
  assign n4911 = (n_n9284 & n4909_1) | ((n_n9284 | n4909_1) & (n7102 | n7103));
  assign n4912 = (n_n8707 & n4911) | ((n_n8707 | n4911) & (n7104 | n7105));
  assign n4913 = n6226 | n6227 | n6228 | n7105;
  assign n4914_1 = (n_n8354 & n4915) | ((n_n8354 | n4915) & (n7116 | n7117));
  assign n4915 = (n_n9448 & n4872) | ((n_n9448 | n4872) & (n7114 | n7115));
  assign n4916 = n6212 | n6213 | n6214 | n7117;
  assign n4917 = n6863 | n6864;
  assign n4918 = n6254 | n6255 | n6256 | n7099;
  assign n4919_1 = (n_n9353 & n4912) | ((n_n9353 | n4912) & (n7106 | n7107));
  assign n4920 = (n_n9353 & (n4912 | n4938)) | n4918 | (n4912 & n4938);
  assign n4921 = n6268 | n6269 | n6270 | n7109;
  assign n4922 = (n_n9416 & n4895) | ((n_n9416 | n4895) & (n7108 | n7109));
  assign n4923 = n6867 | n6868;
  assign n4924_1 = (n_n8923 & (~n_n8603 | n_n8798)) | (n_n8603 & ~n_n8923 & ~n_n8798);
  assign n4925 = n6869 | n6870;
  assign n4926 = n6871 | n6872;
  assign n4927 = (~n_n8911 & ~n_n8933 & ~n_n8978 & ~n5000) | (n_n8978 & (n_n8911 | n_n8933 | n5000));
  assign n4928 = (~n_n9034 & ~n_n9031 & ~n_n8993 & ~n5005) | (n_n9034 & (n_n9031 | n_n8993 | n5005));
  assign n4929_1 = n6873 | n6874;
  assign n4930 = (~n6992 & ~n6993 & (n6999 | n7000)) | (~n6999 & ~n7000 & (n6992 | n6993));
  assign n4931 = n6296 | n6297 | n6298 | n7093;
  assign n4932 = (n_n8419 & n4914_1) | ((n_n8419 | n4914_1) & (n7118 | n7119));
  assign n4933 = n6289 | n6290 | n6291 | n7115;
  assign n4934_1 = (n_n9537 & n4922) | ((n_n9537 | n4922) & (n7110 | n7111));
  assign n4935 = n6275 | n6276 | n6277 | n7111;
  assign n4936 = n6240 | n6241 | n6242 | n7103;
  assign n4937 = n6219 | n6220 | n6221 | n7113;
  assign n4938 = n6247 | n6248 | n6249 | n7107;
  assign n4939_1 = n6875 | n6876;
  assign n4940 = (~n_n8913 & ~n_n8964 & ~n_n9011 & ~n4968) | (n_n9011 & (n_n8913 | n_n8964 | n4968));
  assign n4941 = n6877 | n6878;
  assign n4942 = n6879 | n6880;
  assign n4943 = ~n_n9031 ^ (n_n8993 | n5005);
  assign n4944_1 = n6881 | n6882;
  assign n4945 = (n_n8869 & (~n_n8603 | n_n8923 | n_n8798)) | (n_n8603 & ~n_n8923 & ~n_n8798 & ~n_n8869);
  assign n4946 = n6883 | n6884;
  assign n4947 = (~n_n8631 & ~n_n8847 & ~n_n8561 & ~n4999_1) | (n_n8847 & (n_n8631 | n_n8561 | n4999_1));
  assign n4948 = n6885 | n6886;
  assign n4949_1 = nsr1_2 & (nlc1_2 ? n_n7476 : ~preset_0_0_);
  assign n4950 = n6887 | n6888;
  assign n4951 = n6205 | n6206 | n6207 | n7119;
  assign n4952 = (~n7157 & ~n7158 & (n7164 | n7165)) | (~n7164 & ~n7165 & (n7157 | n7158));
  assign n4953 = n_n9247 & ~n_n7306 & n_n9248;
  assign n4954_1 = (~n6978 & ~n6979 & (n6985 | n6986)) | (~n6985 & ~n6986 & (n6978 | n6979));
  assign n4955 = (n6992 | n6993) & (n6999 | n7000);
  assign n4956 = ~ndn2_2 & ~nlc1_2 & preset_0_0_ & nsr1_2;
  assign n4957 = nsr3_13 ? ndn3_12 : nsr3_14;
  assign n4958 = (nen3_36 & ~ndn3_36) | (~ndn3_4 & ndn3_2);
  assign n4959_1 = (~ndn3_29 & ndn3_28) | (nen3_39 & ~ndn3_39);
  assign n4960 = (ndn3_42 & ~ndn3_44) | (~ndn3_34 & nen3_34);
  assign n4961 = (~ndn3_19 & nen3_19) | (~ndn3_28 & nen3_28);
  assign n4962 = (ndn3_39 & ~ndn3_40) | (ndn3_25 & ~ndn3_26);
  assign n4963 = (~ndn3_42 & ndn3_40) | (ndn3_29 & ~ndn3_32);
  assign n4964_1 = (~ndn3_17 & ndn3_16) | (~ndn3_27 & ndn3_26);
  assign n4965 = (~n6922 & ~n6923 & (n6929 | n6930)) | (~n6929 & ~n6930 & (n6922 | n6923));
  assign n4966 = (~n7048 & ~n7049 & (n7055 | n7056)) | (~n7055 & ~n7056 & (n7048 | n7049));
  assign n4967 = n_n8930 ? n_n8929 : (n6897 | n6898);
  assign n4968 = n_n8631 | n_n8847 | n_n8561 | n4999_1;
  assign n4969_1 = (n4992 & n4993) | ((n6527 | n6528) & (~n4992 ^ ~n4993));
  assign n4970 = (~n7006 & ~n7007 & (n7013 | n7014)) | (~n7013 & ~n7014 & (n7006 | n7007));
  assign n4971 = (~n6936 & ~n6937 & (n6943 | n6944)) | (~n6943 & ~n6944 & (n6936 | n6937));
  assign n4972 = (n4990 & n4991) | ((n6545 | n6546) & (~n4990 ^ ~n4991));
  assign n4973 = (~n6964 & ~n6965 & (n6971 | n6972)) | (~n6971 & ~n6972 & (n6964 | n6965));
  assign n4974_1 = n4957 | n7086 | n7087 | n7088;
  assign n4975 = ~n_n8668 & (~n_n9198 | (~n4967 & n4974_1));
  assign n4976 = (n4983 & n4984_1) | ((n6433 | n6434) & (~n4983 ^ ~n4984_1));
  assign n4977 = (~n7020 & ~n7021 & (n7027 | n7028)) | (~n7027 & ~n7028 & (n7020 | n7021));
  assign n4978 = n6665 | n6666 | n6935 | n6937;
  assign n4979_1 = n6651 | n6652 | n6942 | n6944;
  assign n4980 = (~n7076 & ~n7077 & (n7083 | n7084)) | (~n7083 & ~n7084 & (n7076 | n7077));
  assign n4981 = n6593 | n6594 | n6977 | n6979;
  assign n4982 = n6607 | n6608 | n6984 | n6986;
  assign n4983 = n6465 | n6466 | n7033 | n7035;
  assign n4984_1 = n6417 | n6418 | n7040 | n7042;
  assign n4985 = (~n7129 & ~n7130 & (n7136 | n7137)) | (~n7136 & ~n7137 & (n7129 | n7130));
  assign n4986 = (n5003 & n5006) | ((n6352 | n6353) & (~n5003 ^ ~n5006));
  assign n4987 = (~n7034 & ~n7035 & (n7041 | n7042)) | (~n7041 & ~n7042 & (n7034 | n7035));
  assign n4988 = n6387 | n6388 | n7019 | n7021;
  assign n4989_1 = n6401 | n6402 | n7026 | n7028;
  assign n4990 = n6637 | n6638 | n6949 | n6951;
  assign n4991 = n6529 | n6530 | n6956 | n6958;
  assign n4992 = n6711 | n6712 | n6905 | n6907;
  assign n4993 = n6511 | n6512 | n6914 | n6916;
  assign n4994_1 = n6163 | n6164 | n7128 | n7130;
  assign n4995 = n6147 | n6148 | n7135 | n7137;
  assign n4996 = (~n6950 & ~n6951 & (n6957 | n6958)) | (~n6957 & ~n6958 & (n6950 | n6951));
  assign n4997 = (~n7143 & ~n7144 & (n7150 | n7151)) | (~n7150 & ~n7151 & (n7143 | n7144));
  assign n4998 = n6198 | n6199 | n6200 | n7120;
  assign n4999_1 = n_n9034 | n_n9031 | n_n8993 | n5005;
  assign n5000 = ~n_n8603 | n_n8923 | n_n8798 | n_n8869;
  assign n5001 = n_n9247 ? n7085 : (n4967 & n7089);
  assign n5002 = (~n7062 & ~n7063 & (n7069 | n7070)) | (~n7069 & ~n7070 & (n7062 | n7063));
  assign n5003 = n6322 | n6323 | n7075 | n7077;
  assign n5004_1 = (~n6906 & ~n6907 & (n6915 | n6916)) | (~n6915 & ~n6916 & (n6906 | n6907));
  assign n5005 = n_n8911 | n_n8933 | n_n8978 | n5000;
  assign n5006 = n6338 | n6339 | n7082 | n7084;
  assign n5007 = n6497 | n6498 | n7005 | n7007;
  assign n5008 = n6481 | n6482 | n7012 | n7014;
  assign n5009_1 = ~preset & n_n8580 & (ndn3_34 | ~nen3_34);
  assign n5010 = ~preset & n_n8428 & (ndn3_46 | ~ndn3_44);
  assign n5011 = ~ndn3_46 & ~preset & n_n9333 & ndn3_44;
  assign n5012 = ~preset & n_n9145 & (ngfdn_3 | ~ndn3_46);
  assign n5013 = n_n9629 & ndn3_46 & ~preset & ~ngfdn_3;
  assign n5014_1 = ~preset & n_n8811 & (ndn3_17 | ~ndn3_16);
  assign n5015 = ~preset & n_n7844 & (~nen3_36 | ndn3_36);
  assign n5016 = ~preset & n4876 & (~n4985 ^ ~n4986);
  assign n5017 = ~preset & n_n9131 & (~ndn3_17 | ndn3_18);
  assign n5018 = ~preset & n_n8948 & (ngfdn_3 | ~ndn3_46);
  assign n5019_1 = ~ndn3_2 & ~preset & psv26_3_3_ & n4949_1;
  assign n5020 = ~preset & n_n9405 & (ndn3_2 | ~n4949_1);
  assign n5021 = ~preset & n_n7928 & (nsr3_35 | ndn3_35);
  assign n5022 = ~preset & n_n7453 & (~ndn3_25 | ndn3_26);
  assign n5023 = ~preset & n_n7485 & (~ndn3_25 | ndn3_26);
  assign n5024_1 = ~preset & n4851 & (~n4971 ^ ~n4972);
  assign n5025 = ~preset & n_n9345 & (~ndn3_9 | ndn3_11);
  assign n5026 = ~preset & n_n7788 & (ndn3_37 | nsr3_37);
  assign n5027 = ~preset & n_n8078 & (nsr3_35 | ndn3_35);
  assign n5028 = ~preset & n_n7288 & (~ngfdn_3 | ndn3_50);
  assign n5029_1 = ~ndn3_50 & n_n9282 & ~preset & ngfdn_3;
  assign n5030 = ~preset & n_n7862 & (~ndn3_39 | ndn3_40);
  assign n5031 = ~ndn3_2 & ~preset & psv18_9_9_ & n4949_1;
  assign n5032 = ~preset & n_n6976 & (ndn3_2 | ~n4949_1);
  assign n5033 = ~preset & n_n7344 & (~ngfdn_3 | ndn3_50);
  assign n5034_1 = ~ndn3_50 & ~preset & ngfdn_3 & n_n9570;
  assign n5035 = ~preset & n_n9590 & (nsr3_38 | ndn3_38);
  assign n5036 = ~preset & n_n7203 & (ndn3_46 | ~ndn3_44);
  assign n5037 = ~ndn3_46 & ~preset & n_n9125 & ndn3_44;
  assign n5038 = ~ndn3_2 & ~preset & psv38_14_14_ & n4949_1;
  assign n5039_1 = ~preset & n_n8139 & (ndn3_2 | ~n4949_1);
  assign n5040 = ~preset & n_n8991 & (~nen3_39 | ndn3_39);
  assign n5041 = ~preset & n_n8895 & (ngfdn_3 | ~ndn3_46);
  assign n5042 = ndn3_46 & n_n7570 & ~preset & ~ngfdn_3;
  assign n5043 = ~preset & n_n7920 & (nsr3_38 | ndn3_38);
  assign n5044_1 = ~preset & n_n7156 & (~ndn3_42 | ndn3_44);
  assign n5045 = ~ndn3_44 & ndn3_42 & ~preset & n_n8609;
  assign n5046 = ~preset & n_n6974 & (~ndn3_39 | ndn3_40);
  assign n5047 = ~preset & n_n7500 & (~nen3_22 | ndn3_22);
  assign n5048 = ~ndn3_22 & ~preset & nen3_22 & n_n9460;
  assign n5049_1 = ~preset & n_n9048 & (~ndn3_17 | ndn3_18);
  assign n5050 = ~preset & n4877 & (~n4954_1 ^ ~n4955);
  assign n5051 = ~ndn3_2 & ~preset & psv38_7_7_ & n4949_1;
  assign n5052 = ~preset & n_n9262 & (ndn3_2 | ~n4949_1);
  assign n5053 = ~preset & n_n7076 & (~nen3_22 | ndn3_22);
  assign n5054_1 = ~ndn3_22 & ~preset & nen3_22 & n_n8462;
  assign n5055 = ~preset & n_n9632 & (~ndn3_42 | ndn3_44);
  assign n5056 = ~preset & n_n9505 & (ndn3_37 | nsr3_37);
  assign n5057 = ~ndn3_2 & ~preset & psv18_7_7_ & n4949_1;
  assign n5058 = ~preset & n_n9594 & (ndn3_2 | ~n4949_1);
  assign n5059_1 = ~ndn3_2 & ~preset & psv18_13_13_ & n4949_1;
  assign n5060 = ~preset & n_n7886 & (ndn3_2 | ~n4949_1);
  assign n5061 = ~preset & n_n9269 & (ndn3_4 | ~ndn3_2);
  assign n5062 = ~preset & n4874_1 & (~n4969_1 ^ ~n4970);
  assign n5063 = ~preset & n_n7111 & (~ngfdn_3 | ndn3_50);
  assign n5064_1 = ~ndn3_50 & ~preset & ngfdn_3 & n_n9028;
  assign n5065 = ~ndn3_2 & ~preset & psv2_7_7_ & n4949_1;
  assign n5066 = ~preset & n_n9606 & (ndn3_2 | ~n4949_1);
  assign n5067 = ~preset & n_n7927 & (ndn3_42 | ~ndn3_40);
  assign n5068 = ~preset & n_n8206 & (~ndn3_39 | ndn3_40);
  assign n5069_1 = ~preset & n_n7601 & (ndn3_27 | ~ndn3_26);
  assign n5070 = ~preset & n4859_1 & (~n4971 ^ ~n4972);
  assign n5071 = ~preset & n_n9392 & (nsr3_38 | ndn3_38);
  assign n5072 = ~preset & n_n9133 & (~ndn3_9 | ndn3_11);
  assign n5073 = ~preset & n_n7874 & (nsr3_35 | ndn3_35);
  assign n5074_1 = n7212 & ((n4915 & n4916) | (n_n8354 & (n4915 | n4916)));
  assign n5075 = ~n_n8419 & n4857 & (~n4914_1 ^ ~n4951);
  assign n5076 = ~n4951 & ~n4914_1 & n_n8419 & n4856;
  assign n5077 = ~n5001 & ~preset & n_n8419;
  assign n5078 = ~preset & n_n7664 & (~nen3_36 | ndn3_36);
  assign n5079_1 = ~preset & n4876 & (~n4976 ^ ~n4977);
  assign n5080 = ~preset & n_n9051 & (ndn3_9 | ~ndn3_7);
  assign n5081 = ~preset & n4852 & (~n4954_1 ^ ~n4955);
  assign n5082 = ~preset & n_n9077 & (ndn3_27 | ~ndn3_26);
  assign n5083 = ~ndn3_2 & ~preset & psv13_7_7_ & n4949_1;
  assign n5084_1 = ~preset & n_n9604 & (ndn3_2 | ~n4949_1);
  assign n5085 = ~preset & n_n8937 & (ndn3_29 | ~ndn3_28);
  assign n5086 = ~preset & n4869_1 & (~n4969_1 ^ ~n4970);
  assign n5087 = ~ndn3_2 & ~preset & psv39_9_9_ & n4949_1;
  assign n5088 = ~preset & n_n8416 & (ndn3_2 | ~n4949_1);
  assign n5089_1 = ~preset & n_n7653 & (nsr3_20 | ndn3_20);
  assign n5090 = ~ndn3_2 & ~preset & psv33_9_9_ & n4949_1;
  assign n5091 = ~preset & n_n9348 & (ndn3_2 | ~n4949_1);
  assign n5092 = ~preset & n_n7136 & (~ndn3_39 | ndn3_40);
  assign n5093 = ~ndn3_2 & ~preset & psv26_6_6_ & n4949_1;
  assign n5094_1 = ~preset & n_n8051 & (ndn3_2 | ~n4949_1);
  assign n5095 = ~preset & n_n8850 & (ngfdn_3 | ~ndn3_46);
  assign n5096 = ndn3_46 & n_n9573 & ~preset & ~ngfdn_3;
  assign n5097 = n4950 & (n5975 | (n4975 & n7176));
  assign n5098 = n4856 & (n_n8561 ^ ~n4999_1);
  assign n5099_1 = ~preset & n_n8058 & (~ndn3_17 | ndn3_18);
  assign n5100 = ~ndn3_2 & ~preset & psv26_15_15_ & n4949_1;
  assign n5101 = ~preset & n_n8192 & (ndn3_2 | ~n4949_1);
  assign n5102 = ~preset & n_n7949 & (nsr3_38 | ndn3_38);
  assign n5103 = ~preset & n_n7792 & (ndn3_9 | ~ndn3_7);
  assign n5104_1 = ~ndn3_2 & ~preset & psv18_4_4_ & n4949_1;
  assign n5105 = ~preset & n_n9232 & (ndn3_2 | ~n4949_1);
  assign n5106 = ~ndn3_2 & ~preset & psv13_12_12_ & n4949_1;
  assign n5107 = ~preset & n_n7815 & (ndn3_2 | ~n4949_1);
  assign n5108 = ~ndn3_2 & ~preset & psv2_6_6_ & n4949_1;
  assign n5109_1 = ~preset & n_n7881 & (ndn3_2 | ~n4949_1);
  assign n5110 = ~ndn3_2 & ~preset & psv18_0_0_ & n4949_1;
  assign n5111 = ~preset & n_n8033 & (ndn3_2 | ~n4949_1);
  assign n5112 = ~preset & n_n9525 & (nsr3_14 | ndn3_14);
  assign n5113 = ~ndn3_2 & ~preset & psv2_0_0_ & n4949_1;
  assign n5114_1 = ~preset & n_n8770 & (ndn3_2 | ~n4949_1);
  assign n5115 = n4949_1 & ~ndn3_2 & pinp_6_6_ & ~preset;
  assign n5116 = ~preset & n_n7644 & (ndn3_2 | ~n4949_1);
  assign n5117 = ~preset & n_n8151 & (ndn3_19 | ~nen3_19);
  assign n5118 = ~preset & n4865 & (~n4976 ^ ~n4977);
  assign n5119_1 = ~preset & n_n8226 & (ndn3_17 | ~ndn3_16);
  assign n5120 = ~preset & n_n8841 & (ndn3_23 | nsr3_23);
  assign n5121 = ~preset & n_n8280 & (ndn3_19 | ~nen3_19);
  assign n5122 = ~preset & n4865 & (~n4985 ^ ~n4986);
  assign n5123 = ~preset & n_n7846 & (ndn3_23 | nsr3_23);
  assign n5124_1 = ~preset & n_n7678 & (ndn3_42 | ~ndn3_40);
  assign n5125 = n_n7862 & ndn3_40 & ~preset & ~ndn3_42;
  assign n5126 = ~preset & n_n7666 & (ndn3_27 | ~ndn3_26);
  assign n5127 = ~preset & n4859_1 & (~n4976 ^ ~n4977);
  assign n5128 = ~preset & n_n9520 & (~nen3_22 | ndn3_22);
  assign n5129_1 = ~ndn3_2 & ~preset & psv39_8_8_ & n4949_1;
  assign n5130 = ~preset & n_n7956 & (ndn3_2 | ~n4949_1);
  assign n5131 = ~preset & n_n7732 & (ndn3_30 | nsr3_30);
  assign n5132 = ~preset & n_n7859 & (ndn3_28 | ~nen3_28);
  assign n5133 = n4949_1 & ~ndn3_2 & pinp_12_12_ & ~preset;
  assign n5134_1 = ~preset & n_n8108 & (ndn3_2 | ~n4949_1);
  assign n5135 = ~preset & n_n9026 & (~nen3_22 | ndn3_22);
  assign n5136 = ~ndn3_22 & ~preset & nen3_22 & n_n7236;
  assign n5137 = ~ndn3_2 & ~preset & psv38_12_12_ & n4949_1;
  assign n5138 = ~preset & n_n8088 & (ndn3_2 | ~n4949_1);
  assign n5139_1 = ~ndn3_2 & ~preset & psv38_13_13_ & n4949_1;
  assign n5140 = ~preset & n_n9225 & (ndn3_2 | ~n4949_1);
  assign n5141 = ~preset & n_n8102 & (ndn3_42 | ~ndn3_40);
  assign n5142 = ndn3_40 & n_n9542 & ~preset & ~ndn3_42;
  assign n5143 = ~preset & n_n9347 & (ndn3_4 | ~ndn3_2);
  assign n5144_1 = ~preset & n_n7130 & (ngfdn_3 | ~ndn3_46);
  assign n5145 = ndn3_46 & n_n7527 & ~preset & ~ngfdn_3;
  assign n5146 = ~preset & n_n7444 & (ndn3_46 | ~ndn3_44);
  assign n5147 = ~preset & n_n9542 & (~ndn3_39 | ndn3_40);
  assign n5148 = n4846 & (n4997 ^ (n6083 | n6084_1));
  assign n5149_1 = ~preset & n_n8371 & (ndn3_42 | ~ndn3_40);
  assign n5150 = ndn3_40 & n_n9452 & ~preset & ~ndn3_42;
  assign n5151 = ~preset & n_n9455 & (~nen3_36 | ndn3_36);
  assign n5152 = ~preset & n_n9261 & (~nen3_36 | ndn3_36);
  assign n5153 = ~preset & n4876 & (~n4969_1 ^ ~n4970);
  assign n5154_1 = ~preset & n_n7022 & (ndn3_42 | ~ndn3_40);
  assign n5155 = ~ndn3_42 & ~preset & n_n8959 & ndn3_40;
  assign n5156 = ~preset & n_n8303 & (ndn3_42 | ~ndn3_40);
  assign n5157 = ~ndn3_42 & ~preset & n_n8957 & ndn3_40;
  assign n5158 = ~preset & n_n9593 & (ndn3_28 | ~nen3_28);
  assign n5159_1 = ~preset & n4892 & (~n4969_1 ^ ~n4970);
  assign n5160 = ~preset & n_n7435 & (~ndn3_42 | ndn3_44);
  assign n5161 = ~ndn3_44 & ~preset & ndn3_42 & n_n7927;
  assign n5162 = ~preset & n_n9313 & (ndn3_28 | ~nen3_28);
  assign n5163 = ~preset & n4892 & (~n4954_1 ^ ~n4955);
  assign n5164_1 = ~preset & n_n9522 & (ndn3_23 | nsr3_23);
  assign n5165 = ~preset & n_n9488 & (nsr3_35 | ndn3_35);
  assign n5166 = ~preset & n_n9237 & (~ndn3_42 | ndn3_44);
  assign n5167 = ~preset & n_n9239 & (~ndn3_42 | ndn3_44);
  assign n5168 = ~preset & n_n9452 & (~ndn3_39 | ndn3_40);
  assign n5169_1 = ~preset & n_n9498 & (ndn3_13 | nsr3_13);
  assign n5170 = ~preset & n_n8439 & (~ndn3_42 | ndn3_44);
  assign n5171 = ~ndn3_44 & ndn3_42 & ~preset & n_n7757;
  assign n5172 = ~preset & n_n8146 & (~ndn3_42 | ndn3_44);
  assign n5173 = ~ndn3_44 & ndn3_42 & ~preset & n_n8024;
  assign n5174_1 = ~preset & n_n9376 & (ngfdn_3 | ~ndn3_46);
  assign n5175 = ndn3_46 & n_n8436 & ~preset & ~ngfdn_3;
  assign n5176 = n4948 & (n5975 | (n4975 & n7176));
  assign n5177 = n4856 & n4947;
  assign n5178 = ~preset & n_n7843 & (~ngfdn_3 | ndn3_50);
  assign n5179_1 = ~ndn3_50 & ~preset & ngfdn_3 & n_n8256;
  assign n5180 = ~ndn3_2 & ~preset & psv18_8_8_ & n4949_1;
  assign n5181 = ~preset & n_n8966 & (ndn3_2 | ~n4949_1);
  assign n5182 = ~preset & n_n7674 & (ndn3_46 | ~ndn3_44);
  assign n5183 = n_n9237 & ndn3_44 & ~preset & ~ndn3_46;
  assign n5184_1 = ~preset & n_n8727 & (ndn3_17 | ~ndn3_16);
  assign n5185 = ~preset & n_n6910 & (ndn3_46 | ~ndn3_44);
  assign n5186 = n_n9239 & ndn3_44 & ~preset & ~ndn3_46;
  assign n5187 = ~preset & n_n9081 & (nsr3_38 | ndn3_38);
  assign n5188 = ~ndn3_2 & ~preset & psv26_10_10_ & n4949_1;
  assign n5189_1 = ~preset & n_n7688 & (ndn3_2 | ~n4949_1);
  assign n5190 = ~preset & n_n9338 & (ndn3_25 | ~ndn3_22);
  assign n5191 = ~preset & n_n9061 & (nsr3_38 | ndn3_38);
  assign n5192 = ~preset & n_n7686 & (~nen3_16 | ndn3_16);
  assign n5193 = ~preset & n4875 & (~n4976 ^ ~n4977);
  assign n5194_1 = ~ndn3_2 & ~preset & psv33_12_12_ & n4949_1;
  assign n5195 = ~preset & n_n8267 & (ndn3_2 | ~n4949_1);
  assign n5196 = ~ndn3_2 & ~preset & psv39_10_10_ & n4949_1;
  assign n5197 = ~preset & n_n8116 & (ndn3_2 | ~n4949_1);
  assign n5198 = ~preset & n_n8296 & (~ndn3_9 | ndn3_11);
  assign n5199_1 = ~preset & n4847 & (~n4971 ^ ~n4972);
  assign n5200 = ~preset & n_n8344 & (ndn3_13 | nsr3_13);
  assign n5201 = ~preset & n_n8326 & (ndn3_37 | nsr3_37);
  assign n5202 = n4949_1 & ~ndn3_2 & pinp_0_0_ & ~preset;
  assign n5203 = ~preset & n_n8011 & (ndn3_2 | ~n4949_1);
  assign n5204_1 = ~preset & n_n8583 & (ndn3_17 | ~ndn3_16);
  assign n5205 = n4946 & (n5975 | (n4975 & n7176));
  assign n5206 = n4856 & (n_n8993 ^ ~n5005);
  assign n5207 = n4944_1 & (n5975 | (n4975 & n7176));
  assign n5208 = n4856 & n4945;
  assign n5209_1 = ~preset & n_n8628 & (~ndn3_29 | ndn3_32);
  assign n5210 = ~preset & n4880 & (~n4976 ^ ~n4977);
  assign n5211 = ~ndn3_2 & ~preset & psv18_10_10_ & n4949_1;
  assign n5212 = ~preset & n_n8586 & (ndn3_2 | ~n4949_1);
  assign n5213 = ~preset & n_n9340 & (ndn3_23 | nsr3_23);
  assign n5214_1 = ~ndn3_2 & ~preset & psv18_12_12_ & n4949_1;
  assign n5215 = ~preset & n_n8408 & (ndn3_2 | ~n4949_1);
  assign n5216 = ~ndn3_2 & ~preset & psv26_7_7_ & n4949_1;
  assign n5217 = ~preset & n_n9603 & (ndn3_2 | ~n4949_1);
  assign n5218 = ~preset & n_n7682 & (nsr3_35 | ndn3_35);
  assign n5219_1 = ~ndn3_2 & ~preset & psv26_1_1_ & n4949_1;
  assign n5220 = ~preset & n_n9322 & (ndn3_2 | ~n4949_1);
  assign n5221 = ~ndn3_2 & ~preset & psv33_0_0_ & n4949_1;
  assign n5222 = ~preset & n_n7511 & (ndn3_2 | ~n4949_1);
  assign n5223 = ~preset & n_n7121 & (~ndn3_39 | ndn3_40);
  assign n5224_1 = ~ndn3_40 & n_n7626 & ~preset & ndn3_39;
  assign n5225 = ~preset & n_n8468 & (~ndn3_42 | ndn3_44);
  assign n5226 = n4861 & (n4997 ^ (n6083 | n6084_1));
  assign n5227 = n4942 & (n5975 | (n4975 & n7176));
  assign n5228 = n4856 & (~n_n9031 ^ (n_n8993 | n5005));
  assign n5229_1 = ~preset & n_n9424 & (~ndn3_39 | ndn3_40);
  assign n5230 = ~ndn3_40 & ~preset & ndn3_39 & n_n7346;
  assign n5231 = ~preset & n_n9404 & (ndn3_7 | ~ndn3_4);
  assign n5232 = ~preset & n_n9402 & (nsr3_13 | ndn3_15);
  assign n5233 = ~preset & n_n8361 & (~ndn3_39 | ndn3_40);
  assign n5234_1 = ~ndn3_40 & ndn3_39 & ~preset & n_n9611;
  assign n5235 = ~preset & n_n7366 & (~ndn3_39 | ndn3_40);
  assign n5236 = ~ndn3_40 & ndn3_39 & ~preset & n_n9613;
  assign n5237 = ~preset & n_n9344 & (nsr3_14 | ndn3_14);
  assign n5238 = ~preset & n_n7083 & (ndn3_46 | ~ndn3_44);
  assign n5239_1 = ~preset & n_n8188 & (~ndn3_42 | ndn3_44);
  assign n5240 = n4861 & (n5004_1 ^ (n6527 | n6528));
  assign n5241 = ~preset & n_n9178 & (nsr3_14 | ndn3_14);
  assign n5242 = ~preset & n_n8644 & (~ndn3_39 | ndn3_40);
  assign n5243 = ~ndn3_40 & ndn3_39 & ~preset & n_n8543;
  assign n5244_1 = ~preset & n_n8670 & (~ndn3_42 | ndn3_44);
  assign n5245 = ~ndn3_2 & ~preset & psv33_3_3_ & n4949_1;
  assign n5246 = ~preset & n_n9136 & (ndn3_2 | ~n4949_1);
  assign n5247 = ~preset & n_n9390 & (ndn3_34 | ~nen3_34);
  assign n5248 = ~preset & n_n8789 & (ndn3_4 | ~ndn3_2);
  assign n5249_1 = ~preset & n_n9046 & (ndn3_27 | ~ndn3_26);
  assign n5250 = ~preset & n4859_1 & (~n4954_1 ^ ~n4955);
  assign n5251 = ~preset & n_n8938 & (~ndn3_25 | ndn3_26);
  assign n5252 = ~preset & n4851 & (~n4969_1 ^ ~n4970);
  assign n5253 = ~preset & n_n7402 & (ndn3_46 | ~ndn3_44);
  assign n5254_1 = ~ndn3_46 & ~preset & n_n9635 & ndn3_44;
  assign n5255 = ~ndn3_2 & ~preset & psv26_13_13_ & n4949_1;
  assign n5256 = ~preset & n_n9067 & (ndn3_2 | ~n4949_1);
  assign n5257 = ~preset & n_n7715 & (~ndn3_42 | ndn3_44);
  assign n5258 = ~ndn3_44 & ndn3_42 & ~preset & n_n9486;
  assign n5259_1 = ~preset & n_n6980 & (~nen3_22 | ndn3_22);
  assign n5260 = ~ndn3_22 & nen3_22 & ~preset & n_n9273;
  assign n5261 = ~ndn3_2 & ~preset & psv38_6_6_ & n4949_1;
  assign n5262 = ~preset & n_n8779 & (ndn3_2 | ~n4949_1);
  assign n5263 = n4941 & (n5975 | (n4975 & n7176));
  assign n5264_1 = n4856 & n4940;
  assign n5265 = ~preset & n_n8729 & (ndn3_17 | ~ndn3_16);
  assign n5266 = ~preset & n4882 & (~n4971 ^ ~n4972);
  assign n5267 = ~preset & n_n8916 & (ndn3_46 | ~ndn3_44);
  assign n5268 = ndn3_44 & n_n8670 & ~preset & ~ndn3_46;
  assign n5269_1 = ~ndn3_2 & ~preset & psv2_4_4_ & n4949_1;
  assign n5270 = ~preset & n_n7827 & (ndn3_2 | ~n4949_1);
  assign n5271 = ~ndn3_2 & ~preset & psv13_10_10_ & n4949_1;
  assign n5272 = ~preset & n_n9119 & (ndn3_2 | ~n4949_1);
  assign n5273 = ~ndn3_2 & ~preset & psv2_2_2_ & n4949_1;
  assign n5274_1 = ~preset & n_n7744 & (ndn3_2 | ~n4949_1);
  assign n5275 = ~preset & n_n8909 & (nsr3_14 | ndn3_14);
  assign n5276 = ~ndn3_2 & ~preset & psv13_0_0_ & n4949_1;
  assign n5277 = ~preset & n_n8619 & (ndn3_2 | ~n4949_1);
  assign n5278 = ~preset & n_n8535 & (nsr3_14 | ndn3_14);
  assign n5279_1 = ~preset & n_n9255 & (~ndn3_19 | ndn3_21);
  assign n5280 = ~preset & n4885 & (~n4976 ^ ~n4977);
  assign n5281 = ~preset & n_n7969 & (nsr3_14 | ndn3_14);
  assign n5282 = ~preset & n_n9493 & (~nen3_22 | ndn3_22);
  assign n5283 = ~preset & n_n8657 & (nsr3_20 | ndn3_20);
  assign n5284_1 = ~preset & n_n8636 & (ndn3_37 | nsr3_37);
  assign n5285 = ~preset & n_n8477 & (ndn3_37 | nsr3_37);
  assign n5286 = ~ndn3_2 & ~preset & psv2_13_13_ & n4949_1;
  assign n5287 = ~preset & n_n7890 & (ndn3_2 | ~n4949_1);
  assign n5288 = n4939_1 & (n5975 | (n4975 & n7176));
  assign n5289_1 = n4856 & (~n_n8603 ^ ~n_n8798);
  assign n5290 = ~ndn3_2 & ~preset & psv38_10_10_ & n4949_1;
  assign n5291 = ~preset & n_n7665 & (ndn3_2 | ~n4949_1);
  assign n5292 = n7208 & n4856 & n5001;
  assign n5293 = ~n5001 & ~preset & n_n9353;
  assign n5294_1 = ~preset & n_n9139 & (ndn3_19 | ~nen3_19);
  assign n5295 = ~preset & n4865 & (~n4969_1 ^ ~n4970);
  assign n5296 = ~preset & n_n8839 & (ndn3_28 | ~nen3_28);
  assign n5297 = ~preset & n_n8185 & (~nen3_22 | ndn3_22);
  assign n5298 = ~ndn3_22 & n_n9304 & ~preset & nen3_22;
  assign n5299_1 = ~preset & n_n9155 & (~ndn3_39 | ndn3_40);
  assign n5300 = ~preset & n_n9508 & (ngfdn_3 | ~ndn3_46);
  assign n5301 = n1270 & (n4980 ^ (n6352 | n6353));
  assign n5302 = ~preset & n_n9126 & (~ndn3_29 | ndn3_32);
  assign n5303 = ~preset & n_n9629 & (ndn3_46 | ~ndn3_44);
  assign n5304_1 = n4853 & (n4997 ^ (n6083 | n6084_1));
  assign n5305 = ~preset & n_n9317 & (~nen3_16 | ndn3_16);
  assign n5306 = ~preset & n4875 & (~n4954_1 ^ ~n4955);
  assign n5307 = ~preset & n_n9600 & (nsr3_13 | ndn3_15);
  assign n5308 = ~preset & n4881 & (~n4969_1 ^ ~n4970);
  assign n5309_1 = n7207 & ((n4922 & n4935) | (n_n9537 & (n4922 | n4935)));
  assign n5310 = ~n_n8821 & n4857 & (~n4934_1 ^ ~n4937);
  assign n5311 = ~n4937 & ~n4934_1 & n_n8821 & n4856;
  assign n5312 = ~n5001 & ~preset & n_n8821;
  assign n5313 = ~preset & n_n7074 & (~ndn3_42 | ndn3_44);
  assign n5314_1 = ~ndn3_44 & ndn3_42 & ~preset & n_n9355;
  assign n5315 = ~preset & n_n8249 & (ndn3_42 | ~ndn3_40);
  assign n5316 = ~ndn3_2 & ~preset & psv26_4_4_ & n4949_1;
  assign n5317 = ~preset & n_n8617 & (ndn3_2 | ~n4949_1);
  assign n5318 = ~preset & n_n7069 & (~ngfdn_3 | ndn3_50);
  assign n5319_1 = ~ndn3_50 & n_n7324 & ~preset & ngfdn_3;
  assign n5320 = ~ndn3_2 & ~preset & psv33_1_1_ & n4949_1;
  assign n5321 = ~preset & n_n9053 & (ndn3_2 | ~n4949_1);
  assign n5322 = ~preset & n_n9129 & (ndn3_27 | ~ndn3_26);
  assign n5323 = ~preset & n_n9320 & (ndn3_13 | nsr3_13);
  assign n5324_1 = ~ndn3_2 & ~preset & psv13_15_15_ & n4949_1;
  assign n5325 = ~preset & n_n8502 & (ndn3_2 | ~n4949_1);
  assign n5326 = ~ndn3_2 & ~preset & psv18_6_6_ & n4949_1;
  assign n5327 = ~preset & n_n9230 & (ndn3_2 | ~n4949_1);
  assign n5328 = ~ndn3_2 & ~preset & psv38_4_4_ & n4949_1;
  assign n5329_1 = ~preset & n_n7600 & (ndn3_2 | ~n4949_1);
  assign n5330 = ~preset & n_n8221 & (nsr3_14 | ndn3_14);
  assign n5331 = ~preset & n_n9595 & (ndn3_25 | ~ndn3_22);
  assign n5332 = ~preset & n4889_1 & (~n4969_1 ^ ~n4970);
  assign n5333 = ~preset & n_n7642 & (~ndn3_9 | ndn3_11);
  assign n5334_1 = n4949_1 & ~ndn3_2 & pinp_8_8_ & ~preset;
  assign n5335 = ~preset & n_n7697 & (ndn3_2 | ~n4949_1);
  assign n5336 = ~preset & n_n7108 & (~ndn3_39 | ndn3_40);
  assign n5337 = ~ndn3_40 & ndn3_39 & ~preset & n_n8794;
  assign n5338 = ~preset & n_n7810 & (~nen3_16 | ndn3_16);
  assign n5339_1 = ~preset & n_n7781 & (ngfdn_3 | ~ndn3_46);
  assign n5340 = n1270 & (n4987 ^ (n6433 | n6434));
  assign n5341 = ~preset & n_n7606 & (ngfdn_3 | ~ndn3_46);
  assign n5342 = ~preset & n_n9460 & (~ndn3_19 | ndn3_21);
  assign n5343 = ~preset & n4885 & (~n4985 ^ ~n4986);
  assign n5344_1 = ~preset & n_n8473 & (ndn3_25 | ~ndn3_22);
  assign n5345 = ~preset & n_n8224 & (ndn3_29 | ~ndn3_28);
  assign n5346 = ~ndn3_2 & ~preset & psv39_2_2_ & n4949_1;
  assign n5347 = ~preset & n_n7837 & (ndn3_2 | ~n4949_1);
  assign n5348 = ~preset & n_n8581 & (~ndn3_25 | ndn3_26);
  assign n5349_1 = ~preset & n_n8213 & (~ndn3_19 | ndn3_21);
  assign n5350 = ~preset & n4885 & (~n4969_1 ^ ~n4970);
  assign n5351 = ~preset & n_n9092 & (ndn3_30 | nsr3_30);
  assign n5352 = ~preset & n_n8781 & (~nen3_22 | ndn3_22);
  assign n5353 = ~ndn3_22 & ~preset & nen3_22 & n_n9255;
  assign n5354_1 = ~preset & n_n7990 & (nsr3_35 | ndn3_35);
  assign n5355 = ~preset & n_n8470 & (~ndn3_42 | ndn3_44);
  assign n5356 = ~preset & n_n9394 & (ndn3_30 | nsr3_30);
  assign n5357 = ~preset & n_n9355 & (ndn3_42 | ~ndn3_40);
  assign n5358 = n4863 & (n4997 ^ (n6083 | n6084_1));
  assign n5359_1 = ~preset & n_n7739 & (~nen3_22 | ndn3_22);
  assign n5360 = n7202 & (n_n8930 | ~n4967 | ~n7089);
  assign n5361 = n7203 & n7089 & ~n_n8930 & n4967;
  assign n5362 = ~preset & n_n7728 & (~nen3_22 | ndn3_22);
  assign n5363 = ~preset & n_n8045 & (ndn3_42 | ~ndn3_40);
  assign n5364_1 = n_n7136 & ndn3_40 & ~preset & ~ndn3_42;
  assign n5365 = ~preset & n_n9128 & (~nen3_36 | ndn3_36);
  assign n5366 = ~preset & n_n9159 & (ndn3_28 | ~nen3_28);
  assign n5367 = ~preset & n_n9591 & (nsr3_35 | ndn3_35);
  assign n5368 = ~preset & n_n9393 & (nsr3_35 | ndn3_35);
  assign n5369_1 = ~preset & n_n8263 & (~ngfdn_3 | ndn3_50);
  assign n5370 = ~ndn3_50 & n_n8081 & ~preset & ngfdn_3;
  assign n5371 = ~preset & n_n7848 & (~ndn3_9 | ndn3_11);
  assign n5372 = ~preset & n4847 & (~n4985 ^ ~n4986);
  assign n5373 = ~preset & n_n7626 & (~nen3_39 | ndn3_39);
  assign n5374_1 = ~preset & n4854_1 & (~n4971 ^ ~n4972);
  assign n5375 = ~preset & n_n9421 & (ndn3_46 | ~ndn3_44);
  assign n5376 = ~ndn3_46 & ~preset & n_n7691 & ndn3_44;
  assign n5377 = ~preset & n_n7849 & (ndn3_9 | ~ndn3_7);
  assign n5378 = ~preset & n4852 & (~n4985 ^ ~n4986);
  assign n5379_1 = ~preset & n_n7873 & (nsr3_38 | ndn3_38);
  assign n5380 = ~ndn3_2 & ~preset & psv33_14_14_ & n4949_1;
  assign n5381 = ~preset & n_n7914 & (ndn3_2 | ~n4949_1);
  assign n5382 = ~preset & n_n7668 & (ndn3_9 | ~ndn3_7);
  assign n5383 = ~preset & n4852 & (~n4976 ^ ~n4977);
  assign n5384_1 = ~preset & n_n7925 & (ndn3_30 | nsr3_30);
  assign n5385 = ~preset & n_n8256 & (ngfdn_3 | ~ndn3_46);
  assign n5386 = ~preset & n_n7711 & (ndn3_23 | nsr3_23);
  assign n5387 = ~preset & n_n7971 & (ndn3_4 | ~ndn3_2);
  assign n5388 = ~preset & n_n8064 & (nsr3_20 | ndn3_20);
  assign n5389_1 = ~preset & n_n7932 & (~nen3_22 | ndn3_22);
  assign n5390 = ~preset & n_n8233 & (nsr3_13 | ndn3_15);
  assign n5391 = ~preset & n4881 & (~n4971 ^ ~n4972);
  assign n5392 = ~preset & n_n8003 & (ndn3_25 | ~ndn3_22);
  assign n5393 = n7201 & ((n4895 & n4921) | (n_n9416 & (n4895 | n4921)));
  assign n5394_1 = ~n_n9537 & n4857 & (~n4922 ^ ~n4935);
  assign n5395 = ~n4935 & ~n4922 & n_n9537 & n4856;
  assign n5396 = ~n5001 & ~preset & n_n9537;
  assign n5397 = n7200 & ((n4870 & n4871) | (n_n9638 & (n4870 | n4871)));
  assign n5398 = ~n_n9448 & n4857 & (~n4872 ^ ~n4933);
  assign n5399_1 = ~n4933 & ~n4872 & n_n9448 & n4856;
  assign n5400 = ~n5001 & ~preset & n_n9448;
  assign n5401 = ~preset & n_n9221 & (ndn3_46 | ~ndn3_44);
  assign n5402 = ~preset & n_n9104 & (~ndn3_39 | ndn3_40);
  assign n5403 = ~preset & n_n8277 & (~ndn3_29 | ndn3_32);
  assign n5404_1 = ~preset & n4880 & (~n4985 ^ ~n4986);
  assign n5405 = ~preset & n_n8743 & (ndn3_19 | ~nen3_19);
  assign n5406 = ~preset & n4865 & (~n4954_1 ^ ~n4955);
  assign n5407 = ~ndn3_2 & ~preset & psv33_2_2_ & n4949_1;
  assign n5408 = ~preset & n_n7554 & (ndn3_2 | ~n4949_1);
  assign n5409_1 = n7199 & ((n4914_1 & n4951) | (n_n8419 & (n4914_1 | n4951)));
  assign n5410 = ~n_n8449 & n4857 & (~n4931 ^ ~n4932);
  assign n5411 = ~n4932 & ~n4931 & n_n8449 & n4856;
  assign n5412 = ~n5001 & ~preset & n_n8449;
  assign n5413 = ~preset & n_n8384 & (~nen3_22 | ndn3_22);
  assign n5414_1 = ~ndn3_22 & ~preset & nen3_22 & n_n8464;
  assign n5415 = ~ndn3_2 & ~preset & psv38_3_3_ & n4949_1;
  assign n5416 = ~preset & n_n9212 & (ndn3_2 | ~n4949_1);
  assign n5417 = ~preset & n_n9050 & (~ndn3_9 | ndn3_11);
  assign n5418 = ~preset & n4847 & (~n4954_1 ^ ~n4955);
  assign n5419_1 = ~preset & n_n9570 & (ngfdn_3 | ~ndn3_46);
  assign n5420 = n1270 & (n5004_1 ^ (n6527 | n6528));
  assign n5421 = ~preset & n_n9028 & (ngfdn_3 | ~ndn3_46);
  assign n5422 = ~preset & n_n9626 & (ngfdn_3 | ~ndn3_46);
  assign n5423 = ~ndn3_2 & ~preset & psv39_7_7_ & n4949_1;
  assign n5424_1 = ~preset & n_n9605 & (ndn3_2 | ~n4949_1);
  assign n5425 = ~preset & n_n6968 & (nsr3_35 | ndn3_35);
  assign n5426 = ~preset & n_n7390 & (~ndn3_39 | ndn3_40);
  assign n5427 = ~ndn3_40 & ~preset & ndn3_39 & n_n7334;
  assign n5428 = ~ndn3_2 & ~preset & psv33_7_7_ & n4949_1;
  assign n5429_1 = ~preset & n_n9270 & (ndn3_2 | ~n4949_1);
  assign n5430 = ~preset & n_n7284 & (ndn3_46 | ~ndn3_44);
  assign n5431 = ~ndn3_46 & ~preset & n_n7898 & ndn3_44;
  assign n5432 = ~preset & n_n9403 & (ndn3_13 | nsr3_13);
  assign n5433 = ~preset & n_n9308 & (ndn3_34 | ~nen3_34);
  assign n5434_1 = ~preset & n4860 & (~n4954_1 ^ ~n4955);
  assign n5435 = ~preset & n_n8584 & (~ndn3_11 | ndn3_12);
  assign n5436 = ~ndn3_2 & ~preset & psv26_14_14_ & n4949_1;
  assign n5437 = ~preset & n_n7946 & (ndn3_2 | ~n4949_1);
  assign n5438 = ~preset & n_n7420 & (~ngfdn_3 | ndn3_50);
  assign n5439_1 = ~ndn3_50 & ngfdn_3 & ~preset & n_n7558;
  assign n5440 = ~ndn3_2 & ~preset & psv18_2_2_ & n4949_1;
  assign n5441 = ~preset & n_n7737 & (ndn3_2 | ~n4949_1);
  assign n5442 = ~ndn3_2 & ~preset & psv39_11_11_ & n4949_1;
  assign n5443 = ~preset & n_n8506 & (ndn3_2 | ~n4949_1);
  assign n5444_1 = ~preset & n_n7598 & (~ndn3_29 | ndn3_32);
  assign n5445 = ~preset & n4880 & (~n4971 ^ ~n4972);
  assign n5446 = ~preset & n_n8328 & (ndn3_37 | nsr3_37);
  assign n5447 = n4929_1 & (n5975 | (n4975 & n7176));
  assign n5448 = n4856 & n4928;
  assign n5449_1 = ~preset & n_n9205 & (~ndn3_25 | ndn3_26);
  assign n5450 = ~preset & n_n8004 & (~nen3_22 | ndn3_22);
  assign n5451 = n4866 & (n4997 ^ (n6083 | n6084_1));
  assign n5452 = ~preset & n_n8061 & (ndn3_42 | ~ndn3_40);
  assign n5453 = ~ndn3_42 & ~preset & n_n9104 & ndn3_40;
  assign n5454_1 = ~ndn3_2 & ~preset & psv39_6_6_ & n4949_1;
  assign n5455 = ~preset & n_n9121 & (ndn3_2 | ~n4949_1);
  assign n5456 = ~preset & n_n8436 & (ndn3_46 | ~ndn3_44);
  assign n5457 = n4853 & (n4987 ^ (n6433 | n6434));
  assign n5458 = ~preset & n_n9309 & (ndn3_42 | ~ndn3_40);
  assign n5459_1 = ~preset & n_n9259 & (~ndn3_42 | ndn3_44);
  assign n5460 = ~preset & n_n7476 & (~nsr1_2 | nlc1_2);
  assign n5461 = ~nlc1_2 & nsr1_2 & ~preset_0_0_ & ~preset;
  assign n5462 = ~ndn3_2 & ~preset & psv26_9_9_ & n4949_1;
  assign n5463 = ~preset & n_n7424 & (ndn3_2 | ~n4949_1);
  assign n5464_1 = ~ndn3_2 & ~preset & psv33_4_4_ & n4949_1;
  assign n5465 = ~preset & n_n7604 & (ndn3_2 | ~n4949_1);
  assign n5466 = ~preset & n_n7649 & (ndn3_27 | ~ndn3_26);
  assign n5467 = ~preset & n_n7976 & (ngfdn_3 | ~ndn3_46);
  assign n5468 = ndn3_46 & n_n8765 & ~preset & ~ngfdn_3;
  assign n5469_1 = ~preset & n_n8898 & (ndn3_34 | ~nen3_34);
  assign n5470 = ~preset & n4860 & (~n4971 ^ ~n4972);
  assign n5471 = ~preset & n_n8222 & (ndn3_34 | ~nen3_34);
  assign n5472 = ~preset & n_n7964 & (ndn3_46 | ~ndn3_44);
  assign n5473 = ~ndn3_46 & ~preset & n_n9041 & ndn3_44;
  assign n5474_1 = ~preset & n_n7706 & (~ndn3_42 | ndn3_44);
  assign n5475 = ~preset & n_n9318 & (~ndn3_11 | ndn3_12);
  assign n5476 = ~preset & n4849_1 & (~n4954_1 ^ ~n4955);
  assign n5477 = n4949_1 & ~ndn3_2 & pinp_7_7_ & ~preset;
  assign n5478 = ~preset & n_n9271 & (ndn3_2 | ~n4949_1);
  assign n5479_1 = ~preset & n_n9042 & (~ndn3_29 | ndn3_32);
  assign n5480 = ~preset & n4880 & (~n4954_1 ^ ~n4955);
  assign n5481 = n4926 & (n5975 | (n4975 & n7176));
  assign n5482 = n4856 & n4927;
  assign n5483 = n4925 & (n5975 | (n4975 & n7176));
  assign n5484_1 = n4856 & ((n_n8923 & (~n_n8603 | n_n8798)) | (n_n8603 & ~n_n8923 & ~n_n8798));
  assign n5485 = n_n9248 & (~n_n9247 | ~n4902) & n7198;
  assign n5486 = ~n4902 & n_n9247 & ~preset & n_n9248;
  assign n5487 = ~preset & n_n9252 & (~ndn3_19 | ndn3_21);
  assign n5488 = ~preset & n4885 & (~n4971 ^ ~n4972);
  assign n5489_1 = ~preset & n_n9576 & (~ndn3_39 | ndn3_40);
  assign n5490 = ~preset & n_n6920 & (ndn3_46 | ~ndn3_44);
  assign n5491 = ndn3_44 & n_n8470 & ~preset & ~ndn3_46;
  assign n5492 = ~ndn3_2 & ~preset & psv38_8_8_ & n4949_1;
  assign n5493 = ~preset & n_n7692 & (ndn3_2 | ~n4949_1);
  assign n5494_1 = ~ndn3_2 & ~preset & psv2_8_8_ & n4949_1;
  assign n5495 = ~preset & n_n9023 & (ndn3_2 | ~n4949_1);
  assign n5496 = ~preset & n_n9059 & (nsr3_38 | ndn3_38);
  assign n5497 = ~preset & n_n7809 & (~nen3_22 | ndn3_22);
  assign n5498 = n4866 & (n4980 ^ (n6352 | n6353));
  assign n5499_1 = ~preset & n_n8889 & (ndn3_28 | ~nen3_28);
  assign n5500 = ~preset & n4892 & (~n4976 ^ ~n4977);
  assign n5501 = ~preset & n_n8253 & (~nen3_36 | ndn3_36);
  assign n5502 = ~preset & n4876 & (~n4971 ^ ~n4972);
  assign n5503 = ~preset & n_n7845 & (ndn3_27 | ~ndn3_26);
  assign n5504_1 = ~preset & n4859_1 & (~n4985 ^ ~n4986);
  assign n5505 = ~preset & n_n8989 & (ndn3_42 | ~ndn3_40);
  assign n5506 = n4863 & (n4987 ^ (n6433 | n6434));
  assign n5507 = ~preset & n_n8223 & (~ndn3_29 | ndn3_32);
  assign n5508 = ~preset & n_n9171 & (~ndn3_42 | ndn3_44);
  assign n5509_1 = ~preset & n_n7879 & (ndn3_13 | nsr3_13);
  assign n5510 = ~preset & n_n9186 & (ndn3_13 | nsr3_13);
  assign n5511 = ~preset & n_n7885 & (nsr3_38 | ndn3_38);
  assign n5512 = ~preset & n_n7966 & (ndn3_37 | nsr3_37);
  assign n5513 = ~preset & n_n8081 & (ngfdn_3 | ~ndn3_46);
  assign n5514_1 = n1270 & (n4997 ^ (n6083 | n6084_1));
  assign n5515 = ~preset & n_n9219 & (ngfdn_3 | ~ndn3_46);
  assign n5516 = ~preset & n_n9043 & (ndn3_37 | nsr3_37);
  assign n5517 = n4923 & (n5975 | (n4975 & n7176));
  assign n5518 = n4856 & (n_n8933 ^ ~n5000);
  assign n5519_1 = ~preset & n_n8100 & (~ndn3_39 | ndn3_40);
  assign n5520 = ~ndn3_40 & ndn3_39 & ~preset & n_n8871;
  assign n5521 = ~preset & n_n9266 & (nsr3_14 | ndn3_14);
  assign n5522 = ~preset & n_n7429 & (ndn3_19 | ~nen3_19);
  assign n5523 = ~preset & n4865 & (~n4971 ^ ~n4972);
  assign n5524_1 = ~preset & n_n8791 & (ndn3_4 | ~ndn3_2);
  assign n5525 = ~preset & n4874_1 & (~n4971 ^ ~n4972);
  assign n5526 = ~preset & n_n7624 & (~nen3_39 | ndn3_39);
  assign n5527 = ~preset & n_n9535 & (~ndn3_42 | ndn3_44);
  assign n5528 = ~ndn3_44 & ndn3_42 & ~preset & n_n9309;
  assign n5529_1 = ~preset & n_n8396 & (ndn3_13 | nsr3_13);
  assign n5530 = ~preset & n_n7813 & (ndn3_7 | ~ndn3_4);
  assign n5531 = ~ndn3_2 & ~preset & psv38_0_0_ & n4949_1;
  assign n5532 = ~preset & n_n7509 & (ndn3_2 | ~n4949_1);
  assign n5533 = ~preset & n_n7980 & (ndn3_30 | nsr3_30);
  assign n5534_1 = ~preset & n_n7667 & (ndn3_23 | nsr3_23);
  assign n5535 = ~preset & n_n7761 & (nsr3_20 | ndn3_20);
  assign n5536 = ~preset & n_n7683 & (ndn3_25 | ~ndn3_22);
  assign n5537 = ~preset & n4889_1 & (~n4976 ^ ~n4977);
  assign n5538 = ~preset & n_n8177 & (ndn3_29 | ~ndn3_28);
  assign n5539_1 = ~preset & n4869_1 & (~n4976 ^ ~n4977);
  assign n5540 = ~preset & n_n7793 & (ndn3_4 | ~ndn3_2);
  assign n5541 = ~ndn3_2 & ~preset & psv2_12_12_ & n4949_1;
  assign n5542 = ~preset & n_n7817 & (ndn3_2 | ~n4949_1);
  assign n5543 = ~preset & n_n7225 & (nsr3_20 | ndn3_20);
  assign n5544_1 = ~preset & n_n7808 & (ndn3_30 | nsr3_30);
  assign n5545 = ~preset & n_n6963 & (ndn3_42 | ~ndn3_40);
  assign n5546 = ~ndn3_42 & ~preset & n_n9155 & ndn3_40;
  assign n5547 = ~preset & n_n7392 & (~nen3_22 | ndn3_22);
  assign n5548 = ~ndn3_22 & ~preset & nen3_22 & n_n9586;
  assign n5549_1 = ~ndn3_2 & ~preset & psv33_8_8_ & n4949_1;
  assign n5550 = ~preset & n_n9302 & (ndn3_2 | ~n4949_1);
  assign n5551 = ~preset & n_n9458 & (ndn3_34 | ~nen3_34);
  assign n5552 = ~preset & n_n8801 & (~ndn3_42 | ndn3_44);
  assign n5553 = ~ndn3_44 & ndn3_42 & ~preset & n_n8247;
  assign n5554_1 = ~ndn3_2 & ~preset & psv18_3_3_ & n4949_1;
  assign n5555 = ~preset & n_n9396 & (ndn3_2 | ~n4949_1);
  assign n5556 = ~preset & n_n7231 & (~nen3_22 | ndn3_22);
  assign n5557 = ~ndn3_22 & ~preset & nen3_22 & n_n8093;
  assign n5558 = ~preset & n_n9312 & (ndn3_30 | nsr3_30);
  assign n5559_1 = ~preset & n_n8856 & (~nen3_22 | ndn3_22);
  assign n5560 = n4866 & (n5004_1 ^ (n6527 | n6528));
  assign n5561 = ~n5975 & n7196 & (~n4975 | ~n7176);
  assign n5562 = ~n6866 & ~n6865 & n_n8603 & ~n4856;
  assign n5563 = n7192 & ((n4893 & n4894_1) | (n_n9434 & (n4893 | n4894_1)));
  assign n5564_1 = ~n_n9416 & n4857 & (~n4895 ^ ~n4921);
  assign n5565 = ~n4921 & ~n4895 & n_n9416 & n4856;
  assign n5566 = ~n5001 & ~preset & n_n9416;
  assign n5567 = ~ndn3_2 & ~preset & psv39_1_1_ & n4949_1;
  assign n5568 = ~preset & n_n9324 & (ndn3_2 | ~n4949_1);
  assign n5569_1 = ~ndn3_2 & ~preset & psv33_5_5_ & n4949_1;
  assign n5570 = ~preset & n_n9182 & (ndn3_2 | ~n4949_1);
  assign n5571 = ~preset & n_n9278 & (~ngfdn_3 | ndn3_50);
  assign n5572 = ~ndn3_50 & ~preset & ngfdn_3 & n_n7781;
  assign n5573 = ~preset & n_n8014 & (ndn3_9 | ~ndn3_7);
  assign n5574_1 = ~preset & n_n8961 & (ndn3_9 | ~ndn3_7);
  assign n5575 = ~ndn3_2 & ~preset & psv13_6_6_ & n4949_1;
  assign n5576 = ~preset & n_n7880 & (ndn3_2 | ~n4949_1);
  assign n5577 = ~ndn3_2 & ~preset & psv13_11_11_ & n4949_1;
  assign n5578 = ~preset & n_n7766 & (ndn3_2 | ~n4949_1);
  assign n5579_1 = ~preset & n_n7687 & (nsr3_13 | ndn3_15);
  assign n5580 = ~preset & n4881 & (~n4976 ^ ~n4977);
  assign n5581 = ~preset & n_n7685 & (nsr3_20 | ndn3_20);
  assign n5582 = ~preset & n_n8281 & (ndn3_17 | ~ndn3_16);
  assign n5583 = ~preset & n4882 & (~n4985 ^ ~n4986);
  assign n5584_1 = n4949_1 & ~ndn3_2 & pinp_2_2_ & ~preset;
  assign n5585 = ~preset & n_n8009 & (ndn3_2 | ~n4949_1);
  assign n5586 = ~preset & n_n7825 & (ndn3_7 | ~ndn3_4);
  assign n5587 = ~preset & n4879_1 & (~n4971 ^ ~n4972);
  assign n5588 = ~preset & n_n7878 & (nsr3_13 | ndn3_15);
  assign n5589_1 = ~preset & n_n7395 & (ndn3_42 | ~ndn3_40);
  assign n5590 = n_n8206 & ndn3_40 & ~preset & ~ndn3_42;
  assign n5591 = ~preset & n_n9327 & (ndn3_28 | ~nen3_28);
  assign n5592 = ~preset & n_n9176 & (ndn3_23 | nsr3_23);
  assign n5593 = ~preset & n_n7756 & (~ndn3_19 | ndn3_21);
  assign n5594_1 = ~preset & n_n8464 & (~ndn3_19 | ndn3_21);
  assign n5595 = ~preset & n_n7734 & (nsr3_35 | ndn3_35);
  assign n5596 = ~ndn3_2 & ~preset & psv26_5_5_ & n4949_1;
  assign n5597 = ~preset & n_n9500 & (ndn3_2 | ~n4949_1);
  assign n5598 = ~preset & n_n7650 & (nsr3_35 | ndn3_35);
  assign n5599_1 = ~preset & n_n7807 & (nsr3_35 | ndn3_35);
  assign n5600 = ~preset & n_n8794 & (~nen3_39 | ndn3_39);
  assign n5601 = ~preset & n_n7360 & (~nen3_22 | ndn3_22);
  assign n5602 = ~ndn3_22 & ~preset & nen3_22 & n_n7756;
  assign n5603 = ~preset & n_n8984 & (~ndn3_11 | ndn3_12);
  assign n5604_1 = ~preset & n_n9599 & (~ndn3_11 | ndn3_12);
  assign n5605 = ~preset & n4849_1 & (~n4969_1 ^ ~n4970);
  assign n5606 = ~ndn3_2 & ~preset & psv13_9_9_ & n4949_1;
  assign n5607 = ~preset & n_n7866 & (ndn3_2 | ~n4949_1);
  assign n5608 = ~preset & n_n8486 & (~ngfdn_3 | ndn3_50);
  assign n5609_1 = ~ndn3_50 & ~preset & ngfdn_3 & n_n9626;
  assign n5610 = ~ndn3_2 & ~preset & psv18_1_1_ & n4949_1;
  assign n5611 = ~preset & n_n9314 & (ndn3_2 | ~n4949_1);
  assign n5612 = ~preset & n_n8073 & (~ndn3_39 | ndn3_40);
  assign n5613 = ~ndn3_40 & n_n7624 & ~preset & ndn3_39;
  assign n5614_1 = ~preset & n_n7896 & (ndn3_46 | ~ndn3_44);
  assign n5615 = n4949_1 & ~ndn3_2 & pinp_9_9_ & ~preset;
  assign n5616 = ~preset & n_n9349 & (ndn3_2 | ~n4949_1);
  assign n5617 = ~ndn3_2 & ~preset & psv13_1_1_ & n4949_1;
  assign n5618 = ~preset & n_n9323 & (ndn3_2 | ~n4949_1);
  assign n5619_1 = ~ndn3_2 & ~preset & pinp_5_5_ & n4949_1;
  assign n5620 = ~preset & n_n9183 & (ndn3_2 | ~n4949_1);
  assign n5621 = ~preset & n_n8854 & (~nen3_22 | ndn3_22);
  assign n5622 = n4949_1 & ~ndn3_2 & pinp_3_3_ & ~preset;
  assign n5623 = ~preset & n_n9137 & (ndn3_2 | ~n4949_1);
  assign n5624_1 = ~preset & n_n9319 & (nsr3_13 | ndn3_15);
  assign n5625 = ~preset & n4881 & (~n4954_1 ^ ~n4955);
  assign n5626 = n7187 & ((n4912 & n4938) | (n_n9353 & (n4912 | n4938)));
  assign n5627 = ~preset & n_n9395 & (ndn3_28 | ~nen3_28);
  assign n5628 = ~preset & n_n7923 & (~ngfdn_3 | ndn3_50);
  assign n5629_1 = ~ndn3_50 & ngfdn_3 & ~preset & n_n7779;
  assign n5630 = ~preset & n_n8833 & (ndn3_13 | nsr3_13);
  assign n5631 = ~preset & n_n8276 & (~ndn3_9 | ndn3_11);
  assign n5632 = ~preset & n4847 & (~n4976 ^ ~n4977);
  assign n5633 = ~preset & n_n7514 & (ndn3_46 | ~ndn3_44);
  assign n5634_1 = ndn3_44 & n_n8188 & ~preset & ~ndn3_46;
  assign n5635 = ~ndn3_2 & ~preset & psv33_15_15_ & n4949_1;
  assign n5636 = ~preset & n_n8456 & (ndn3_2 | ~n4949_1);
  assign n5637 = ~ndn3_2 & ~preset & psv39_13_13_ & n4949_1;
  assign n5638 = ~preset & n_n8504 & (ndn3_2 | ~n4949_1);
  assign n5639_1 = ~preset & n_n7950 & (ndn3_30 | nsr3_30);
  assign n5640 = ~preset & n_n9315 & (ndn3_25 | ~ndn3_22);
  assign n5641 = ~preset & n4889_1 & (~n4954_1 ^ ~n4955);
  assign n5642 = ~preset & n_n8402 & (~ndn3_17 | ndn3_18);
  assign n5643 = ~preset & n_n7684 & (~nen3_22 | ndn3_22);
  assign n5644_1 = ~preset & n_n8552 & (~nen3_36 | ndn3_36);
  assign n5645 = ~ndn3_2 & ~preset & psv39_4_4_ & n4949_1;
  assign n5646 = ~preset & n_n7835 & (ndn3_2 | ~n4949_1);
  assign n5647 = ~ndn3_2 & ~preset & psv2_10_10_ & n4949_1;
  assign n5648 = ~preset & n_n7689 & (ndn3_2 | ~n4949_1);
  assign n5649_1 = ~preset & n_n9494 & (nsr3_20 | ndn3_20);
  assign n5650 = ~preset & n_n8982 & (ndn3_19 | ~nen3_19);
  assign n5651 = ~preset & n_n8095 & (nsr3_35 | ndn3_35);
  assign n5652 = ~preset & n_n8900 & (ndn3_30 | nsr3_30);
  assign n5653 = ~preset & n_n8210 & (nsr3_14 | ndn3_14);
  assign n5654_1 = ~preset & n_n8626 & (ndn3_34 | ~nen3_34);
  assign n5655 = ~preset & n4860 & (~n4985 ^ ~n4986);
  assign n5656 = ~preset & n_n7988 & (nsr3_35 | ndn3_35);
  assign n5657 = ~preset & n_n8906 & (~nen3_39 | ndn3_39);
  assign n5658 = ~preset & n4854_1 & (~n4969_1 ^ ~n4970);
  assign n5659_1 = ~preset & n_n9268 & (ndn3_9 | ~ndn3_7);
  assign n5660 = ~preset & n4852 & (~n4969_1 ^ ~n4970);
  assign n5661 = ~preset & n_n8983 & (ndn3_17 | ~ndn3_16);
  assign n5662 = ~preset & n_n7256 & (ndn3_46 | ~ndn3_44);
  assign n5663 = ~ndn3_46 & ~preset & n_n9171 & ndn3_44;
  assign n5664_1 = ~preset & n_n8939 & (ndn3_17 | ~ndn3_16);
  assign n5665 = ~preset & n4882 & (~n4969_1 ^ ~n4970);
  assign n5666 = ~ndn3_2 & ~preset & psv2_9_9_ & n4949_1;
  assign n5667 = ~preset & n_n8739 & (ndn3_2 | ~n4949_1);
  assign n5668 = ~preset & n_n9366 & (~ndn3_39 | ndn3_40);
  assign n5669_1 = ~ndn3_40 & n_n7464 & ~preset & ndn3_39;
  assign n5670 = ~preset & n_n9310 & (nsr3_38 | ndn3_38);
  assign n5671 = ~preset & n_n7570 & (ndn3_46 | ~ndn3_44);
  assign n5672 = n4853 & (n4980 ^ (n6352 | n6353));
  assign n5673 = ~preset & n_n9470 & (~ndn3_29 | ndn3_32);
  assign n5674_1 = ~preset & n4880 & (~n4969_1 ^ ~n4970);
  assign n5675 = ~preset & n_n9623 & (ndn3_42 | ~ndn3_40);
  assign n5676 = ~preset & n_n9609 & (~ndn3_39 | ndn3_40);
  assign n5677 = ~ndn3_2 & ~preset & psv2_1_1_ & n4949_1;
  assign n5678 = ~preset & n_n9325 & (ndn3_2 | ~n4949_1);
  assign n5679_1 = ~preset & n_n9342 & (~nen3_16 | ndn3_16);
  assign n5680 = n4949_1 & ~ndn3_2 & pinp_1_1_ & ~preset;
  assign n5681 = ~preset & n_n9054 & (ndn3_2 | ~n4949_1);
  assign n5682 = ~preset & n_n7822 & (~nen3_22 | ndn3_22);
  assign n5683 = ~ndn3_2 & ~preset & psv39_5_5_ & n4949_1;
  assign n5684_1 = ~preset & n_n9502 & (ndn3_2 | ~n4949_1);
  assign n5685 = ~preset & n_n8741 & (ndn3_29 | ~ndn3_28);
  assign n5686 = ~preset & n4869_1 & (~n4954_1 ^ ~n4955);
  assign n5687 = ~preset & n_n9371 & (~ndn3_39 | ndn3_40);
  assign n5688 = ~ndn3_40 & ndn3_39 & ~preset & n_n8611;
  assign n5689_1 = ~preset & n_n8980 & (ndn3_34 | ~nen3_34);
  assign n5690 = ~ndn3_2 & ~preset & psv26_2_2_ & n4949_1;
  assign n5691 = ~preset & n_n7743 & (ndn3_2 | ~n4949_1);
  assign n5692 = ~preset & n_n9429 & (~ngfdn_3 | ndn3_50);
  assign n5693 = ~ndn3_50 & n_n7217 & ~preset & ngfdn_3;
  assign n5694_1 = ~preset & n_n6961 & (~ndn3_42 | ndn3_44);
  assign n5695 = ~ndn3_44 & ndn3_42 & ~preset & n_n8989;
  assign n5696 = ~preset & n_n8809 & (~ndn3_25 | ndn3_26);
  assign n5697 = ~preset & n_n8340 & (ndn3_46 | ~ndn3_44);
  assign n5698 = ndn3_44 & n_n8468 & ~preset & ~ndn3_46;
  assign n5699_1 = ~ndn3_2 & ~preset & psv39_14_14_ & n4949_1;
  assign n5700 = ~preset & n_n7936 & (ndn3_2 | ~n4949_1);
  assign n5701 = ~preset & n_n8430 & (~ndn3_39 | ndn3_40);
  assign n5702 = ~ndn3_40 & ndn3_39 & ~preset & n_n9106;
  assign n5703 = ~preset & n_n9596 & (~nen3_22 | ndn3_22);
  assign n5704_1 = ~preset & n_n7876 & (~nen3_16 | ndn3_16);
  assign n5705 = n4917 & (n5975 | (n4975 & n7176));
  assign n5706 = n4856 & (~n_n8911 ^ (n_n8933 | n5000));
  assign n5707 = ~preset & n_n7887 & (ndn3_25 | ~ndn3_22);
  assign n5708 = ~preset & n4889_1 & (~n4985 ^ ~n4986);
  assign n5709_1 = ~preset & n_n8760 & (ndn3_4 | ~ndn3_2);
  assign n5710 = ~preset & n4874_1 & (~n4976 ^ ~n4977);
  assign n5711 = ~preset & n_n9264 & (ndn3_23 | nsr3_23);
  assign n5712 = ~ndn3_2 & ~preset & psv39_0_0_ & n4949_1;
  assign n5713 = ~preset & n_n7657 & (ndn3_2 | ~n4949_1);
  assign n5714_1 = ~preset & n_n9102 & (~ndn3_39 | ndn3_40);
  assign n5715 = n4846 & (n4987 ^ (n6433 | n6434));
  assign n5716 = ~preset & n_n9316 & (nsr3_20 | ndn3_20);
  assign n5717 = ~preset & n_n7929 & (ndn3_30 | nsr3_30);
  assign n5718 = ~preset & n_n7962 & (~ndn3_39 | ndn3_40);
  assign n5719_1 = n4846 & (n4996 ^ (n6545 | n6546));
  assign n5720 = ~ndn3_2 & ~preset & psv18_14_14_ & n4949_1;
  assign n5721 = ~preset & n_n7930 & (ndn3_2 | ~n4949_1);
  assign n5722 = ~preset & n_n8864 & (~ndn3_29 | ndn3_32);
  assign n5723 = n7186 & ((n4872 & n4933) | (n_n9448 & (n4872 | n4933)));
  assign n5724_1 = ~n_n8354 & n4857 & (~n4915 ^ ~n4916);
  assign n5725 = ~n4916 & ~n4915 & n_n8354 & n4856;
  assign n5726 = ~n5001 & ~preset & n_n8354;
  assign n5727 = ~preset & n_n7789 & (~nen3_36 | ndn3_36);
  assign n5728 = ~preset & n_n8543 & (~nen3_39 | ndn3_39);
  assign n5729_1 = ~preset & n4854_1 & (~n4976 ^ ~n4977);
  assign n5730 = ~preset & n_n8480 & (ndn3_37 | nsr3_37);
  assign n5731 = ~preset & n_n9487 & (nsr3_38 | ndn3_38);
  assign n5732 = ~preset & n_n7967 & (~nen3_36 | ndn3_36);
  assign n5733 = ~preset & n_n8744 & (ndn3_17 | ~ndn3_16);
  assign n5734_1 = ~preset & n4882 & (~n4954_1 ^ ~n4955);
  assign n5735 = ~preset & n_n8022 & (ndn3_42 | ~ndn3_40);
  assign n5736 = n4863 & (n4980 ^ (n6352 | n6353));
  assign n5737 = ~preset & n_n9592 & (ndn3_30 | nsr3_30);
  assign n5738 = ~preset & n_n8808 & (ndn3_29 | ~ndn3_28);
  assign n5739_1 = ~preset & n_n9044 & (~nen3_36 | ndn3_36);
  assign n5740 = ~preset & n4876 & (~n4954_1 ^ ~n4955);
  assign n5741 = ~ndn3_2 & ~preset & psv39_3_3_ & n4949_1;
  assign n5742 = ~preset & n_n9407 & (ndn3_2 | ~n4949_1);
  assign n5743 = ~preset & n_n9132 & (nsr3_14 | ndn3_14);
  assign n5744_1 = ~preset & n_n9337 & (ndn3_27 | ~ndn3_26);
  assign n5745 = ~preset & n_n8589 & (ngfdn_3 | ~ndn3_46);
  assign n5746 = n_n9221 & ndn3_46 & ~preset & ~ngfdn_3;
  assign n5747 = ~preset & n_n7603 & (~ndn3_17 | ndn3_18);
  assign n5748 = ~preset & n4877 & (~n4971 ^ ~n4972);
  assign n5749_1 = n4908 & (n5975 | (n4975 & n7176));
  assign n5750 = n4856 & ((~n_n8913 & ~n_n8964 & ~n4968) | (n_n8964 & (n_n8913 | n4968)));
  assign n5751 = ~ndn3_2 & ~preset & psv38_2_2_ & n4949_1;
  assign n5752 = ~preset & n_n8638 & (ndn3_2 | ~n4949_1);
  assign n5753 = ~preset & n_n7017 & (~nen3_22 | ndn3_22);
  assign n5754_1 = ~ndn3_22 & ~preset & nen3_22 & n_n9087;
  assign n5755 = ~preset & n_n9397 & (ndn3_25 | ~ndn3_22);
  assign n5756 = ~preset & n_n8519 & (nsr3_13 | ndn3_15);
  assign n5757 = ~preset & n_n9368 & (~nen3_22 | ndn3_22);
  assign n5758 = ~preset & n_n8750 & (ndn3_42 | ~ndn3_40);
  assign n5759_1 = ~ndn3_42 & ~preset & n_n7962 & ndn3_40;
  assign n5760 = ~preset & n_n7968 & (ndn3_23 | nsr3_23);
  assign n5761 = n4949_1 & ~ndn3_2 & pinp_14_14_ & ~preset;
  assign n5762 = ~preset & n_n8000 & (ndn3_2 | ~n4949_1);
  assign n5763 = n4949_1 & ~ndn3_2 & pinp_11_11_ & ~preset;
  assign n5764_1 = ~preset & n_n8986 & (ndn3_2 | ~n4949_1);
  assign n5765 = ~preset & n_n7820 & (ndn3_28 | ~nen3_28);
  assign n5766 = ~preset & n4892 & (~n4971 ^ ~n4972);
  assign n5767 = ~preset & n_n9333 & (~ndn3_42 | ndn3_44);
  assign n5768 = n4861 & (n4987 ^ (n6433 | n6434));
  assign n5769_1 = ~preset & n_n9047 & (ndn3_23 | nsr3_23);
  assign n5770 = ~preset & n_n8810 & (ndn3_19 | ~nen3_19);
  assign n5771 = ~preset & n_n8381 & (nsr3_14 | ndn3_14);
  assign n5772 = ~preset & n_n9041 & (~ndn3_42 | ndn3_44);
  assign n5773 = ~preset & n_n8093 & (~ndn3_19 | ndn3_21);
  assign n5774_1 = ~preset & n4885 & (~n4954_1 ^ ~n4955);
  assign n5775 = ~preset & n_n7102 & (ndn3_42 | ~ndn3_40);
  assign n5776 = ~ndn3_42 & ~preset & n_n9609 & ndn3_40;
  assign n5777 = n7180 & ((n4931 & n4932) | (n_n8449 & (n4931 | n4932)));
  assign n5778 = ~n_n8549 & n4857 & (~n4905 ^ ~n4906);
  assign n5779_1 = ~n4906 & ~n4905 & n_n8549 & n4856;
  assign n5780 = ~n5001 & ~preset & n_n8549;
  assign n5781 = ~preset & n_n7681 & (nsr3_38 | ndn3_38);
  assign n5782 = ~preset & n_n9346 & (ndn3_9 | ~ndn3_7);
  assign n5783 = ~ndn3_2 & ~preset & psv38_9_9_ & n4949_1;
  assign n5784_1 = ~preset & n_n9336 & (ndn3_2 | ~n4949_1);
  assign n5785 = ~preset & n_n9134 & (ndn3_9 | ~ndn3_7);
  assign n5786 = ~ndn3_2 & ~preset & psv18_5_5_ & n4949_1;
  assign n5787 = ~preset & n_n9491 & (ndn3_2 | ~n4949_1);
  assign n5788 = ~preset & n_n9334 & (~ndn3_29 | ndn3_32);
  assign n5789_1 = ~ndn3_2 & ~preset & psv38_1_1_ & n4949_1;
  assign n5790 = ~preset & n_n9045 & (ndn3_2 | ~n4949_1);
  assign n5791 = ~preset & n_n9282 & (ngfdn_3 | ~ndn3_46);
  assign n5792 = ~preset & n_n8697 & (ndn3_23 | nsr3_23);
  assign n5793 = ~preset & n_n7875 & (nsr3_20 | ndn3_20);
  assign n5794_1 = ~preset & n_n9036 & (ndn3_42 | ~ndn3_40);
  assign n5795 = ~preset & n_n7527 & (ndn3_46 | ~ndn3_44);
  assign n5796 = ~preset & n_n7454 & (ndn3_19 | ~nen3_19);
  assign n5797 = ~preset & n_n8369 & (~ngfdn_3 | ndn3_50);
  assign n5798 = ~ndn3_50 & ~preset & ngfdn_3 & n_n9508;
  assign n5799_1 = ~preset & n_n9263 & (ndn3_27 | ~ndn3_26);
  assign n5800 = ~preset & n4859_1 & (~n4969_1 ^ ~n4970);
  assign n5801 = ~preset & n_n8153 & (~ndn3_11 | ndn3_12);
  assign n5802 = ~preset & n4849_1 & (~n4976 ^ ~n4977);
  assign n5803 = ~preset & n_n9004 & (ngfdn_3 | ~ndn3_46);
  assign n5804_1 = ndn3_46 & n_n8951 & ~preset & ~ngfdn_3;
  assign n5805 = ~preset & n_n8049 & (~ndn3_42 | ndn3_44);
  assign n5806 = ~ndn3_44 & ndn3_42 & ~preset & n_n9589;
  assign n5807 = ~preset & n_n9148 & (~ngfdn_3 | ndn3_50);
  assign n5808 = ~ndn3_50 & ~preset & ngfdn_3 & n_n7606;
  assign n5809_1 = ~preset & n_n7498 & (~ndn3_42 | ndn3_44);
  assign n5810 = ~ndn3_44 & ndn3_42 & ~preset & n_n9391;
  assign n5811 = ~preset & n_n7824 & (~ndn3_11 | ndn3_12);
  assign n5812 = ~preset & n4849_1 & (~n4971 ^ ~n4972);
  assign n5813 = ~preset & n_n7777 & (~nen3_22 | ndn3_22);
  assign n5814_1 = ~ndn3_22 & ~preset & nen3_22 & n_n9100;
  assign n5815 = ~ndn3_2 & ~preset & psv13_4_4_ & n4949_1;
  assign n5816 = ~preset & n_n7826 & (ndn3_2 | ~n4949_1);
  assign n5817 = ~preset & n_n8777 & (~ndn3_39 | ndn3_40);
  assign n5818 = ~ndn3_40 & ~preset & ndn3_39 & n_n8858;
  assign n5819_1 = ~ndn3_2 & ~preset & psv33_10_10_ & n4949_1;
  assign n5820 = ~preset & n_n9300 & (ndn3_2 | ~n4949_1);
  assign n5821 = ~preset & n_n7847 & (~ndn3_17 | ndn3_18);
  assign n5822 = ~preset & n4877 & (~n4985 ^ ~n4986);
  assign n5823 = ~preset & n_n7760 & (~nen3_22 | ndn3_22);
  assign n5824_1 = ~preset & n_n8466 & (ngfdn_3 | ~ndn3_46);
  assign n5825 = ~preset & n_n7911 & (ndn3_23 | nsr3_23);
  assign n5826 = ~preset & n_n8582 & (ndn3_19 | ~nen3_19);
  assign n5827 = ~preset & n_n7790 & (ndn3_27 | ~ndn3_26);
  assign n5828 = ~preset & n_n8279 & (~ndn3_25 | ndn3_26);
  assign n5829_1 = ~preset & n4851 & (~n4985 ^ ~n4986);
  assign n5830 = ~ndn3_2 & ~preset & psv2_11_11_ & n4949_1;
  assign n5831 = ~preset & n_n9387 & (ndn3_2 | ~n4949_1);
  assign n5832 = ~preset & n_n9589 & (ndn3_42 | ~ndn3_40);
  assign n5833 = ~preset & n_n8951 & (ndn3_46 | ~ndn3_44);
  assign n5834_1 = ~preset & n_n9573 & (ndn3_46 | ~ndn3_44);
  assign n5835 = n4853 & (n4996 ^ (n6545 | n6546));
  assign n5836 = ~preset & n_n8659 & (nsr3_14 | ndn3_14);
  assign n5837 = ~preset & n_n8681 & (ndn3_42 | ~ndn3_40);
  assign n5838 = ~ndn3_42 & ~preset & n_n8996 & ndn3_40;
  assign n5839_1 = ~preset & n_n8042 & (nsr3_14 | ndn3_14);
  assign n5840 = ~preset & n_n8941 & (ndn3_29 | ~ndn3_28);
  assign n5841 = ~ndn3_2 & ~preset & psv33_6_6_ & n4949_1;
  assign n5842 = ~preset & n_n7643 & (ndn3_2 | ~n4949_1);
  assign n5843 = ~preset & n_n7775 & (ngfdn_3 | ~ndn3_46);
  assign n5844_1 = n_n7083 & ndn3_46 & ~preset & ~ngfdn_3;
  assign n5845 = ~preset & n_n9096 & (ngfdn_3 | ~ndn3_46);
  assign n5846 = ndn3_46 & n_n8258 & ~preset & ~ngfdn_3;
  assign n5847 = ~preset & n_n9189 & (ndn3_13 | nsr3_13);
  assign n5848 = ~preset & n_n9341 & (~ndn3_17 | ndn3_18);
  assign n5849_1 = ~preset & n_n8260 & (ndn3_13 | nsr3_13);
  assign n5850 = ~preset & n_n7918 & (nsr3_38 | ndn3_38);
  assign n5851 = ~preset & n_n8996 & (~ndn3_39 | ndn3_40);
  assign n5852 = ~preset & n_n7806 & (nsr3_38 | ndn3_38);
  assign n5853 = ~preset & n_n8024 & (ndn3_42 | ~ndn3_40);
  assign n5854_1 = ~preset & n_n8678 & (~ndn3_42 | ndn3_44);
  assign n5855 = ~ndn3_44 & ndn3_42 & ~preset & n_n7948;
  assign n5856 = ~preset & n_n9432 & (~ndn3_42 | ndn3_44);
  assign n5857 = ~ndn3_44 & ndn3_42 & ~preset & n_n9036;
  assign n5858 = ~ndn3_2 & ~preset & psv38_5_5_ & n4949_1;
  assign n5859_1 = ~preset & n_n9174 & (ndn3_2 | ~n4949_1);
  assign n5860 = ~preset & n_n7757 & (ndn3_42 | ~ndn3_40);
  assign n5861 = ~preset & n_n7831 & (ndn3_30 | nsr3_30);
  assign n5862 = ~ndn3_2 & ~preset & psv13_5_5_ & n4949_1;
  assign n5863 = ~preset & n_n9501 & (ndn3_2 | ~n4949_1);
  assign n5864_1 = ~preset & n_n8445 & (nsr3_38 | ndn3_38);
  assign n5865 = ~ndn3_2 & ~preset & psv2_3_3_ & n4949_1;
  assign n5866 = ~preset & n_n9408 & (ndn3_2 | ~n4949_1);
  assign n5867 = ~preset & n_n9489 & (ndn3_30 | nsr3_30);
  assign n5868 = ~preset & n_n7821 & (ndn3_25 | ~ndn3_22);
  assign n5869_1 = ~preset & n4889_1 & (~n4971 ^ ~n4972);
  assign n5870 = ~preset & n_n7217 & (ngfdn_3 | ~ndn3_46);
  assign n5871 = ~preset & n_n9321 & (ndn3_7 | ~ndn3_4);
  assign n5872 = ~preset & n4879_1 & (~n4954_1 ^ ~n4955);
  assign n5873 = ~preset & n_n8843 & (nsr3_20 | ndn3_20);
  assign n5874_1 = ~preset & n_n7641 & (ndn3_23 | nsr3_23);
  assign n5875 = ~preset & n_n8258 & (ndn3_46 | ~ndn3_44);
  assign n5876 = ~preset & n_n8247 & (ndn3_42 | ~ndn3_40);
  assign n5877 = ~preset & n_n8957 & (~ndn3_39 | ndn3_40);
  assign n5878 = ~preset & n_n8959 & (~ndn3_39 | ndn3_40);
  assign n5879_1 = n4846 & (n5004_1 ^ (n6527 | n6528));
  assign n5880 = ~ndn3_2 & ~preset & psv26_8_8_ & n4949_1;
  assign n5881 = ~preset & n_n7954 & (ndn3_2 | ~n4949_1);
  assign n5882 = ~preset & n_n9601 & (ndn3_13 | nsr3_13);
  assign n5883 = ~preset & n_n9465 & (~ndn3_42 | ndn3_44);
  assign n5884_1 = ~ndn3_44 & ndn3_42 & ~preset & n_n8022;
  assign n5885 = ~ndn3_2 & ~preset & psv26_0_0_ & n4949_1;
  assign n5886 = ~preset & n_n7656 & (ndn3_2 | ~n4949_1);
  assign n5887 = ~preset & n_n8998 & (~ndn3_25 | ndn3_26);
  assign n5888 = ~preset & n_n8282 & (~ndn3_11 | ndn3_12);
  assign n5889_1 = ~preset & n4849_1 & (~n4985 ^ ~n4986);
  assign n5890 = ~preset & n_n7546 & (ngfdn_3 | ~ndn3_46);
  assign n5891 = ~ngfdn_3 & ~preset & n_n9235 & ndn3_46;
  assign n5892 = ~preset & n_n7174 & (ndn3_46 | ~ndn3_44);
  assign n5893 = n_n9632 & ndn3_44 & ~preset & ~ndn3_46;
  assign n5894_1 = ~preset & n_n8742 & (~ndn3_25 | ndn3_26);
  assign n5895 = ~preset & n4851 & (~n4954_1 ^ ~n4955);
  assign n5896 = ~preset & n_n8006 & (ndn3_7 | ~ndn3_4);
  assign n5897 = ~ndn3_2 & ~preset & psv13_13_13_ & n4949_1;
  assign n5898 = ~preset & n_n8414 & (ndn3_2 | ~n4949_1);
  assign n5899_1 = ~ndn3_2 & ~preset & psv13_8_8_ & n4949_1;
  assign n5900 = ~preset & n_n7955 & (ndn3_2 | ~n4949_1);
  assign n5901 = ~preset & n_n7160 & (~ndn3_39 | ndn3_40);
  assign n5902 = ~ndn3_40 & ndn3_39 & ~preset & n_n8906;
  assign n5903 = ~ndn3_2 & ~preset & psv33_13_13_ & n4949_1;
  assign n5904_1 = ~preset & n_n9098 & (ndn3_2 | ~n4949_1);
  assign n5905 = ~preset & n_n7640 & (~ndn3_29 | ndn3_32);
  assign n5906 = ~preset & n_n7803 & (ndn3_7 | ~ndn3_4);
  assign n5907 = ~preset & n4879_1 & (~n4976 ^ ~n4977);
  assign n5908 = ~ndn3_2 & ~preset & psv33_11_11_ & n4949_1;
  assign n5909_1 = ~preset & n_n8086 & (ndn3_2 | ~n4949_1);
  assign n5910 = ~preset & n_n9339 & (~nen3_22 | ndn3_22);
  assign n5911 = n4866 & (n4987 ^ (n6433 | n6434));
  assign n5912 = n4949_1 & ~ndn3_2 & pinp_4_4_ & ~preset;
  assign n5913 = ~preset & n_n8736 & (ndn3_2 | ~n4949_1);
  assign n5914_1 = ~preset & n_n8005 & (~nen3_16 | ndn3_16);
  assign n5915 = ~preset & n_n7823 & (~nen3_16 | ndn3_16);
  assign n5916 = ~preset & n4875 & (~n4971 ^ ~n4972);
  assign n5917 = ~preset & n_n8545 & (~ndn3_25 | ndn3_26);
  assign n5918 = ~preset & n4851 & (~n4976 ^ ~n4977);
  assign n5919_1 = ~preset & n_n8219 & (nsr3_20 | ndn3_20);
  assign n5920 = ~preset & n_n7236 & (~ndn3_19 | ndn3_21);
  assign n5921 = ~preset & n_n7428 & (ndn3_29 | ~ndn3_28);
  assign n5922 = ~preset & n4869_1 & (~n4971 ^ ~n4972);
  assign n5923 = ~preset & n_n9597 & (nsr3_20 | ndn3_20);
  assign n5924_1 = n4949_1 & ~ndn3_2 & pinp_10_10_ & ~preset;
  assign n5925 = ~preset & n_n8110 & (ndn3_2 | ~n4949_1);
  assign n5926 = ~preset & n_n9391 & (ndn3_42 | ~ndn3_40);
  assign n5927 = n4863 & (n4996 ^ (n6545 | n6546));
  assign n5928 = ~preset & n_n7758 & (ndn3_30 | nsr3_30);
  assign n5929_1 = ~preset & n_n8278 & (ndn3_29 | ~ndn3_28);
  assign n5930 = ~preset & n4869_1 & (~n4985 ^ ~n4986);
  assign n5931 = ~preset & n_n9125 & (~ndn3_42 | ndn3_44);
  assign n5932 = n4861 & (n4996 ^ (n6545 | n6546));
  assign n5933 = ~preset & n_n9169 & (ndn3_42 | ~ndn3_40);
  assign n5934_1 = n_n6974 & ndn3_40 & ~preset & ~ndn3_42;
  assign n5935 = ~ndn3_2 & ~preset & psv38_15_15_ & n4949_1;
  assign n5936 = ~preset & n_n9223 & (ndn3_2 | ~n4949_1);
  assign n5937 = ~preset & n_n9135 & (ndn3_4 | ~ndn3_2);
  assign n5938 = ~preset & n_n7898 & (~ndn3_42 | ndn3_44);
  assign n5939_1 = ~preset & n_n8765 & (ndn3_46 | ~ndn3_44);
  assign n5940 = ~preset & n_n7908 & (ndn3_37 | nsr3_37);
  assign n5941 = ~preset & n_n7462 & (~ngfdn_3 | ndn3_50);
  assign n5942 = ~ndn3_50 & n_n9219 & ~preset & ngfdn_3;
  assign n5943 = ~preset & n_n7384 & (ndn3_46 | ~ndn3_44);
  assign n5944_1 = ~preset & n_n9613 & (~nen3_39 | ndn3_39);
  assign n5945 = ~preset & n4854_1 & (~n4985 ^ ~n4986);
  assign n5946 = ~ndn3_2 & ~preset & psv13_3_3_ & n4949_1;
  assign n5947 = ~preset & n_n9406 & (ndn3_2 | ~n4949_1);
  assign n5948 = ~preset & n_n9611 & (~nen3_39 | ndn3_39);
  assign n5949_1 = ~preset & n_n7324 & (ngfdn_3 | ~ndn3_46);
  assign n5950 = ~preset & n_n9335 & (ndn3_37 | nsr3_37);
  assign n5951 = ~preset & n_n9127 & (ndn3_37 | nsr3_37);
  assign n5952 = ~ngfdn_3 & nsr1_2 & (~preset_0_0_ | nlc1_2);
  assign n5953 = ~preset & n_n9400 & (~nen3_16 | ndn3_16);
  assign n5954_1 = ~preset & n_n9343 & (nsr3_13 | ndn3_15);
  assign n5955 = ~preset & n_n7054 & (ndn3_42 | ~ndn3_40);
  assign n5956 = ~ndn3_42 & ~preset & n_n9576 & ndn3_40;
  assign n5957 = ~preset & n_n7948 & (ndn3_42 | ~ndn3_40);
  assign n5958 = ~preset & n_n7783 & (ndn3_46 | ~ndn3_44);
  assign n5959_1 = n4853 & (n5004_1 ^ (n6527 | n6528));
  assign n5960 = ~preset & n_n7602 & (ndn3_23 | nsr3_23);
  assign n5961 = ~preset & n_n7740 & (nsr3_20 | ndn3_20);
  assign n5962 = ~preset & n_n7691 & (~ndn3_42 | ndn3_44);
  assign n5963 = ~preset & n_n9483 & (~ngfdn_3 | ndn3_50);
  assign n5964_1 = ~ndn3_50 & ~preset & ngfdn_3 & n_n8948;
  assign n5965 = ~preset & n_n9049 & (nsr3_14 | ndn3_14);
  assign n5966 = ~preset & n_n9588 & (ndn3_34 | ~nen3_34);
  assign n5967 = ~preset & n4860 & (~n4969_1 ^ ~n4970);
  assign n5968 = ~preset & n_n7791 & (~ndn3_9 | ndn3_11);
  assign n5969_1 = ~preset & n_n7857 & (ndn3_46 | ~ndn3_44);
  assign n5970 = ~ndn3_46 & ~preset & n_n7706 & ndn3_44;
  assign n5971 = n4900 & (n5975 | (n4975 & n7176));
  assign n5972 = n4856 & (~n_n8631 ^ (n_n8561 | n4999_1));
  assign n5973 = n4897 & (n5975 | (n4975 & n7176));
  assign n5974_1 = n4856 & (n_n8913 ^ ~n4968);
  assign n5975 = n7089 & n4967 & ~preset & ~n_n9247;
  assign n5976 = ~ndn3_2 & ~preset & psv13_14_14_ & n4949_1;
  assign n5977 = ~preset & n_n8114 & (ndn3_2 | ~n4949_1);
  assign n5978 = ~ndn3_2 & ~preset & psv39_15_15_ & n4949_1;
  assign n5979_1 = ~preset & n_n8491 & (ndn3_2 | ~n4949_1);
  assign n5980 = ~preset & n_n8175 & (~nen3_22 | ndn3_22);
  assign n5981 = ~ndn3_22 & ~preset & nen3_22 & n_n9252;
  assign n5982 = ~preset & n_n9257 & (ndn3_13 | nsr3_13);
  assign n5983 = ~preset & n_n8091 & (~ngfdn_3 | ndn3_50);
  assign n5984_1 = ~ndn3_50 & n_n8466 & ~preset & ngfdn_3;
  assign n5985 = ~preset & n_n8066 & (nsr3_14 | ndn3_14);
  assign n5986 = ~ndn3_2 & ~preset & psv13_2_2_ & n4949_1;
  assign n5987 = ~preset & n_n8053 & (ndn3_2 | ~n4949_1);
  assign n5988 = ~preset & n_n7811 & (nsr3_13 | ndn3_15);
  assign n5989_1 = ~preset & n_n7934 & (ndn3_13 | nsr3_13);
  assign n5990 = ~preset & n_n7735 & (ndn3_30 | nsr3_30);
  assign n5991 = ~preset & n_n7651 & (ndn3_30 | nsr3_30);
  assign n5992 = ~preset & n_n9412 & (~ndn3_19 | ndn3_21);
  assign n5993 = ~preset & n_n9398 & (~nen3_22 | ndn3_22);
  assign n5994_1 = n4866 & (n4996 ^ (n6545 | n6546));
  assign n5995 = ~preset & n_n9064 & (nsr3_20 | ndn3_20);
  assign n5996 = ~ndn3_2 & ~preset & psv2_15_15_ & n4949_1;
  assign n5997 = ~preset & n_n8007 & (ndn3_2 | ~n4949_1);
  assign n5998 = n4949_1 & ~ndn3_2 & pinp_15_15_ & ~preset;
  assign n5999_1 = ~preset & n_n8482 & (ndn3_2 | ~n4949_1);
  assign n6000 = ~ndn3_2 & ~preset & psv2_14_14_ & n4949_1;
  assign n6001 = ~preset & n_n7937 & (ndn3_2 | ~n4949_1);
  assign n6002 = n4949_1 & ~ndn3_2 & pinp_13_13_ & ~preset;
  assign n6003 = ~preset & n_n7850 & (ndn3_2 | ~n4949_1);
  assign n6004_1 = n7175 & ((n4918 & n4919_1) | (n_n9512 & (n4918 | n4919_1)));
  assign n6005 = ~n_n9434 & n4857 & (~n4893 ^ ~n4894_1);
  assign n6006 = ~n4894_1 & ~n4893 & n_n9434 & n4856;
  assign n6007 = ~n5001 & ~preset & n_n9434;
  assign n6008 = ~preset & n_n9399 & (nsr3_20 | ndn3_20);
  assign n6009_1 = ~preset & n_n8333 & (ndn3_28 | ~nen3_28);
  assign n6010 = ~preset & n4892 & (~n4985 ^ ~n4986);
  assign n6011 = ~ndn3_2 & ~preset & psv18_11_11_ & n4949_1;
  assign n6012 = ~preset & n_n7759 & (ndn3_2 | ~n4949_1);
  assign n6013 = ~preset & n_n8661 & (nsr3_14 | ndn3_14);
  assign n6014_1 = ~preset & n_n8132 & (ndn3_42 | ~ndn3_40);
  assign n6015 = ~ndn3_42 & ~preset & n_n8150 & ndn3_40;
  assign n6016 = ~preset & n_n8488 & (~nen3_22 | ndn3_22);
  assign n6017 = ~ndn3_22 & n_n9412 & ~preset & nen3_22;
  assign n6018 = ~preset & n_n7953 & (ndn3_13 | nsr3_13);
  assign n6019_1 = ~preset & n_n7179 & (ngfdn_3 | ~ndn3_46);
  assign n6020 = ndn3_46 & n_n7783 & ~preset & ~ngfdn_3;
  assign n6021 = ~preset & n_n9265 & (~ndn3_17 | ndn3_18);
  assign n6022 = ~preset & n4877 & (~n4969_1 ^ ~n4970);
  assign n6023 = ~preset & n_n9052 & (ndn3_4 | ~ndn3_2);
  assign n6024_1 = ~preset & n4874_1 & (~n4954_1 ^ ~n4955);
  assign n6025 = ~preset & n_n9106 & (~nen3_39 | ndn3_39);
  assign n6026 = ~preset & n4854_1 & (~n4954_1 ^ ~n4955);
  assign n6027 = ~preset & n_n8702 & (~nen3_22 | ndn3_22);
  assign n6028 = ~ndn3_22 & ~preset & nen3_22 & n_n8213;
  assign n6029_1 = ~preset & n_n7190 & (~ndn3_42 | ndn3_44);
  assign n6030 = ~ndn3_44 & ndn3_42 & ~preset & n_n8249;
  assign n6031 = ~preset & n_n9635 & (~ndn3_42 | ndn3_44);
  assign n6032 = n4861 & (n4980 ^ (n6352 | n6353));
  assign n6033 = ~preset & n_n8001 & (nsr3_38 | ndn3_38);
  assign n6034_1 = ~preset & n_n9000 & (ndn3_25 | ~ndn3_22);
  assign n6035 = ~preset & n_n9598 & (~nen3_16 | ndn3_16);
  assign n6036 = ~preset & n4875 & (~n4969_1 ^ ~n4970);
  assign n6037 = ~preset & n_n8786 & (ndn3_7 | ~ndn3_4);
  assign n6038 = ~preset & n_n9602 & (ndn3_7 | ~ndn3_4);
  assign n6039_1 = ~preset & n4879_1 & (~n4969_1 ^ ~n4970);
  assign n6040 = ~preset & n_n8981 & (ndn3_29 | ~ndn3_28);
  assign n6041 = ~preset & n_n8308 & (ndn3_46 | ~ndn3_44);
  assign n6042 = ~preset & n_n8609 & (ndn3_42 | ~ndn3_40);
  assign n6043 = n4863 & (n5004_1 ^ (n6527 | n6528));
  assign n6044_1 = ~preset & n_n8699 & (nsr3_20 | ndn3_20);
  assign n6045 = ~preset & n_n8533 & (ndn3_23 | nsr3_23);
  assign n6046 = ~preset & n_n9273 & (~ndn3_19 | ndn3_21);
  assign n6047 = ~preset & n_n9311 & (nsr3_35 | ndn3_35);
  assign n6048 = ~preset & n_n7148 & (~ndn3_42 | ndn3_44);
  assign n6049_1 = ~ndn3_44 & ndn3_42 & ~preset & n_n9623;
  assign n6050 = ~preset & n_n8227 & (~ndn3_11 | ndn3_12);
  assign n6051 = ~preset & n_n7970 & (~ndn3_9 | ndn3_11);
  assign n6052 = ~preset & n_n7581 & (~nen3_22 | ndn3_22);
  assign n6053 = ~ndn3_22 & ~preset & nen3_22 & n_n9351;
  assign n6054_1 = ~preset & n_n9008 & (ndn3_9 | ~ndn3_7);
  assign n6055 = ~preset & n4852 & (~n4971 ^ ~n4972);
  assign n6056 = ~ndn3_2 & ~preset & psv26_12_12_ & n4949_1;
  assign n6057 = ~preset & n_n7814 & (ndn3_2 | ~n4949_1);
  assign n6058 = ~preset & n_n7877 & (~ndn3_11 | ndn3_12);
  assign n6059_1 = ~ndn3_2 & ~preset & psv26_11_11_ & n4949_1;
  assign n6060 = ~preset & n_n7765 & (ndn3_2 | ~n4949_1);
  assign n6061 = ~preset & n_n8758 & (ndn3_7 | ~ndn3_4);
  assign n6062 = ~preset & n4879_1 & (~n4985 ^ ~n4986);
  assign n6063 = ~preset & n_n7332 & (~ndn3_39 | ndn3_40);
  assign n6064_1 = ~ndn3_40 & ~preset & ndn3_39 & n_n8991;
  assign n6065 = ~ndn3_2 & ~preset & psv39_12_12_ & n4949_1;
  assign n6066 = ~preset & n_n7816 & (ndn3_2 | ~n4949_1);
  assign n6067 = ~preset & n_n7812 & (ndn3_13 | nsr3_13);
  assign n6068 = ~preset & n_n8394 & (ndn3_13 | nsr3_13);
  assign n6069_1 = ~preset & n_n8152 & (ndn3_17 | ~ndn3_16);
  assign n6070 = ~preset & n4882 & (~n4976 ^ ~n4977);
  assign n6071 = ~preset & n_n8597 & (~ndn3_17 | ndn3_18);
  assign n6072 = ~preset & n4877 & (~n4976 ^ ~n4977);
  assign n6073 = ~preset & n_n7889 & (nsr3_13 | ndn3_15);
  assign n6074_1 = ~preset & n4881 & (~n4985 ^ ~n4986);
  assign n6075 = ~preset & n_n7888 & (~nen3_16 | ndn3_16);
  assign n6076 = ~preset & n4875 & (~n4985 ^ ~n4986);
  assign n6077 = ~preset & n_n8225 & (ndn3_19 | ~nen3_19);
  assign n6078 = ~preset & n_n7599 & (ndn3_37 | nsr3_37);
  assign n6079_1 = ~preset & n_n7558 & (ngfdn_3 | ~ndn3_46);
  assign n6080 = n1270 & (n4996 ^ (n6545 | n6546));
  assign n6081 = ~preset & n_n8377 & (ndn3_7 | ~ndn3_4);
  assign n6082 = ~preset & n_n8208 & (~ndn3_17 | ndn3_18);
  assign n6083 = n4952 & ((n4994_1 & n4995) | (n4986 & (~n4994_1 ^ ~n4995)));
  assign n6084_1 = (n7157 | n7158) & (n7164 | n7165);
  assign n6085 = n_n9568 & ((nen3_22 & ~ndn3_22) | n6899);
  assign n6086 = n_n8772 & (n6900 | (~ndn3_17 & ndn3_16));
  assign n6087 = n_n7914 & ~ndn3_7 & ndn3_4;
  assign n6088 = n_n7913 & ndn3_11 & ~ndn3_12;
  assign n6089_1 = ndn3_40 & n_n7908 & ~ndn3_42;
  assign n6090 = ndn3_26 & ~ndn3_27 & n_n7932;
  assign n6091 = n_n9632 & ~ngfdn_3 & ndn3_46;
  assign n6092 = n_n8535 & nen3_16 & ~ndn3_16;
  assign n6093 = ~ndn3_32 & ndn3_29 & n_n7910;
  assign n6094_1 = ~ndn3_40 & n_n7909 & ndn3_39;
  assign n6095 = n_n7912 & ndn3_19 & ~ndn3_21;
  assign n6096 = n_n7911 & ~ndn3_25 & ndn3_22;
  assign n6097 = ndn3_44 & n_n8512 & ~ndn3_46;
  assign n6098 = n_n8106 & ndn3_17 & ~ndn3_18;
  assign n6099 = n_n7935 & ((nen3_16 & ~ndn3_16) | n6908);
  assign n6100 = n_n7936 & ((~ndn3_25 & ndn3_22) | n6909);
  assign n6101 = ndn3_2 & n_n7937 & ~ndn3_4;
  assign n6102 = n_n7928 & nen3_39 & ~ndn3_39;
  assign n6103 = ndn3_7 & ~ndn3_9 & n_n8114;
  assign n6104 = ndn3_46 & ~ngfdn_3 & n_n9108;
  assign n6105 = n_n7946 & ndn3_9 & ~ndn3_11;
  assign n6106 = n_n7933 & ndn3_19 & ~ndn3_21;
  assign n6107 = nen3_28 & n_n7931 & ~ndn3_28;
  assign n6108 = n_n7927 & ~ndn3_46 & ndn3_44;
  assign n6109 = ~ndn3_44 & n_n8445 & ndn3_42;
  assign n6110 = nen3_34 & ~ndn3_34 & n_n8425;
  assign n6111 = ~ndn3_36 & nen3_36 & n_n7929;
  assign n6112 = n_n8516 & ndn3_17 & ~ndn3_18;
  assign n6113 = n_n8219 & nen3_22 & ~ndn3_22;
  assign n6114 = ~ndn3_15 & n_n7934 & ~nsr3_13;
  assign n6115 = n_n7971 & ((nen3_22 & ~ndn3_22) | n6899);
  assign n6116 = n_n8014 & ((~ndn3_17 & ndn3_16) | n6900);
  assign n6117 = ndn3_4 & ~ndn3_7 & n_n8456;
  assign n6118 = ~ndn3_12 & n_n7970 & ndn3_11;
  assign n6119 = ndn3_40 & n_n7966 & ~ndn3_42;
  assign n6120 = ndn3_26 & ~ndn3_27 & n_n8004;
  assign n6121 = n_n8468 & ~ngfdn_3 & ndn3_46;
  assign n6122 = n_n7969 & nen3_16 & ~ndn3_16;
  assign n6123 = ~ndn3_32 & ndn3_29 & n_n9077;
  assign n6124 = ~ndn3_40 & n_n7967 & ndn3_39;
  assign n6125 = ~ndn3_21 & n_n8208 & ndn3_19;
  assign n6126 = n_n7968 & ~ndn3_25 & ndn3_22;
  assign n6127 = ndn3_44 & n_n8864 & ~ndn3_46;
  assign n6128 = n_n8519 & ndn3_17 & ~ndn3_18;
  assign n6129 = n_n8006 & (n6908 | (nen3_16 & ~ndn3_16));
  assign n6130 = n_n8491 & (n6909 | (~ndn3_25 & ndn3_22));
  assign n6131 = ndn3_2 & n_n8007 & ~ndn3_4;
  assign n6132 = n_n8078 & nen3_39 & ~ndn3_39;
  assign n6133 = n_n8502 & ~ndn3_9 & ndn3_7;
  assign n6134 = n_n8580 & ~ngfdn_3 & ndn3_46;
  assign n6135 = n_n8192 & ndn3_9 & ~ndn3_11;
  assign n6136 = ~ndn3_21 & n_n8005 & ndn3_19;
  assign n6137 = nen3_28 & ~ndn3_28 & n_n8003;
  assign n6138 = ndn3_44 & ~ndn3_46 & n_n9355;
  assign n6139 = ~ndn3_44 & n_n8001 & ndn3_42;
  assign n6140 = nen3_34 & ~ndn3_34 & n_n8839;
  assign n6141 = ~ndn3_36 & nen3_36 & n_n8900;
  assign n6142 = n_n8584 & ndn3_17 & ~ndn3_18;
  assign n6143 = n_n8064 & nen3_22 & ~ndn3_22;
  assign n6144 = n_n8344 & ~nsr3_13 & ~ndn3_15;
  assign n6145 = ~preset & n_n8775 & (ndn3_4 | ~ndn3_2);
  assign n6146 = ~preset & n4874_1 & (~n4985 ^ ~n4986);
  assign n6147 = n_n8758 & (n6908 | (nen3_16 & ~ndn3_16));
  assign n6148 = n_n8504 & ((~ndn3_25 & ndn3_22) | n6909);
  assign n6149 = ndn3_2 & ~ndn3_4 & n_n7890;
  assign n6150 = ~ndn3_39 & nen3_39 & n_n7988;
  assign n6151 = ndn3_7 & ~ndn3_9 & n_n8414;
  assign n6152 = ndn3_46 & ~ngfdn_3 & n_n8626;
  assign n6153 = n_n9067 & ndn3_9 & ~ndn3_11;
  assign n6154 = ~ndn3_21 & n_n7888 & ndn3_19;
  assign n6155 = nen3_28 & ~ndn3_28 & n_n7887;
  assign n6156 = ndn3_44 & n_n9623 & ~ndn3_46;
  assign n6157 = ~ndn3_44 & n_n7885 & ndn3_42;
  assign n6158 = nen3_34 & n_n8333 & ~ndn3_34;
  assign n6159 = n_n9092 & nen3_36 & ~ndn3_36;
  assign n6160 = n_n8282 & ndn3_17 & ~ndn3_18;
  assign n6161 = ~ndn3_22 & nen3_22 & n_n9064;
  assign n6162 = ~ndn3_15 & n_n8394 & ~nsr3_13;
  assign n6163 = n_n8775 & (n6899 | (nen3_22 & ~ndn3_22));
  assign n6164 = n_n7849 & ((~ndn3_17 & ndn3_16) | n6900);
  assign n6165 = ndn3_4 & n_n9098 & ~ndn3_7;
  assign n6166 = n_n7848 & ndn3_11 & ~ndn3_12;
  assign n6167 = ndn3_40 & n_n8480 & ~ndn3_42;
  assign n6168 = ndn3_26 & ~ndn3_27 & n_n9520;
  assign n6169 = n_n8470 & ~ngfdn_3 & ndn3_46;
  assign n6170 = n_n8909 & nen3_16 & ~ndn3_16;
  assign n6171 = ~ndn3_32 & ndn3_29 & n_n7845;
  assign n6172 = n_n7844 & ndn3_39 & ~ndn3_40;
  assign n6173 = ~ndn3_21 & n_n7847 & ndn3_19;
  assign n6174 = n_n7846 & ~ndn3_25 & ndn3_22;
  assign n6175 = ndn3_44 & ~ndn3_46 & n_n8277;
  assign n6176 = ~ndn3_18 & n_n7889 & ndn3_17;
  assign n6177 = ~preset & n_n7452 & (ndn3_29 | ~ndn3_28);
  assign n6178 = n7123 & ((n4934_1 & n4937) | (n_n8821 & (n4934_1 | n4937)));
  assign n6179 = ~n_n9638 & n4857 & (~n4870 ^ ~n4871);
  assign n6180 = ~n4871 & ~n4870 & n_n9638 & n4856;
  assign n6181 = ~n5001 & ~preset & n_n9638;
  assign n6182 = ~preset & n_n7522 & (ndn3_42 | ~ndn3_40);
  assign n6183 = ~ndn3_42 & ~preset & n_n9102 & ndn3_40;
  assign n6184 = ~preset & n_n9235 & (ndn3_46 | ~ndn3_44);
  assign n6185 = ~preset & n_n9486 & (ndn3_42 | ~ndn3_40);
  assign n6186 = ~preset & n_n9130 & (ndn3_23 | nsr3_23);
  assign n6187 = ~ndn3_2 & ~preset & psv38_11_11_ & n4949_1;
  assign n6188 = ~preset & n_n7709 & (ndn3_2 | ~n4949_1);
  assign n6189 = ~preset & n_n7819 & (nsr3_35 | ndn3_35);
  assign n6190 = ~ndn3_2 & ~preset & psv18_15_15_ & n4949_1;
  assign n6191 = ~preset & n_n8002 & (ndn3_2 | ~n4949_1);
  assign n6192 = ~preset & n_n9467 & (ndn3_34 | ~nen3_34);
  assign n6193 = ~preset & n4860 & (~n4976 ^ ~n4977);
  assign n6194 = ~preset & n_n9548 & (ngfdn_3 | ~ndn3_46);
  assign n6195 = ndn3_46 & n_n7384 & ~preset & ~ngfdn_3;
  assign n6196 = ~preset & n_n7707 & (ndn3_37 | nsr3_37);
  assign n6197 = ~n5001 & ~preset & n_n8557;
  assign n6198 = n_n8584 & (nsr3_13 ? ndn3_12 : nsr3_14);
  assign n6199 = nsr3_20 & ndn3_17 & n_n8583;
  assign n6200 = nsr3_35 & ndn3_29 & n_n8941;
  assign n6201 = nen3_34 & n_n8864 & nsr3_37;
  assign n6202 = ndn3_26 & nsr3_30 & n_n8581;
  assign n6203 = n_n8580 & nsr3_38 & nen3_36;
  assign n6204 = ndn3_19 & nsr3_23 & n_n8582;
  assign n6205 = n_n8227 & (nsr3_13 ? ndn3_12 : nsr3_14);
  assign n6206 = n_n8226 & ndn3_17 & nsr3_20;
  assign n6207 = n_n8224 & ndn3_29 & nsr3_35;
  assign n6208 = nen3_34 & n_n8223 & nsr3_37;
  assign n6209 = ndn3_26 & nsr3_30 & n_n9205;
  assign n6210 = n_n8222 & nsr3_38 & nen3_36;
  assign n6211 = ndn3_19 & n_n8225 & nsr3_23;
  assign n6212 = n_n8203 & (nsr3_13 ? ndn3_12 : nsr3_14);
  assign n6213 = nsr3_20 & ndn3_17 & n_n9019;
  assign n6214 = n_n8201 & ndn3_29 & nsr3_35;
  assign n6215 = nen3_34 & n_n9110 & nsr3_37;
  assign n6216 = ndn3_26 & nsr3_30 & n_n9615;
  assign n6217 = n_n9516 & nsr3_38 & nen3_36;
  assign n6218 = ndn3_19 & n_n8202 & nsr3_23;
  assign n6219 = n_n7951 & (nsr3_13 ? ndn3_12 : nsr3_14);
  assign n6220 = nsr3_20 & ndn3_17 & n_n8753;
  assign n6221 = nsr3_35 & ndn3_29 & n_n7474;
  assign n6222 = nen3_34 & n_n9518 & nsr3_37;
  assign n6223 = ndn3_26 & nsr3_30 & n_n9286;
  assign n6224 = n_n7947 & nsr3_38 & nen3_36;
  assign n6225 = n_n7588 & nsr3_23 & ndn3_19;
  assign n6226 = n_n9141 & (nsr3_13 ? ndn3_12 : nsr3_14);
  assign n6227 = nsr3_20 & ndn3_17 & n_n7375;
  assign n6228 = nsr3_35 & n_n7373 & ndn3_29;
  assign n6229 = nen3_34 & n_n8499 & nsr3_37;
  assign n6230 = ndn3_26 & nsr3_30 & n_n7487;
  assign n6231 = n_n8135 & nsr3_38 & nen3_36;
  assign n6232 = n_n7374 & nsr3_23 & ndn3_19;
  assign n6233 = n_n9015 & (nsr3_13 ? ndn3_12 : nsr3_14);
  assign n6234 = nsr3_20 & ndn3_17 & n_n8104;
  assign n6235 = n_n8828 & ndn3_29 & nsr3_35;
  assign n6236 = nen3_34 & n_n7670 & nsr3_37;
  assign n6237 = ndn3_26 & n_n7341 & nsr3_30;
  assign n6238 = nen3_36 & n_n8862 & nsr3_38;
  assign n6239 = n_n7342 & nsr3_23 & ndn3_19;
  assign n6240 = n_n9318 & (nsr3_13 ? ndn3_12 : nsr3_14);
  assign n6241 = nsr3_20 & ndn3_17 & n_n8744;
  assign n6242 = nsr3_35 & ndn3_29 & n_n8741;
  assign n6243 = nen3_34 & n_n9042 & nsr3_37;
  assign n6244 = ndn3_26 & n_n8742 & nsr3_30;
  assign n6245 = n_n9308 & nsr3_38 & nen3_36;
  assign n6246 = n_n8743 & nsr3_23 & ndn3_19;
  assign n6247 = n_n9401 & (nsr3_13 ? ndn3_12 : nsr3_14);
  assign n6248 = n_n8811 & ndn3_17 & nsr3_20;
  assign n6249 = nsr3_35 & ndn3_29 & n_n8808;
  assign n6250 = nen3_34 & n_n9126 & nsr3_37;
  assign n6251 = ndn3_26 & nsr3_30 & n_n8809;
  assign n6252 = n_n9390 & nsr3_38 & nen3_36;
  assign n6253 = n_n8810 & nsr3_23 & ndn3_19;
  assign n6254 = n_n7824 & (nsr3_13 ? ndn3_12 : nsr3_14);
  assign n6255 = nsr3_20 & ndn3_17 & n_n8729;
  assign n6256 = nsr3_35 & ndn3_29 & n_n7428;
  assign n6257 = nen3_34 & n_n7598 & nsr3_37;
  assign n6258 = n_n7485 & nsr3_30 & ndn3_26;
  assign n6259 = n_n8898 & nsr3_38 & nen3_36;
  assign n6260 = n_n7429 & nsr3_23 & ndn3_19;
  assign n6261 = n_n9496 & (nsr3_13 ? ndn3_12 : nsr3_14);
  assign n6262 = nsr3_20 & ndn3_17 & n_n8884;
  assign n6263 = n_n8881 & ndn3_29 & nsr3_35;
  assign n6264 = nen3_34 & n_n9473 & nsr3_37;
  assign n6265 = ndn3_26 & n_n8882 & nsr3_30;
  assign n6266 = nen3_36 & n_n9485 & nsr3_38;
  assign n6267 = ndn3_19 & n_n8883 & nsr3_23;
  assign n6268 = n_n7877 & (nsr3_13 ? ndn3_12 : nsr3_14);
  assign n6269 = nsr3_20 & ndn3_17 & n_n8727;
  assign n6270 = nsr3_35 & n_n7452 & ndn3_29;
  assign n6271 = nen3_34 & n_n7640 & nsr3_37;
  assign n6272 = n_n7453 & nsr3_30 & ndn3_26;
  assign n6273 = n_n9458 & nsr3_38 & nen3_36;
  assign n6274 = ndn3_19 & nsr3_23 & n_n7454;
  assign n6275 = n_n9599 & (nsr3_13 ? ndn3_12 : nsr3_14);
  assign n6276 = nsr3_20 & ndn3_17 & n_n8939;
  assign n6277 = n_n8937 & ndn3_29 & nsr3_35;
  assign n6278 = nen3_34 & n_n9470 & nsr3_37;
  assign n6279 = ndn3_26 & nsr3_30 & n_n8938;
  assign n6280 = nen3_36 & n_n9588 & nsr3_38;
  assign n6281 = n_n9139 & nsr3_23 & ndn3_19;
  assign n6282 = n_n8984 & (nsr3_13 ? ndn3_12 : nsr3_14);
  assign n6283 = nsr3_20 & ndn3_17 & n_n8983;
  assign n6284 = nsr3_35 & n_n8981 & ndn3_29;
  assign n6285 = nen3_34 & n_n9334 & nsr3_37;
  assign n6286 = ndn3_26 & n_n8998 & nsr3_30;
  assign n6287 = n_n8980 & nsr3_38 & nen3_36;
  assign n6288 = n_n8982 & nsr3_23 & ndn3_19;
  assign n6289 = n_n8153 & (nsr3_13 ? ndn3_12 : nsr3_14);
  assign n6290 = nsr3_20 & n_n8152 & ndn3_17;
  assign n6291 = n_n8177 & ndn3_29 & nsr3_35;
  assign n6292 = nen3_34 & nsr3_37 & n_n8628;
  assign n6293 = ndn3_26 & n_n8545 & nsr3_30;
  assign n6294 = nen3_36 & n_n9467 & nsr3_38;
  assign n6295 = n_n8151 & nsr3_23 & ndn3_19;
  assign n6296 = n_n8282 & (nsr3_13 ? ndn3_12 : nsr3_14);
  assign n6297 = nsr3_20 & ndn3_17 & n_n8281;
  assign n6298 = nsr3_35 & ndn3_29 & n_n8278;
  assign n6299 = nen3_34 & n_n8277 & nsr3_37;
  assign n6300 = ndn3_26 & n_n8279 & nsr3_30;
  assign n6301 = n_n8626 & nsr3_38 & nen3_36;
  assign n6302 = n_n8280 & nsr3_23 & ndn3_19;
  assign n6303 = n_n8516 & (nsr3_13 ? ndn3_12 : nsr3_14);
  assign n6304 = nsr3_20 & ndn3_17 & n_n8515;
  assign n6305 = n_n8513 & ndn3_29 & nsr3_35;
  assign n6306 = nen3_34 & n_n8512 & nsr3_37;
  assign n6307 = ndn3_26 & nsr3_30 & n_n9203;
  assign n6308 = n_n9108 & nsr3_38 & nen3_36;
  assign n6309 = n_n8514 & nsr3_23 & ndn3_19;
  assign n6310 = ~preset & n_n6991 & (ngfdn_3 | ~ndn3_46);
  assign n6311 = ndn3_46 & n_n7896 & ~preset & ~ngfdn_3;
  assign n6312 = ~preset & n_n7271 & (ngfdn_3 | ~ndn3_46);
  assign n6313 = ~ngfdn_3 & ~preset & n_n8308 & ndn3_46;
  assign n6314 = ~preset & n_n7252 & (ngfdn_3 | ~ndn3_46);
  assign n6315 = n_n7444 & ndn3_46 & ~preset & ~ngfdn_3;
  assign n6316 = ~preset & n_n8871 & (~nen3_39 | ndn3_39);
  assign n6317 = ~preset & n_n8592 & (ndn3_46 | ~ndn3_44);
  assign n6318 = ~ndn3_46 & ~preset & n_n9259 & ndn3_44;
  assign n6319 = ~preset & n_n9401 & (~ndn3_11 | ndn3_12);
  assign n6320 = ~preset & n_n8150 & (~ndn3_39 | ndn3_40);
  assign n6321 = n4846 & (n4980 ^ (n6352 | n6353));
  assign n6322 = n_n7813 & ((nen3_16 & ~ndn3_16) | n6908);
  assign n6323 = n_n7816 & (n6909 | (~ndn3_25 & ndn3_22));
  assign n6324 = ndn3_2 & n_n7817 & ~ndn3_4;
  assign n6325 = ~ndn3_39 & nen3_39 & n_n7807;
  assign n6326 = n_n7815 & ~ndn3_9 & ndn3_7;
  assign n6327 = ndn3_46 & ~ngfdn_3 & n_n8222;
  assign n6328 = ~ndn3_11 & n_n7814 & ndn3_9;
  assign n6329 = n_n7810 & ndn3_19 & ~ndn3_21;
  assign n6330 = nen3_28 & ~ndn3_28 & n_n8473;
  assign n6331 = ndn3_44 & n_n8022 & ~ndn3_46;
  assign n6332 = ~ndn3_44 & n_n7806 & ndn3_42;
  assign n6333 = nen3_34 & ~ndn3_34 & n_n7859;
  assign n6334 = ~ndn3_36 & nen3_36 & n_n7808;
  assign n6335 = ~ndn3_18 & n_n8227 & ndn3_17;
  assign n6336 = n_n8657 & nen3_22 & ~ndn3_22;
  assign n6337 = ~ndn3_15 & n_n7812 & ~nsr3_13;
  assign n6338 = n_n7793 & ((nen3_22 & ~ndn3_22) | n6899);
  assign n6339 = n_n7792 & ((~ndn3_17 & ndn3_16) | n6900);
  assign n6340 = n_n8267 & ~ndn3_7 & ndn3_4;
  assign n6341 = ~ndn3_12 & n_n7791 & ndn3_11;
  assign n6342 = n_n7788 & ~ndn3_42 & ndn3_40;
  assign n6343 = ndn3_26 & ~ndn3_27 & n_n7809;
  assign n6344 = ndn3_46 & n_n9635 & ~ngfdn_3;
  assign n6345 = n_n9525 & nen3_16 & ~ndn3_16;
  assign n6346 = ~ndn3_32 & ndn3_29 & n_n7790;
  assign n6347 = ~ndn3_40 & n_n7789 & ndn3_39;
  assign n6348 = n_n8402 & ndn3_19 & ~ndn3_21;
  assign n6349 = n_n8841 & ~ndn3_25 & ndn3_22;
  assign n6350 = ndn3_44 & n_n8223 & ~ndn3_46;
  assign n6351 = ~ndn3_18 & ndn3_17 & n_n7811;
  assign n6352 = (n7062 | n7063) & (n7069 | n7070);
  assign n6353 = n5002 & ((n4988 & n4989_1) | (n4976 & (n4988 ^ n4989_1)));
  assign n6354 = ~ndn3_2 & ~preset & psv2_5_5_ & n4949_1;
  assign n6355 = ~preset & n_n9503 & (ndn3_2 | ~n4949_1);
  assign n6356 = ~preset & n_n7779 & (ngfdn_3 | ~ndn3_46);
  assign n6357 = n_n7764 & ((nen3_16 & ~ndn3_16) | n6908);
  assign n6358 = n_n8506 & ((~ndn3_25 & ndn3_22) | n6909);
  assign n6359 = ndn3_2 & n_n9387 & ~ndn3_4;
  assign n6360 = n_n7990 & nen3_39 & ~ndn3_39;
  assign n6361 = n_n7766 & ~ndn3_9 & ndn3_7;
  assign n6362 = n_n9516 & ~ngfdn_3 & ndn3_46;
  assign n6363 = ~ndn3_11 & n_n7765 & ndn3_9;
  assign n6364 = n_n7762 & ndn3_19 & ~ndn3_21;
  assign n6365 = n_n8852 & ~ndn3_28 & nen3_28;
  assign n6366 = ndn3_44 & n_n7757 & ~ndn3_46;
  assign n6367 = ~ndn3_44 & n_n7918 & ndn3_42;
  assign n6368 = nen3_34 & n_n9157 & ~ndn3_34;
  assign n6369 = ~ndn3_36 & n_n7758 & nen3_36;
  assign n6370 = n_n8203 & ndn3_17 & ~ndn3_18;
  assign n6371 = n_n7761 & nen3_22 & ~ndn3_22;
  assign n6372 = n_n8396 & ~nsr3_13 & ~ndn3_15;
  assign n6373 = n_n7901 & ((nen3_22 & ~ndn3_22) | n6899);
  assign n6374 = n_n7713 & (n6900 | (~ndn3_17 & ndn3_16));
  assign n6375 = ndn3_4 & n_n8086 & ~ndn3_7;
  assign n6376 = n_n9210 & ndn3_11 & ~ndn3_12;
  assign n6377 = ndn3_40 & n_n7707 & ~ndn3_42;
  assign n6378 = ndn3_26 & n_n7760 & ~ndn3_27;
  assign n6379 = ndn3_46 & ~ngfdn_3 & n_n7706;
  assign n6380 = ~ndn3_16 & n_n8066 & nen3_16;
  assign n6381 = ~ndn3_32 & ndn3_29 & n_n7710;
  assign n6382 = ~ndn3_40 & n_n7708 & ndn3_39;
  assign n6383 = ~ndn3_21 & n_n7712 & ndn3_19;
  assign n6384 = n_n7711 & ~ndn3_25 & ndn3_22;
  assign n6385 = ndn3_44 & n_n9110 & ~ndn3_46;
  assign n6386 = n_n7763 & ndn3_17 & ~ndn3_18;
  assign n6387 = n_n8760 & ((nen3_22 & ~ndn3_22) | n6899);
  assign n6388 = n_n7668 & ((~ndn3_17 & ndn3_16) | n6900);
  assign n6389 = ndn3_4 & n_n9300 & ~ndn3_7;
  assign n6390 = ~ndn3_12 & ndn3_11 & n_n8276;
  assign n6391 = n_n9505 & ~ndn3_42 & ndn3_40;
  assign n6392 = ndn3_26 & ~ndn3_27 & n_n7684;
  assign n6393 = ndn3_46 & ~ngfdn_3 & n_n7898;
  assign n6394 = n_n8221 & nen3_16 & ~ndn3_16;
  assign n6395 = ~ndn3_32 & ndn3_29 & n_n7666;
  assign n6396 = n_n7664 & ndn3_39 & ~ndn3_40;
  assign n6397 = ~ndn3_21 & n_n8597 & ndn3_19;
  assign n6398 = n_n7667 & ~ndn3_25 & ndn3_22;
  assign n6399 = n_n8628 & ~ndn3_46 & ndn3_44;
  assign n6400 = n_n7687 & ndn3_17 & ~ndn3_18;
  assign n6401 = n_n7803 & (n6908 | (nen3_16 & ~ndn3_16));
  assign n6402 = n_n8116 & ((~ndn3_25 & ndn3_22) | n6909);
  assign n6403 = ndn3_2 & n_n7689 & ~ndn3_4;
  assign n6404 = n_n7682 & nen3_39 & ~ndn3_39;
  assign n6405 = n_n9119 & ~ndn3_9 & ndn3_7;
  assign n6406 = ndn3_46 & n_n9467 & ~ngfdn_3;
  assign n6407 = n_n7688 & ndn3_9 & ~ndn3_11;
  assign n6408 = n_n7686 & ndn3_19 & ~ndn3_21;
  assign n6409 = nen3_28 & ~ndn3_28 & n_n7683;
  assign n6410 = ndn3_44 & n_n8024 & ~ndn3_46;
  assign n6411 = ~ndn3_44 & n_n7681 & ndn3_42;
  assign n6412 = nen3_34 & ~ndn3_34 & n_n8889;
  assign n6413 = n_n7732 & nen3_36 & ~ndn3_36;
  assign n6414 = n_n8153 & ndn3_17 & ~ndn3_18;
  assign n6415 = n_n7685 & nen3_22 & ~ndn3_22;
  assign n6416 = ~ndn3_15 & n_n9257 & ~nsr3_13;
  assign n6417 = n_n8786 & (n6908 | (nen3_16 & ~ndn3_16));
  assign n6418 = n_n8416 & ((~ndn3_25 & ndn3_22) | n6909);
  assign n6419 = ndn3_2 & n_n8739 & ~ndn3_4;
  assign n6420 = n_n6968 & nen3_39 & ~ndn3_39;
  assign n6421 = n_n7866 & ~ndn3_9 & ndn3_7;
  assign n6422 = ndn3_46 & ~ngfdn_3 & n_n8980;
  assign n6423 = n_n7424 & ndn3_9 & ~ndn3_11;
  assign n6424 = n_n9342 & ndn3_19 & ~ndn3_21;
  assign n6425 = n_n9338 & ~ndn3_28 & nen3_28;
  assign n6426 = ndn3_44 & n_n8989 & ~ndn3_46;
  assign n6427 = n_n7920 & ndn3_42 & ~ndn3_44;
  assign n6428 = nen3_34 & ~ndn3_34 & n_n9159;
  assign n6429 = ~ndn3_36 & n_n7831 & nen3_36;
  assign n6430 = n_n8984 & ndn3_17 & ~ndn3_18;
  assign n6431 = n_n7225 & nen3_22 & ~ndn3_22;
  assign n6432 = n_n8833 & ~nsr3_13 & ~ndn3_15;
  assign n6433 = (n7048 | n7049) & (n7055 | n7056);
  assign n6434 = n4966 & ((n5007 & n5008) | (n4969_1 & (~n5007 ^ ~n5008)));
  assign n6435 = n_n8375 & ((nen3_16 & ~ndn3_16) | n6908);
  assign n6436 = n_n7956 & ((~ndn3_25 & ndn3_22) | n6909);
  assign n6437 = ndn3_2 & n_n9023 & ~ndn3_4;
  assign n6438 = ~ndn3_39 & nen3_39 & n_n8095;
  assign n6439 = ndn3_7 & ~ndn3_9 & n_n7955;
  assign n6440 = ndn3_46 & ~ngfdn_3 & n_n7947;
  assign n6441 = ~ndn3_11 & ndn3_9 & n_n7954;
  assign n6442 = n_n9021 & ndn3_19 & ~ndn3_21;
  assign n6443 = nen3_28 & n_n9618 & ~ndn3_28;
  assign n6444 = ndn3_44 & n_n7948 & ~ndn3_46;
  assign n6445 = n_n7949 & ndn3_42 & ~ndn3_44;
  assign n6446 = nen3_34 & n_n8891 & ~ndn3_34;
  assign n6447 = ~ndn3_36 & nen3_36 & n_n7950;
  assign n6448 = ~ndn3_18 & ndn3_17 & n_n7951;
  assign n6449 = n_n8843 & nen3_22 & ~ndn3_22;
  assign n6450 = ~ndn3_15 & n_n7953 & ~nsr3_13;
  assign n6451 = n_n7696 & ((nen3_22 & ~ndn3_22) | n6899);
  assign n6452 = n_n7695 & ((~ndn3_17 & ndn3_16) | n6900);
  assign n6453 = ndn3_4 & ~ndn3_7 & n_n9302;
  assign n6454 = n_n7694 & ndn3_11 & ~ndn3_12;
  assign n6455 = ndn3_40 & ~ndn3_42 & n_n8326;
  assign n6456 = ndn3_26 & ~ndn3_27 & n_n8854;
  assign n6457 = ndn3_46 & ~ngfdn_3 & n_n7691;
  assign n6458 = ~ndn3_16 & nen3_16 & n_n8659;
  assign n6459 = ~ndn3_32 & ndn3_29 & n_n7693;
  assign n6460 = ~ndn3_40 & n_n8410 & ndn3_39;
  assign n6461 = ~ndn3_21 & n_n8599 & ndn3_19;
  assign n6462 = n_n8697 & ~ndn3_25 & ndn3_22;
  assign n6463 = ndn3_44 & n_n9518 & ~ndn3_46;
  assign n6464 = n_n7952 & ndn3_17 & ~ndn3_18;
  assign n6465 = n_n9347 & ((nen3_22 & ~ndn3_22) | n6899);
  assign n6466 = n_n9346 & (n6900 | (~ndn3_17 & ndn3_16));
  assign n6467 = n_n9348 & ~ndn3_7 & ndn3_4;
  assign n6468 = n_n9345 & ndn3_11 & ~ndn3_12;
  assign n6469 = ndn3_40 & n_n9335 & ~ndn3_42;
  assign n6470 = ndn3_26 & n_n9339 & ~ndn3_27;
  assign n6471 = ndn3_46 & ~ngfdn_3 & n_n9333;
  assign n6472 = n_n9344 & nen3_16 & ~ndn3_16;
  assign n6473 = ~ndn3_32 & ndn3_29 & n_n9337;
  assign n6474 = ~ndn3_40 & ndn3_39 & n_n9455;
  assign n6475 = ~ndn3_21 & n_n9341 & ndn3_19;
  assign n6476 = n_n9340 & ~ndn3_25 & ndn3_22;
  assign n6477 = ndn3_44 & n_n9334 & ~ndn3_46;
  assign n6478 = ~ndn3_18 & ndn3_17 & n_n9343;
  assign n6479 = ~preset & n_n9267 & (~ndn3_9 | ndn3_11);
  assign n6480 = ~preset & n4847 & (~n4969_1 ^ ~n4970);
  assign n6481 = n_n9602 & (n6908 | (nen3_16 & ~ndn3_16));
  assign n6482 = n_n9605 & ((~ndn3_25 & ndn3_22) | n6909);
  assign n6483 = n_n9606 & ~ndn3_4 & ndn3_2;
  assign n6484 = n_n9591 & nen3_39 & ~ndn3_39;
  assign n6485 = n_n9604 & ~ndn3_9 & ndn3_7;
  assign n6486 = ndn3_46 & ~ngfdn_3 & n_n9588;
  assign n6487 = n_n9603 & ndn3_9 & ~ndn3_11;
  assign n6488 = ~ndn3_21 & n_n9598 & ndn3_19;
  assign n6489 = nen3_28 & ~ndn3_28 & n_n9595;
  assign n6490 = ndn3_44 & n_n9589 & ~ndn3_46;
  assign n6491 = n_n9590 & ndn3_42 & ~ndn3_44;
  assign n6492 = nen3_34 & ~ndn3_34 & n_n9593;
  assign n6493 = ~ndn3_36 & nen3_36 & n_n9592;
  assign n6494 = n_n9599 & ndn3_17 & ~ndn3_18;
  assign n6495 = n_n9597 & nen3_22 & ~ndn3_22;
  assign n6496 = ~ndn3_15 & n_n9601 & ~nsr3_13;
  assign n6497 = n_n9269 & ((nen3_22 & ~ndn3_22) | n6899);
  assign n6498 = n_n9268 & (n6900 | (~ndn3_17 & ndn3_16));
  assign n6499 = n_n9270 & ~ndn3_7 & ndn3_4;
  assign n6500 = ~ndn3_12 & n_n9267 & ndn3_11;
  assign n6501 = ndn3_40 & n_n9260 & ~ndn3_42;
  assign n6502 = ndn3_26 & n_n9596 & ~ndn3_27;
  assign n6503 = ndn3_46 & ~ngfdn_3 & n_n9259;
  assign n6504 = n_n9266 & nen3_16 & ~ndn3_16;
  assign n6505 = ~ndn3_32 & ndn3_29 & n_n9263;
  assign n6506 = ~ndn3_40 & ndn3_39 & n_n9261;
  assign n6507 = ~ndn3_21 & n_n9265 & ndn3_19;
  assign n6508 = n_n9264 & ~ndn3_25 & ndn3_22;
  assign n6509 = ndn3_44 & n_n9470 & ~ndn3_46;
  assign n6510 = n_n9600 & ndn3_17 & ~ndn3_18;
  assign n6511 = n_n8377 & (n6908 | (nen3_16 & ~ndn3_16));
  assign n6512 = n_n9121 & ((~ndn3_25 & ndn3_22) | n6909);
  assign n6513 = n_n7881 & ~ndn3_4 & ndn3_2;
  assign n6514 = n_n7874 & nen3_39 & ~ndn3_39;
  assign n6515 = n_n7880 & ~ndn3_9 & ndn3_7;
  assign n6516 = ndn3_46 & ~ngfdn_3 & n_n9458;
  assign n6517 = n_n8051 & ndn3_9 & ~ndn3_11;
  assign n6518 = n_n7876 & ndn3_19 & ~ndn3_21;
  assign n6519 = nen3_28 & n_n9000 & ~ndn3_28;
  assign n6520 = ndn3_44 & n_n8609 & ~ndn3_46;
  assign n6521 = ~ndn3_44 & n_n7873 & ndn3_42;
  assign n6522 = nen3_34 & n_n9327 & ~ndn3_34;
  assign n6523 = ~ndn3_36 & nen3_36 & n_n7980;
  assign n6524 = ~ndn3_18 & n_n7877 & ndn3_17;
  assign n6525 = n_n7875 & nen3_22 & ~ndn3_22;
  assign n6526 = n_n7879 & ~nsr3_13 & ~ndn3_15;
  assign n6527 = n4965 & ((n4978 & n4979_1) | (n4972 & (~n4978 ^ ~n4979_1)));
  assign n6528 = (n6922 | n6923) & (n6929 | n6930);
  assign n6529 = n_n9404 & ((nen3_16 & ~ndn3_16) | n6908);
  assign n6530 = n_n9407 & ((~ndn3_25 & ndn3_22) | n6909);
  assign n6531 = ndn3_2 & n_n9408 & ~ndn3_4;
  assign n6532 = n_n9393 & nen3_39 & ~ndn3_39;
  assign n6533 = ndn3_7 & ~ndn3_9 & n_n9406;
  assign n6534 = n_n9390 & ~ngfdn_3 & ndn3_46;
  assign n6535 = n_n9405 & ndn3_9 & ~ndn3_11;
  assign n6536 = ~ndn3_21 & n_n9400 & ndn3_19;
  assign n6537 = nen3_28 & ~ndn3_28 & n_n9397;
  assign n6538 = ndn3_44 & n_n9391 & ~ndn3_46;
  assign n6539 = n_n9392 & ndn3_42 & ~ndn3_44;
  assign n6540 = nen3_34 & n_n9395 & ~ndn3_34;
  assign n6541 = ~ndn3_36 & nen3_36 & n_n9394;
  assign n6542 = ~ndn3_18 & n_n9401 & ndn3_17;
  assign n6543 = ~ndn3_22 & nen3_22 & n_n9399;
  assign n6544 = n_n9403 & ~nsr3_13 & ~ndn3_15;
  assign n6545 = (n6964 | n6965) & (n6971 | n6972);
  assign n6546 = n4973 & ((n4981 & n4982) | (n4955 & (~n4981 ^ ~n4982)));
  assign n6547 = n_n7742 & (n6908 | (nen3_16 & ~ndn3_16));
  assign n6548 = n_n7837 & ((~ndn3_25 & ndn3_22) | n6909);
  assign n6549 = ndn3_2 & ~ndn3_4 & n_n7744;
  assign n6550 = ~ndn3_39 & nen3_39 & n_n7734;
  assign n6551 = ndn3_7 & ~ndn3_9 & n_n8053;
  assign n6552 = n_n8135 & ~ngfdn_3 & ndn3_46;
  assign n6553 = n_n7743 & ndn3_9 & ~ndn3_11;
  assign n6554 = n_n7741 & ndn3_19 & ~ndn3_21;
  assign n6555 = nen3_28 & n_n7738 & ~ndn3_28;
  assign n6556 = ndn3_44 & n_n8247 & ~ndn3_46;
  assign n6557 = ~ndn3_44 & n_n9059 & ndn3_42;
  assign n6558 = nen3_34 & n_n7736 & ~ndn3_34;
  assign n6559 = ~ndn3_36 & n_n7735 & nen3_36;
  assign n6560 = ~ndn3_18 & n_n9141 & ndn3_17;
  assign n6561 = ~ndn3_22 & nen3_22 & n_n7740;
  assign n6562 = ~ndn3_15 & n_n9189 & ~nsr3_13;
  assign n6563 = n_n7655 & ((nen3_16 & ~ndn3_16) | n6908);
  assign n6564 = n_n7657 & ((~ndn3_25 & ndn3_22) | n6909);
  assign n6565 = n_n8770 & ~ndn3_4 & ndn3_2;
  assign n6566 = ~ndn3_39 & nen3_39 & n_n7650;
  assign n6567 = n_n8619 & ~ndn3_9 & ndn3_7;
  assign n6568 = ndn3_46 & ~ngfdn_3 & n_n8862;
  assign n6569 = ~ndn3_11 & ndn3_9 & n_n7656;
  assign n6570 = ~ndn3_21 & n_n7654 & ndn3_19;
  assign n6571 = nen3_28 & ~ndn3_28 & n_n7652;
  assign n6572 = ndn3_44 & ~ndn3_46 & n_n8249;
  assign n6573 = n_n9061 & ndn3_42 & ~ndn3_44;
  assign n6574 = nen3_34 & ~ndn3_34 & n_n9075;
  assign n6575 = ~ndn3_36 & n_n7651 & nen3_36;
  assign n6576 = ~ndn3_18 & ndn3_17 & n_n9015;
  assign n6577 = n_n7653 & nen3_22 & ~ndn3_22;
  assign n6578 = ~ndn3_15 & n_n8260 & ~nsr3_13;
  assign n6579 = n_n8641 & ((nen3_22 & ~ndn3_22) | n6899);
  assign n6580 = n_n9566 & (n6900 | (~ndn3_17 & ndn3_16));
  assign n6581 = n_n7511 & ~ndn3_7 & ndn3_4;
  assign n6582 = n_n8075 & ndn3_11 & ~ndn3_12;
  assign n6583 = ndn3_40 & ~ndn3_42 & n_n8477;
  assign n6584 = ndn3_26 & ~ndn3_27 & n_n7728;
  assign n6585 = n_n8670 & ~ngfdn_3 & ndn3_46;
  assign n6586 = ~ndn3_16 & nen3_16 & n_n8210;
  assign n6587 = n_n8526 & ndn3_29 & ~ndn3_32;
  assign n6588 = ~ndn3_40 & n_n7995 & ndn3_39;
  assign n6589 = n_n7510 & ndn3_19 & ~ndn3_21;
  assign n6590 = n_n9522 & ~ndn3_25 & ndn3_22;
  assign n6591 = ndn3_44 & n_n7670 & ~ndn3_46;
  assign n6592 = n_n7661 & ndn3_17 & ~ndn3_18;
  assign n6593 = n_n9052 & (n6899 | (nen3_22 & ~ndn3_22));
  assign n6594 = n_n9051 & ((~ndn3_17 & ndn3_16) | n6900);
  assign n6595 = n_n9053 & ~ndn3_7 & ndn3_4;
  assign n6596 = n_n9050 & ndn3_11 & ~ndn3_12;
  assign n6597 = ndn3_40 & n_n9043 & ~ndn3_42;
  assign n6598 = ndn3_26 & n_n9368 & ~ndn3_27;
  assign n6599 = ndn3_46 & ~ngfdn_3 & n_n9041;
  assign n6600 = ~ndn3_16 & n_n9049 & nen3_16;
  assign n6601 = ~ndn3_32 & ndn3_29 & n_n9046;
  assign n6602 = ~ndn3_40 & n_n9044 & ndn3_39;
  assign n6603 = n_n9048 & ndn3_19 & ~ndn3_21;
  assign n6604 = n_n9047 & ~ndn3_25 & ndn3_22;
  assign n6605 = ndn3_44 & n_n9042 & ~ndn3_46;
  assign n6606 = n_n9319 & ndn3_17 & ~ndn3_18;
  assign n6607 = n_n9321 & (n6908 | (nen3_16 & ~ndn3_16));
  assign n6608 = n_n9324 & ((~ndn3_25 & ndn3_22) | n6909);
  assign n6609 = ndn3_2 & n_n9325 & ~ndn3_4;
  assign n6610 = ~ndn3_39 & n_n9311 & nen3_39;
  assign n6611 = n_n9323 & ~ndn3_9 & ndn3_7;
  assign n6612 = ndn3_46 & ~ngfdn_3 & n_n9308;
  assign n6613 = n_n9322 & ndn3_9 & ~ndn3_11;
  assign n6614 = n_n9317 & ndn3_19 & ~ndn3_21;
  assign n6615 = nen3_28 & ~ndn3_28 & n_n9315;
  assign n6616 = ndn3_44 & n_n9309 & ~ndn3_46;
  assign n6617 = ~ndn3_44 & n_n9310 & ndn3_42;
  assign n6618 = nen3_34 & ~ndn3_34 & n_n9313;
  assign n6619 = ~ndn3_36 & nen3_36 & n_n9312;
  assign n6620 = n_n9318 & ndn3_17 & ~ndn3_18;
  assign n6621 = n_n9316 & nen3_22 & ~ndn3_22;
  assign n6622 = n_n9320 & ~nsr3_13 & ~ndn3_15;
  assign n6623 = n_n7553 & ((nen3_22 & ~ndn3_22) | n6899);
  assign n6624 = n_n9563 & ((~ndn3_17 & ndn3_16) | n6900);
  assign n6625 = n_n7554 & ~ndn3_7 & ndn3_4;
  assign n6626 = ~ndn3_12 & n_n8298 & ndn3_11;
  assign n6627 = ndn3_40 & ~ndn3_42 & n_n8636;
  assign n6628 = ndn3_26 & ~ndn3_27 & n_n7739;
  assign n6629 = n_n9239 & ~ngfdn_3 & ndn3_46;
  assign n6630 = ~ndn3_16 & nen3_16 & n_n8381;
  assign n6631 = ~ndn3_32 & n_n7552 & ndn3_29;
  assign n6632 = ~ndn3_40 & ndn3_39 & n_n7993;
  assign n6633 = ~ndn3_21 & n_n8035 & ndn3_19;
  assign n6634 = ndn3_22 & n_n8533 & ~ndn3_25;
  assign n6635 = ndn3_44 & n_n8499 & ~ndn3_46;
  assign n6636 = ~ndn3_18 & ndn3_17 & n_n9528;
  assign n6637 = n_n9135 & ((nen3_22 & ~ndn3_22) | n6899);
  assign n6638 = n_n9134 & (n6900 | (~ndn3_17 & ndn3_16));
  assign n6639 = n_n9136 & ~ndn3_7 & ndn3_4;
  assign n6640 = n_n9133 & ndn3_11 & ~ndn3_12;
  assign n6641 = ndn3_40 & n_n9127 & ~ndn3_42;
  assign n6642 = ndn3_26 & n_n9398 & ~ndn3_27;
  assign n6643 = ndn3_46 & ~ngfdn_3 & n_n9125;
  assign n6644 = ~ndn3_16 & nen3_16 & n_n9132;
  assign n6645 = ~ndn3_32 & ndn3_29 & n_n9129;
  assign n6646 = ~ndn3_40 & ndn3_39 & n_n9128;
  assign n6647 = n_n9131 & ndn3_19 & ~ndn3_21;
  assign n6648 = ndn3_22 & n_n9130 & ~ndn3_25;
  assign n6649 = ndn3_44 & ~ndn3_46 & n_n9126;
  assign n6650 = n_n9402 & ndn3_17 & ~ndn3_18;
  assign n6651 = n_n8791 & ((nen3_22 & ~ndn3_22) | n6899);
  assign n6652 = n_n9008 & (n6900 | (~ndn3_17 & ndn3_16));
  assign n6653 = n_n7604 & ~ndn3_7 & ndn3_4;
  assign n6654 = n_n8296 & ndn3_11 & ~ndn3_12;
  assign n6655 = ndn3_40 & n_n7599 & ~ndn3_42;
  assign n6656 = ndn3_26 & n_n7822 & ~ndn3_27;
  assign n6657 = n_n9237 & ~ngfdn_3 & ndn3_46;
  assign n6658 = ~ndn3_16 & nen3_16 & n_n8042;
  assign n6659 = n_n7601 & ndn3_29 & ~ndn3_32;
  assign n6660 = ~ndn3_40 & ndn3_39 & n_n8253;
  assign n6661 = ~ndn3_21 & ndn3_19 & n_n7603;
  assign n6662 = ndn3_22 & ~ndn3_25 & n_n7602;
  assign n6663 = ndn3_44 & n_n7598 & ~ndn3_46;
  assign n6664 = n_n8233 & ndn3_17 & ~ndn3_18;
  assign n6665 = n_n7825 & ((nen3_16 & ~ndn3_16) | n6908);
  assign n6666 = n_n7835 & ((~ndn3_25 & ndn3_22) | n6909);
  assign n6667 = ndn3_2 & ~ndn3_4 & n_n7827;
  assign n6668 = ~ndn3_39 & n_n7819 & nen3_39;
  assign n6669 = ndn3_7 & ~ndn3_9 & n_n7826;
  assign n6670 = ndn3_46 & ~ngfdn_3 & n_n8898;
  assign n6671 = n_n8617 & ndn3_9 & ~ndn3_11;
  assign n6672 = ~ndn3_21 & n_n7823 & ndn3_19;
  assign n6673 = nen3_28 & n_n7821 & ~ndn3_28;
  assign n6674 = ndn3_44 & n_n9036 & ~ndn3_46;
  assign n6675 = n_n9081 & ndn3_42 & ~ndn3_44;
  assign n6676 = nen3_34 & n_n7820 & ~ndn3_34;
  assign n6677 = ~ndn3_36 & nen3_36 & n_n7925;
  assign n6678 = n_n7824 & ndn3_17 & ~ndn3_18;
  assign n6679 = ~ndn3_22 & n_n8699 & nen3_22;
  assign n6680 = n_n9186 & ~nsr3_13 & ~ndn3_15;
  assign n6681 = n_n9499 & ((nen3_16 & ~ndn3_16) | n6908);
  assign n6682 = n_n9502 & ((~ndn3_25 & ndn3_22) | n6909);
  assign n6683 = ndn3_2 & n_n9503 & ~ndn3_4;
  assign n6684 = n_n9488 & nen3_39 & ~ndn3_39;
  assign n6685 = ndn3_7 & ~ndn3_9 & n_n9501;
  assign n6686 = ndn3_46 & n_n9485 & ~ngfdn_3;
  assign n6687 = n_n9500 & ndn3_9 & ~ndn3_11;
  assign n6688 = n_n9495 & ndn3_19 & ~ndn3_21;
  assign n6689 = nen3_28 & n_n9492 & ~ndn3_28;
  assign n6690 = ndn3_44 & n_n9486 & ~ndn3_46;
  assign n6691 = ~ndn3_44 & n_n9487 & ndn3_42;
  assign n6692 = nen3_34 & ~ndn3_34 & n_n9490;
  assign n6693 = ~ndn3_36 & n_n9489 & nen3_36;
  assign n6694 = n_n9496 & ndn3_17 & ~ndn3_18;
  assign n6695 = n_n9494 & nen3_22 & ~ndn3_22;
  assign n6696 = n_n9498 & ~nsr3_13 & ~ndn3_15;
  assign n6697 = n_n9181 & ((nen3_22 & ~ndn3_22) | n6899);
  assign n6698 = n_n9180 & (n6900 | (~ndn3_17 & ndn3_16));
  assign n6699 = ndn3_4 & ~ndn3_7 & n_n9182;
  assign n6700 = n_n9179 & ndn3_11 & ~ndn3_12;
  assign n6701 = ndn3_40 & n_n9172 & ~ndn3_42;
  assign n6702 = ndn3_26 & ~ndn3_27 & n_n9493;
  assign n6703 = ndn3_46 & ~ngfdn_3 & n_n9171;
  assign n6704 = n_n9178 & nen3_16 & ~ndn3_16;
  assign n6705 = ~ndn3_32 & ndn3_29 & n_n9175;
  assign n6706 = ~ndn3_40 & ndn3_39 & n_n9173;
  assign n6707 = n_n9177 & ndn3_19 & ~ndn3_21;
  assign n6708 = n_n9176 & ~ndn3_25 & ndn3_22;
  assign n6709 = ndn3_44 & n_n9473 & ~ndn3_46;
  assign n6710 = n_n9497 & ndn3_17 & ~ndn3_18;
  assign n6711 = n_n8789 & ((nen3_22 & ~ndn3_22) | n6899);
  assign n6712 = n_n8961 & ((~ndn3_17 & ndn3_16) | n6900);
  assign n6713 = ndn3_4 & n_n7643 & ~ndn3_7;
  assign n6714 = n_n7642 & ndn3_11 & ~ndn3_12;
  assign n6715 = ndn3_40 & n_n8328 & ~ndn3_42;
  assign n6716 = ndn3_26 & ~ndn3_27 & n_n8856;
  assign n6717 = n_n8188 & ~ngfdn_3 & ndn3_46;
  assign n6718 = ~ndn3_16 & n_n8661 & nen3_16;
  assign n6719 = ~ndn3_32 & ndn3_29 & n_n7649;
  assign n6720 = ~ndn3_40 & n_n8552 & ndn3_39;
  assign n6721 = n_n8058 & ndn3_19 & ~ndn3_21;
  assign n6722 = n_n7641 & ~ndn3_25 & ndn3_22;
  assign n6723 = ndn3_44 & n_n7640 & ~ndn3_46;
  assign n6724 = n_n7878 & ndn3_17 & ~ndn3_18;
  assign n6725 = ~preset & n_n7726 & (~ndn3_39 | ndn3_40);
  assign n6726 = ~ndn3_40 & ndn3_39 & ~preset & n_n7376;
  assign n6727 = ~preset & n_n9260 & (ndn3_37 | nsr3_37);
  assign n6728 = ~preset & n_n9172 & (ndn3_37 | nsr3_37);
  assign n6729 = nsr3_14 & ~nsr3_13 & n_n8649;
  assign n6730 = nsr3_20 & ndn3_17 & n_n8648;
  assign n6731 = n_n8650 & nsr3_13 & ndn3_12;
  assign n6732 = n_n8796 & ndn3_29 & nsr3_35;
  assign n6733 = nen3_34 & n_n8647 & nsr3_37;
  assign n6734 = ndn3_26 & n_n9242 & nsr3_30;
  assign n6735 = n_n8646 & nsr3_38 & nen3_36;
  assign n6736 = n_n9013 & nsr3_23 & ndn3_19;
  assign n6737 = n_n7629 & ~nsr3_13 & nsr3_14;
  assign n6738 = n_n7628 & ndn3_17 & nsr3_20;
  assign n6739 = n_n7630 & nsr3_13 & ndn3_12;
  assign n6740 = nsr3_35 & n_n8613 & ndn3_29;
  assign n6741 = nen3_34 & n_n8875 & nsr3_37;
  assign n6742 = ndn3_26 & nsr3_30 & n_n8141;
  assign n6743 = n_n7627 & nsr3_38 & nen3_36;
  assign n6744 = ndn3_19 & nsr3_23 & n_n7983;
  assign n6745 = n_n9165 & ~nsr3_13 & nsr3_14;
  assign n6746 = nsr3_20 & ndn3_17 & n_n9164;
  assign n6747 = n_n9166 & nsr3_13 & ndn3_12;
  assign n6748 = n_n9161 & ndn3_29 & nsr3_35;
  assign n6749 = nen3_34 & n_n9160 & nsr3_37;
  assign n6750 = ndn3_26 & nsr3_30 & n_n9162;
  assign n6751 = n_n9578 & nsr3_38 & nen3_36;
  assign n6752 = n_n9163 & nsr3_23 & ndn3_19;
  assign n6753 = nsr3_14 & ~nsr3_13 & n_n8240;
  assign n6754 = nsr3_20 & ndn3_17 & n_n8239;
  assign n6755 = n_n8241 & nsr3_13 & ndn3_12;
  assign n6756 = n_n8312 & ndn3_29 & nsr3_35;
  assign n6757 = nen3_34 & n_n8236 & nsr3_37;
  assign n6758 = ndn3_26 & n_n8237 & nsr3_30;
  assign n6759 = nen3_36 & nsr3_38 & n_n8235;
  assign n6760 = n_n8238 & nsr3_23 & ndn3_19;
  assign n6761 = n_n8574 & ~nsr3_13 & nsr3_14;
  assign n6762 = nsr3_20 & n_n8573 & ndn3_17;
  assign n6763 = n_n8575 & nsr3_13 & ndn3_12;
  assign n6764 = nsr3_35 & ndn3_29 & n_n8572;
  assign n6765 = nen3_34 & n_n8571 & nsr3_37;
  assign n6766 = ndn3_26 & nsr3_30 & n_n8970;
  assign n6767 = n_n8570 & nsr3_38 & nen3_36;
  assign n6768 = ndn3_19 & n_n9150 & nsr3_23;
  assign n6769 = nsr3_14 & n_n9362 & ~nsr3_13;
  assign n6770 = nsr3_20 & ndn3_17 & n_n9552;
  assign n6771 = n_n9363 & nsr3_13 & ndn3_12;
  assign n6772 = n_n9359 & ndn3_29 & nsr3_35;
  assign n6773 = nen3_34 & n_n9358 & nsr3_37;
  assign n6774 = ndn3_26 & nsr3_30 & n_n9360;
  assign n6775 = n_n9357 & nsr3_38 & nen3_36;
  assign n6776 = ndn3_19 & n_n9361 & nsr3_23;
  assign n6777 = n_n9292 & ~nsr3_13 & nsr3_14;
  assign n6778 = nsr3_20 & ndn3_17 & n_n9291;
  assign n6779 = ndn3_12 & n_n9410 & nsr3_13;
  assign n6780 = n_n9289 & ndn3_29 & nsr3_35;
  assign n6781 = nen3_34 & n_n9539 & nsr3_37;
  assign n6782 = ndn3_26 & n_n9290 & nsr3_30;
  assign n6783 = n_n9296 & nsr3_38 & nen3_36;
  assign n6784 = n_n9298 & nsr3_23 & ndn3_19;
  assign n6785 = nsr3_14 & ~nsr3_13 & n_n8273;
  assign n6786 = nsr3_20 & ndn3_17 & n_n8272;
  assign n6787 = ndn3_12 & nsr3_13 & n_n8274;
  assign n6788 = nsr3_35 & ndn3_29 & n_n8348;
  assign n6789 = nen3_34 & n_n8269 & nsr3_37;
  assign n6790 = ndn3_26 & n_n8270 & nsr3_30;
  assign n6791 = nen3_36 & n_n8508 & nsr3_38;
  assign n6792 = n_n8271 & nsr3_23 & ndn3_19;
  assign n6793 = nsr3_14 & n_n9560 & ~nsr3_13;
  assign n6794 = nsr3_20 & ndn3_17 & n_n9559;
  assign n6795 = ndn3_12 & n_n9561 & nsr3_13;
  assign n6796 = n_n9556 & ndn3_29 & nsr3_35;
  assign n6797 = nen3_34 & n_n9555 & nsr3_37;
  assign n6798 = ndn3_26 & n_n9557 & nsr3_30;
  assign n6799 = nen3_36 & n_n9554 & nsr3_38;
  assign n6800 = n_n9558 & nsr3_23 & ndn3_19;
  assign n6801 = nsr3_14 & ~nsr3_13 & n_n9510;
  assign n6802 = nsr3_20 & ndn3_17 & n_n7854;
  assign n6803 = ndn3_12 & n_n8037 & nsr3_13;
  assign n6804 = n_n7852 & ndn3_29 & nsr3_35;
  assign n6805 = nen3_34 & nsr3_37 & n_n8756;
  assign n6806 = ndn3_26 & nsr3_30 & n_n8972;
  assign n6807 = n_n8171 & nsr3_38 & nen3_36;
  assign n6808 = n_n7853 & nsr3_23 & ndn3_19;
  assign n6809 = nsr3_14 & ~nsr3_13 & n_n7771;
  assign n6810 = n_n7770 & ndn3_17 & nsr3_20;
  assign n6811 = n_n7961 & nsr3_13 & ndn3_12;
  assign n6812 = nsr3_35 & ndn3_29 & n_n9331;
  assign n6813 = nen3_34 & n_n7768 & nsr3_37;
  assign n6814 = ndn3_26 & nsr3_30 & n_n7769;
  assign n6815 = nen3_36 & n_n8173 & nsr3_38;
  assign n6816 = n_n8803 & nsr3_23 & ndn3_19;
  assign n6817 = nsr3_14 & n_n8199 & ~nsr3_13;
  assign n6818 = nsr3_20 & n_n9280 & ndn3_17;
  assign n6819 = n_n8200 & nsr3_13 & ndn3_12;
  assign n6820 = n_n8197 & ndn3_29 & nsr3_35;
  assign n6821 = nen3_34 & n_n8710 & nsr3_37;
  assign n6822 = ndn3_26 & nsr3_30 & n_n8366;
  assign n6823 = nen3_36 & n_n8196 & nsr3_38;
  assign n6824 = n_n8198 & nsr3_23 & ndn3_19;
  assign n6825 = n_n9441 & ~nsr3_13 & nsr3_14;
  assign n6826 = nsr3_20 & ndn3_17 & n_n9550;
  assign n6827 = ndn3_12 & n_n9442 & nsr3_13;
  assign n6828 = nsr3_35 & ndn3_29 & n_n9438;
  assign n6829 = nen3_34 & n_n9437 & nsr3_37;
  assign n6830 = ndn3_26 & nsr3_30 & n_n9439;
  assign n6831 = n_n9436 & nsr3_38 & nen3_36;
  assign n6832 = n_n9440 & nsr3_23 & ndn3_19;
  assign n6833 = nsr3_14 & ~nsr3_13 & n_n7584;
  assign n6834 = n_n8447 & ndn3_17 & nsr3_20;
  assign n6835 = n_n8691 & nsr3_13 & ndn3_12;
  assign n6836 = nsr3_35 & ndn3_29 & n_n8968;
  assign n6837 = nen3_34 & n_n7582 & nsr3_37;
  assign n6838 = ndn3_26 & n_n7583 & nsr3_30;
  assign n6839 = n_n8016 & nsr3_38 & nen3_36;
  assign n6840 = n_n7985 & nsr3_23 & ndn3_19;
  assign n6841 = n_n7704 & ~nsr3_13 & nsr3_14;
  assign n6842 = nsr3_20 & ndn3_17 & n_n8685;
  assign n6843 = n_n8577 & nsr3_13 & ndn3_12;
  assign n6844 = n_n9294 & ndn3_29 & nsr3_35;
  assign n6845 = nen3_34 & nsr3_37 & n_n8118;
  assign n6846 = ndn3_26 & n_n7702 & nsr3_30;
  assign n6847 = n_n7701 & nsr3_38 & nen3_36;
  assign n6848 = ndn3_19 & nsr3_23 & n_n7703;
  assign n6849 = nsr3_14 & n_n8531 & ~nsr3_13;
  assign n6850 = nsr3_20 & ndn3_17 & n_n8530;
  assign n6851 = ndn3_12 & nsr3_13 & n_n8615;
  assign n6852 = n_n9275 & ndn3_29 & nsr3_35;
  assign n6853 = nen3_34 & n_n8529 & nsr3_37;
  assign n6854 = ndn3_26 & n_n9244 & nsr3_30;
  assign n6855 = n_n8528 & nsr3_38 & nen3_36;
  assign n6856 = ndn3_19 & nsr3_23 & n_n8935;
  assign n6857 = n6849 | n6850 | n6851 | n6852;
  assign n6858 = n6853 | n6854 | n6855 | n6856;
  assign n6859 = n6753 | n6754 | n6755 | n6756;
  assign n6860 = n6757 | n6758 | n6759 | n6760;
  assign n6861 = n6761 | n6762 | n6763 | n6764;
  assign n6862 = n6765 | n6766 | n6767 | n6768;
  assign n6863 = n6769 | n6770 | n6771 | n6772;
  assign n6864 = n6773 | n6774 | n6775 | n6776;
  assign n6865 = n6833 | n6834 | n6835 | n6836;
  assign n6866 = n6837 | n6838 | n6839 | n6840;
  assign n6867 = n6841 | n6842 | n6843 | n6844;
  assign n6868 = n6845 | n6846 | n6847 | n6848;
  assign n6869 = n6737 | n6738 | n6739 | n6740;
  assign n6870 = n6741 | n6742 | n6743 | n6744;
  assign n6871 = n6809 | n6810 | n6811 | n6812;
  assign n6872 = n6813 | n6814 | n6815 | n6816;
  assign n6873 = n6793 | n6794 | n6795 | n6796;
  assign n6874 = n6797 | n6798 | n6799 | n6800;
  assign n6875 = n6745 | n6746 | n6747 | n6748;
  assign n6876 = n6749 | n6750 | n6751 | n6752;
  assign n6877 = n6729 | n6730 | n6731 | n6732;
  assign n6878 = n6733 | n6734 | n6735 | n6736;
  assign n6879 = n6801 | n6802 | n6803 | n6804;
  assign n6880 = n6805 | n6806 | n6807 | n6808;
  assign n6881 = n6777 | n6778 | n6779 | n6780;
  assign n6882 = n6781 | n6782 | n6783 | n6784;
  assign n6883 = n6825 | n6826 | n6827 | n6828;
  assign n6884 = n6829 | n6830 | n6831 | n6832;
  assign n6885 = n6785 | n6786 | n6787 | n6788;
  assign n6886 = n6789 | n6790 | n6791 | n6792;
  assign n6887 = n6817 | n6818 | n6819 | n6820;
  assign n6888 = n6821 | n6822 | n6823 | n6824;
  assign n6889 = n6857 | n6858 | n6859 | n6860;
  assign n6890 = n6861 | n6862 | n6863 | n6864;
  assign n6891 = n6865 | n6866 | n6867 | n6868;
  assign n6892 = n6869 | n6870 | n6871 | n6872;
  assign n6893 = n6873 | n6874 | n6875 | n6876;
  assign n6894 = n6877 | n6878 | n6879 | n6880;
  assign n6895 = n6881 | n6882 | n6883 | n6884;
  assign n6896 = n6885 | n6886 | n6887 | n6888;
  assign n6897 = n6889 | n6890 | n6891 | n6892;
  assign n6898 = n6893 | n6894 | n6895 | n6896;
  assign n6899 = (~ndn3_9 & ndn3_7) | (ndn3_25 & ~ndn3_26);
  assign n6900 = (ndn3_9 & ~ndn3_11) | (~nsr3_13 & ~ndn3_15);
  assign n6901 = (n_n8779 & n4960) | (n_n7876 & n4961);
  assign n6902 = (n_n7644 & n4958) | (n_n9000 & n4959_1);
  assign n6903 = n6713 | n6714 | n6715 | n6716;
  assign n6904 = n6717 | n6718 | n6719 | n6720;
  assign n6905 = n6721 | n6722 | n6723 | n6724;
  assign n6906 = n6905 | n6711 | n6712;
  assign n6907 = n6901 | n6902 | n6903 | n6904;
  assign n6908 = (~ndn3_19 & nen3_19) | (ndn3_11 & ~ndn3_12);
  assign n6909 = (~ndn3_29 & ndn3_28) | (~ndn3_7 & ndn3_4);
  assign n6910 = (n_n9230 & n4963) | (n_n7878 & n4964_1);
  assign n6911 = n6514 | n6513 | (n_n8856 & n4962);
  assign n6912 = n6515 | n6516 | n6517 | n6518;
  assign n6913 = n6519 | n6520 | n6521 | n6522;
  assign n6914 = n6523 | n6524 | n6525 | n6526;
  assign n6915 = n6914 | n6511 | n6512;
  assign n6916 = n6910 | n6911 | n6912 | n6913;
  assign n6917 = (n_n9491 & n4963) | (n_n9497 & n4964_1);
  assign n6918 = n6684 | n6683 | (n_n9493 & n4962);
  assign n6919 = n6685 | n6686 | n6687 | n6688;
  assign n6920 = n6689 | n6690 | n6691 | n6692;
  assign n6921 = n6693 | n6694 | n6695 | n6696;
  assign n6922 = n6921 | n6681 | n6682;
  assign n6923 = n6917 | n6918 | n6919 | n6920;
  assign n6924 = (n_n9495 & n4961) | (n_n9174 & n4960);
  assign n6925 = (n_n9183 & n4958) | (n_n9492 & n4959_1);
  assign n6926 = n6699 | n6700 | n6701 | n6702;
  assign n6927 = n6703 | n6704 | n6705 | n6706;
  assign n6928 = n6707 | n6708 | n6709 | n6710;
  assign n6929 = n6928 | n6697 | n6698;
  assign n6930 = n6924 | n6925 | n6926 | n6927;
  assign n6931 = (n_n9232 & n4963) | (n_n8233 & n4964_1);
  assign n6932 = n6668 | n6667 | (n_n7822 & n4962);
  assign n6933 = n6669 | n6670 | n6671 | n6672;
  assign n6934 = n6673 | n6674 | n6675 | n6676;
  assign n6935 = n6677 | n6678 | n6679 | n6680;
  assign n6936 = n6935 | n6665 | n6666;
  assign n6937 = n6931 | n6932 | n6933 | n6934;
  assign n6938 = (n_n7600 & n4960) | (n_n7823 & n4961);
  assign n6939 = (n_n7821 & n4959_1) | (n_n8736 & n4958);
  assign n6940 = n6653 | n6654 | n6655 | n6656;
  assign n6941 = n6657 | n6658 | n6659 | n6660;
  assign n6942 = n6661 | n6662 | n6663 | n6664;
  assign n6943 = n6942 | n6651 | n6652;
  assign n6944 = n6938 | n6939 | n6940 | n6941;
  assign n6945 = (n_n9212 & n4960) | (n_n9400 & n4961);
  assign n6946 = (n_n9137 & n4958) | (n_n9397 & n4959_1);
  assign n6947 = n6639 | n6640 | n6641 | n6642;
  assign n6948 = n6643 | n6644 | n6645 | n6646;
  assign n6949 = n6647 | n6648 | n6649 | n6650;
  assign n6950 = n6949 | n6637 | n6638;
  assign n6951 = n6945 | n6946 | n6947 | n6948;
  assign n6952 = (n_n9402 & n4964_1) | (n_n9396 & n4963);
  assign n6953 = n6532 | n6531 | (n_n9398 & n4962);
  assign n6954 = n6533 | n6534 | n6535 | n6536;
  assign n6955 = n6537 | n6538 | n6539 | n6540;
  assign n6956 = n6541 | n6542 | n6543 | n6544;
  assign n6957 = n6956 | n6529 | n6530;
  assign n6958 = n6952 | n6953 | n6954 | n6955;
  assign n6959 = (n_n7741 & n4961) | (n_n8638 & n4960);
  assign n6960 = (n_n8009 & n4958) | (n_n7738 & n4959_1);
  assign n6961 = n6625 | n6626 | n6627 | n6628;
  assign n6962 = n6629 | n6630 | n6631 | n6632;
  assign n6963 = n6633 | n6634 | n6635 | n6636;
  assign n6964 = n6963 | n6623 | n6624;
  assign n6965 = n6959 | n6960 | n6961 | n6962;
  assign n6966 = (n_n7737 & n4963) | (n_n9528 & n4964_1);
  assign n6967 = n6550 | n6549 | (n_n7739 & n4962);
  assign n6968 = n6551 | n6552 | n6553 | n6554;
  assign n6969 = n6555 | n6556 | n6557 | n6558;
  assign n6970 = n6559 | n6560 | n6561 | n6562;
  assign n6971 = n6970 | n6547 | n6548;
  assign n6972 = n6966 | n6967 | n6968 | n6969;
  assign n6973 = (n_n9317 & n4961) | (n_n9045 & n4960);
  assign n6974 = (n_n9315 & n4959_1) | (n_n9054 & n4958);
  assign n6975 = n6595 | n6596 | n6597 | n6598;
  assign n6976 = n6599 | n6600 | n6601 | n6602;
  assign n6977 = n6603 | n6604 | n6605 | n6606;
  assign n6978 = n6977 | n6593 | n6594;
  assign n6979 = n6973 | n6974 | n6975 | n6976;
  assign n6980 = (n_n9314 & n4963) | (n_n9319 & n4964_1);
  assign n6981 = n6610 | n6609 | (n_n9368 & n4962);
  assign n6982 = n6611 | n6612 | n6613 | n6614;
  assign n6983 = n6615 | n6616 | n6617 | n6618;
  assign n6984 = n6619 | n6620 | n6621 | n6622;
  assign n6985 = n6984 | n6607 | n6608;
  assign n6986 = n6980 | n6981 | n6982 | n6983;
  assign n6987 = (n_n7509 & n4960) | (n_n7654 & n4961);
  assign n6988 = (n_n8011 & n4958) | (n_n7652 & n4959_1);
  assign n6989 = n6581 | n6582 | n6583 | n6584;
  assign n6990 = n6585 | n6586 | n6587 | n6588;
  assign n6991 = n6589 | n6590 | n6591 | n6592;
  assign n6992 = n6991 | n6579 | n6580;
  assign n6993 = n6987 | n6988 | n6989 | n6990;
  assign n6994 = (n_n8033 & n4963) | (n_n7661 & n4964_1);
  assign n6995 = n6566 | n6565 | (n_n7728 & n4962);
  assign n6996 = n6567 | n6568 | n6569 | n6570;
  assign n6997 = n6571 | n6572 | n6573 | n6574;
  assign n6998 = n6575 | n6576 | n6577 | n6578;
  assign n6999 = n6998 | n6563 | n6564;
  assign n7000 = n6994 | n6995 | n6996 | n6997;
  assign n7001 = (n_n9262 & n4960) | (n_n9598 & n4961);
  assign n7002 = (n_n9595 & n4959_1) | (n_n9271 & n4958);
  assign n7003 = n6499 | n6500 | n6501 | n6502;
  assign n7004 = n6503 | n6504 | n6505 | n6506;
  assign n7005 = n6507 | n6508 | n6509 | n6510;
  assign n7006 = n7005 | n6497 | n6498;
  assign n7007 = n7001 | n7002 | n7003 | n7004;
  assign n7008 = (n_n9594 & n4963) | (n_n9600 & n4964_1);
  assign n7009 = n6484 | n6483 | (n_n9596 & n4962);
  assign n7010 = n6485 | n6486 | n6487 | n6488;
  assign n7011 = n6489 | n6490 | n6491 | n6492;
  assign n7012 = n6493 | n6494 | n6495 | n6496;
  assign n7013 = n7012 | n6481 | n6482;
  assign n7014 = n7008 | n7009 | n7010 | n7011;
  assign n7015 = (n_n7686 & n4961) | (n_n7665 & n4960);
  assign n7016 = (n_n7683 & n4959_1) | (n_n8110 & n4958);
  assign n7017 = n6389 | n6390 | n6391 | n6392;
  assign n7018 = n6393 | n6394 | n6395 | n6396;
  assign n7019 = n6397 | n6398 | n6399 | n6400;
  assign n7020 = n7019 | n6387 | n6388;
  assign n7021 = n7015 | n7016 | n7017 | n7018;
  assign n7022 = (n_n8586 & n4963) | (n_n7687 & n4964_1);
  assign n7023 = n6404 | n6403 | (n_n7684 & n4962);
  assign n7024 = n6405 | n6406 | n6407 | n6408;
  assign n7025 = n6409 | n6410 | n6411 | n6412;
  assign n7026 = n6413 | n6414 | n6415 | n6416;
  assign n7027 = n7026 | n6401 | n6402;
  assign n7028 = n7022 | n7023 | n7024 | n7025;
  assign n7029 = (n_n9342 & n4961) | (n_n9336 & n4960);
  assign n7030 = (n_n9338 & n4959_1) | (n_n9349 & n4958);
  assign n7031 = n6467 | n6468 | n6469 | n6470;
  assign n7032 = n6471 | n6472 | n6473 | n6474;
  assign n7033 = n6475 | n6476 | n6477 | n6478;
  assign n7034 = n7033 | n6465 | n6466;
  assign n7035 = n7029 | n7030 | n7031 | n7032;
  assign n7036 = (n_n6976 & n4963) | (n_n9343 & n4964_1);
  assign n7037 = n6420 | n6419 | (n_n9339 & n4962);
  assign n7038 = n6421 | n6422 | n6423 | n6424;
  assign n7039 = n6425 | n6426 | n6427 | n6428;
  assign n7040 = n6429 | n6430 | n6431 | n6432;
  assign n7041 = n7040 | n6417 | n6418;
  assign n7042 = n7036 | n7037 | n7038 | n7039;
  assign n7043 = (n_n9021 & n4961) | (n_n7692 & n4960);
  assign n7044 = (n_n7697 & n4958) | (n_n9618 & n4959_1);
  assign n7045 = n6453 | n6454 | n6455 | n6456;
  assign n7046 = n6457 | n6458 | n6459 | n6460;
  assign n7047 = n6461 | n6462 | n6463 | n6464;
  assign n7048 = n7047 | n6451 | n6452;
  assign n7049 = n7043 | n7044 | n7045 | n7046;
  assign n7050 = (n_n8966 & n4963) | (n_n7952 & n4964_1);
  assign n7051 = n6438 | n6437 | (n_n8854 & n4962);
  assign n7052 = n6439 | n6440 | n6441 | n6442;
  assign n7053 = n6443 | n6444 | n6445 | n6446;
  assign n7054 = n6447 | n6448 | n6449 | n6450;
  assign n7055 = n7054 | n6435 | n6436;
  assign n7056 = n7050 | n7051 | n7052 | n7053;
  assign n7057 = (n_n7762 & n4961) | (n_n7709 & n4960);
  assign n7058 = (n_n8852 & n4959_1) | (n_n8986 & n4958);
  assign n7059 = n6375 | n6376 | n6377 | n6378;
  assign n7060 = n6379 | n6380 | n6381 | n6382;
  assign n7061 = n6383 | n6384 | n6385 | n6386;
  assign n7062 = n7061 | n6373 | n6374;
  assign n7063 = n7057 | n7058 | n7059 | n7060;
  assign n7064 = (n_n7763 & n4964_1) | (n_n7759 & n4963);
  assign n7065 = n6360 | n6359 | (n_n7760 & n4962);
  assign n7066 = n6361 | n6362 | n6363 | n6364;
  assign n7067 = n6365 | n6366 | n6367 | n6368;
  assign n7068 = n6369 | n6370 | n6371 | n6372;
  assign n7069 = n7068 | n6357 | n6358;
  assign n7070 = n7064 | n7065 | n7066 | n7067;
  assign n7071 = (n_n8408 & n4963) | (n_n7811 & n4964_1);
  assign n7072 = n6325 | n6324 | (n_n7809 & n4962);
  assign n7073 = n6326 | n6327 | n6328 | n6329;
  assign n7074 = n6330 | n6331 | n6332 | n6333;
  assign n7075 = n6334 | n6335 | n6336 | n6337;
  assign n7076 = n7075 | n6322 | n6323;
  assign n7077 = n7071 | n7072 | n7073 | n7074;
  assign n7078 = (n_n8088 & n4960) | (n_n7810 & n4961);
  assign n7079 = (n_n8108 & n4958) | (n_n8473 & n4959_1);
  assign n7080 = n6340 | n6341 | n6342 | n6343;
  assign n7081 = n6344 | n6345 | n6346 | n6347;
  assign n7082 = n6348 | n6349 | n6350 | n6351;
  assign n7083 = n7082 | n6338 | n6339;
  assign n7084 = n7078 | n7079 | n7080 | n7081;
  assign n7085 = n_n9248 & ~n_n7306;
  assign n7086 = (nsr3_38 & nen3_36) | (nsr3_23 & ndn3_19);
  assign n7087 = (nsr3_37 & nen3_34) | (nsr3_30 & ndn3_26);
  assign n7088 = (ndn3_29 & nsr3_35) | (ndn3_17 & nsr3_20);
  assign n7089 = n4974_1 & n_n9198;
  assign n7090 = n6305 | n6303 | n6304;
  assign n7091 = n6306 | n6307 | n6308 | n6309;
  assign n7092 = n6298 | n6296 | n6297;
  assign n7093 = n6299 | n6300 | n6301 | n6302;
  assign n7094 = n6284 | n6282 | n6283;
  assign n7095 = n6285 | n6286 | n6287 | n6288;
  assign n7096 = n6263 | n6261 | n6262;
  assign n7097 = n6264 | n6265 | n6266 | n6267;
  assign n7098 = n6256 | n6254 | n6255;
  assign n7099 = n6257 | n6258 | n6259 | n6260;
  assign n7100 = n6235 | n6233 | n6234;
  assign n7101 = n6236 | n6237 | n6238 | n6239;
  assign n7102 = n6242 | n6240 | n6241;
  assign n7103 = n6243 | n6244 | n6245 | n6246;
  assign n7104 = n6228 | n6226 | n6227;
  assign n7105 = n6229 | n6230 | n6231 | n6232;
  assign n7106 = n6249 | n6247 | n6248;
  assign n7107 = n6250 | n6251 | n6252 | n6253;
  assign n7108 = n6270 | n6268 | n6269;
  assign n7109 = n6271 | n6272 | n6273 | n6274;
  assign n7110 = n6277 | n6275 | n6276;
  assign n7111 = n6278 | n6279 | n6280 | n6281;
  assign n7112 = n6221 | n6219 | n6220;
  assign n7113 = n6222 | n6223 | n6224 | n6225;
  assign n7114 = n6291 | n6289 | n6290;
  assign n7115 = n6292 | n6293 | n6294 | n6295;
  assign n7116 = n6214 | n6212 | n6213;
  assign n7117 = n6215 | n6216 | n6217 | n6218;
  assign n7118 = n6207 | n6205 | n6206;
  assign n7119 = n6208 | n6209 | n6210 | n6211;
  assign n7120 = n6201 | n6202 | n6203 | n6204;
  assign n7121 = n5001 & ~n_n8557 & n4856;
  assign n7122 = n4856 & n_n8557;
  assign n7123 = n_n9638 & n4856 & (n7094 | n7095);
  assign n7124 = (n_n9225 & n4960) | (n_n7888 & n4961);
  assign n7125 = (n_n7887 & n4959_1) | (n_n7850 & n4958);
  assign n7126 = n6165 | n6166 | n6167 | n6168;
  assign n7127 = n6169 | n6170 | n6171 | n6172;
  assign n7128 = n6173 | n6174 | n6175 | n6176;
  assign n7129 = n7128 | n6163 | n6164;
  assign n7130 = n7124 | n7125 | n7126 | n7127;
  assign n7131 = (n_n7886 & n4963) | (n_n7889 & n4964_1);
  assign n7132 = n6150 | n6149 | (n_n9520 & n4962);
  assign n7133 = n6151 | n6152 | n6153 | n6154;
  assign n7134 = n6155 | n6156 | n6157 | n6158;
  assign n7135 = n6159 | n6160 | n6161 | n6162;
  assign n7136 = n7135 | n6147 | n6148;
  assign n7137 = n7131 | n7132 | n7133 | n7134;
  assign n7138 = (n_n8519 & n4964_1) | (n_n8002 & n4963);
  assign n7139 = n6132 | n6131 | (n_n8004 & n4962);
  assign n7140 = n6133 | n6134 | n6135 | n6136;
  assign n7141 = n6137 | n6138 | n6139 | n6140;
  assign n7142 = n6141 | n6142 | n6143 | n6144;
  assign n7143 = n7142 | n6129 | n6130;
  assign n7144 = n7138 | n7139 | n7140 | n7141;
  assign n7145 = (n_n8005 & n4961) | (n_n9223 & n4960);
  assign n7146 = (n_n8003 & n4959_1) | (n_n8482 & n4958);
  assign n7147 = n6117 | n6118 | n6119 | n6120;
  assign n7148 = n6121 | n6122 | n6123 | n6124;
  assign n7149 = n6125 | n6126 | n6127 | n6128;
  assign n7150 = n7149 | n6115 | n6116;
  assign n7151 = n7145 | n7146 | n7147 | n7148;
  assign n7152 = (n_n8139 & n4960) | (n_n7933 & n4961);
  assign n7153 = (n_n8000 & n4958) | (n_n7931 & n4959_1);
  assign n7154 = n6087 | n6088 | n6089_1 | n6090;
  assign n7155 = n6091 | n6092 | n6093 | n6094_1;
  assign n7156 = n6095 | n6096 | n6097 | n6098;
  assign n7157 = n7156 | n6085 | n6086;
  assign n7158 = n7152 | n7153 | n7154 | n7155;
  assign n7159 = (n_n8106 & n4964_1) | (n_n7930 & n4963);
  assign n7160 = n6102 | n6101 | (n_n7932 & n4962);
  assign n7161 = n6103 | n6104 | n6105 | n6106;
  assign n7162 = n6107 | n6108 | n6109 | n6110;
  assign n7163 = n6111 | n6112 | n6113 | n6114;
  assign n7164 = n7163 | n6099 | n6100;
  assign n7165 = n7159 | n7160 | n7161 | n7162;
  assign n7166 = ~n_n8869 & ~n_n8603 & ~n_n8798;
  assign n7167 = ~n4924_1 & n4953 & (n_n8933 ^ n5000);
  assign n7168 = n7166 & (n_n8911 ^ (n_n8933 | n5000));
  assign n7169 = ~n4927 & n7167;
  assign n7170 = ~n4928 & n7168 & (~n_n8993 ^ ~n5005);
  assign n7171 = ~n4943 & n7169 & (~n_n8561 ^ ~n4999_1);
  assign n7172 = ~n4947 & n7171;
  assign n7173 = ~n4899_1 & n7170 & (~n_n8913 ^ ~n4968);
  assign n7174 = preset | ~n_n9198 | ~n4967 | ~n4974_1;
  assign n7175 = n_n9434 & n4856 & (n7096 | n7097);
  assign n7176 = ~n4967 & ~preset;
  assign n7177 = pdn | preset | (nsr3_23 & ~nak3_13);
  assign n7178 = pdn | preset | (nsr3_13 & ~nak3_13);
  assign n7179 = pdn | preset | (nsr3_38 & ~nak3_13);
  assign n7180 = n_n8549 & n4856 & (n7090 | n7091);
  assign n7181 = n4856 & (n_n8652 ? ~n4910 : (n4910 & n5001));
  assign n7182 = ~n_n8707 & (n4911 ^ (n7104 | n7105));
  assign n7183 = n_n8707 & n4856 & (~n4911 ^ n4913);
  assign n7184 = n7183 | (n4856 & n5001 & n7182);
  assign n7185 = pdn | preset | (nsr3_30 & ~ndn3_26);
  assign n7186 = n_n8354 & n4856 & (n7116 | n7117);
  assign n7187 = n_n9512 & n4856 & (n7098 | n7099);
  assign n7188 = n5001 & n4856 & n4920;
  assign n7189 = n4856 & n_n9512;
  assign n7190 = n5626 | (~preset & n_n9512 & ~n5001);
  assign n7191 = pdn | preset | (nsr3_35 & ~nak3_13);
  assign n7192 = n_n9416 & n4856 & (n7108 | n7109);
  assign n7193 = pdn | (~nak3_13 & (preset | nsr3_14));
  assign n7194 = ~n_n8603 & ~n5975 & (~n4975 | ~n7176);
  assign n7195 = ~n6866 & ~n_n8603 & ~n6865;
  assign n7196 = ~n4856 & n_n8603;
  assign n7197 = ~n4898 & (n7194 | n7195);
  assign n7198 = n4974_1 & n4967 & ~preset & n_n9198;
  assign n7199 = n_n8449 & n4856 & (n7092 | n7093);
  assign n7200 = n_n9448 & n4856 & (n7114 | n7115);
  assign n7201 = n_n9537 & n4856 & (n7110 | n7111);
  assign n7202 = n_n8929 & ~preset;
  assign n7203 = ~preset & (n6897 | n6898);
  assign n7204 = ~n_n9284 & (n4909_1 ^ (n7102 | n7103));
  assign n7205 = n_n9284 & n4856 & (~n4909_1 ^ n4936);
  assign n7206 = n7205 | (n4856 & n5001 & n7204);
  assign n7207 = n_n8821 & n4856 & (n7112 | n7113);
  assign n7208 = ~n_n9353 & (n4912 ^ (n7106 | n7107));
  assign n7209 = n_n9353 & n4856 & (~n4912 ^ n4938);
  assign n7210 = pdn | preset | (nsr3_37 & ~nen3_34);
  assign n7211 = pdn | preset | (~nak3_13 & nsr3_20);
  assign n7212 = n_n8419 & n4856 & (n7118 | n7119);
  always @ (posedge clk) begin
    n_n9280 <= n491;
    n_n9172 <= n496;
    n_n9260 <= n501;
    n_n7726 <= n506;
    n_n8270 <= n511;
    n_n8196 <= n516;
    n_n9150 <= n521;
    n_n9267 <= n526;
    n_n7779 <= n531;
    n_n9503 <= n536;
    n_n8150 <= n541;
    n_n9401 <= n546;
    n_n7341 <= n551;
    n_n9180 <= n556;
    n_n8592 <= n561;
    n_n8871 <= n566;
    n_n7252 <= n571;
    n_n7271 <= n576;
    n_n6991 <= n581;
    n_n8557 <= n586;
    n_n7707 <= n591;
    n_n7552 <= n596;
    ndn3_23 <= n601;
    n_n9548 <= n606;
    n_n9467 <= n611;
    n_n8002 <= n616;
    n_n6950 <= n621;
    n_n8930 <= n626;
    n_n7244 <= n631;
    n_n7819 <= n636;
    n_n8883 <= n641;
    n_n7709 <= n646;
    n_n9580 <= n651;
    n_n9130 <= n656;
    n_n9486 <= n661;
    n_n9235 <= n666;
    n_n7522 <= n671;
    n_n7373 <= n676;
    n_n9085 <= n681;
    n_n9638 <= n686;
    n_n7452 <= n691;
    n_n8775 <= n696;
    n_n7654 <= n701;
    n_n8410 <= n706;
    n_n8208 <= n711;
    n_n8377 <= n716;
    n_n7558 <= n721;
    n_n7599 <= n726;
    n_n8225 <= n731;
    n_n8202 <= n736;
    n_n7670 <= n741;
    n_n7888 <= n746;
    n_n7889 <= n751;
    n_n8597 <= n756;
    n_n8152 <= n761;
    n_n8394 <= n766;
    n_n7812 <= n771;
    n_n7816 <= n776;
    n_n9141 <= n781;
    n_n7332 <= n786;
    n_n8758 <= n791;
    n_n7765 <= n796;
    n_n7877 <= n801;
    n_n7814 <= n806;
    n_n9008 <= n811;
    n_n7581 <= n816;
    n_n7376 <= n821;
    n_n7970 <= n826;
    pover_0_0_ <= n831;
    n_n8599 <= n835;
    n_n8227 <= n840;
    n_n9442 <= n845;
    n_n9485 <= n850;
    n_n7148 <= n855;
    n_n9311 <= n860;
    n_n9273 <= n865;
    ndn3_9 <= n870;
    n_n8613 <= n875;
    n_n8533 <= n880;
    n_n8699 <= n885;
    n_n8609 <= n890;
    n_n8308 <= n895;
    n_n8655 <= n900;
    n_n8981 <= n905;
    n_n7583 <= n910;
    n_n9198 <= n915;
    n_n9602 <= n920;
    n_n8786 <= n925;
    n_n9598 <= n930;
    n_n7738 <= n935;
    n_n8573 <= n940;
    n_n9473 <= n945;
    n_n9000 <= n950;
    n_n8001 <= n955;
    n_n9554 <= n960;
    n_n8508 <= n965;
    n_n9635 <= n970;
    n_n7190 <= n975;
    n_n8702 <= n980;
    n_n9106 <= n985;
    n_n7409 <= n990;
    n_n9437 <= n995;
    n_n9052 <= n1000;
    n_n8647 <= n1005;
    n_n9265 <= n1010;
    n_n7179 <= n1015;
    ndn3_13 <= n1020;
    ndn3_17 <= n1025;
    ndn3_25 <= n1030;
    ndn3_29 <= n1035;
    n_n9539 <= n1040;
    n_n7953 <= n1045;
    n_n8488 <= n1050;
    nen3_22 <= n1055;
    n_n9438 <= n1060;
    n_n8132 <= n1065;
    n_n8661 <= n1070;
    n_n7759 <= n1075;
    n_n8333 <= n1080;
    n_n9399 <= n1085;
    n_n7798 <= n1090;
    n_n9434 <= n1095;
    n_n7910 <= n1100;
    n_n9528 <= n1105;
    n_n7850 <= n1110;
    n_n8251 <= n1115;
    n_n7937 <= n1120;
    n_n8482 <= n1125;
    n_n9290 <= n1130;
    n_n8007 <= n1135;
    n_n7556 <= n1140;
    n_n9064 <= n1145;
    n_n9398 <= n1150;
    n_n9412 <= n1155;
    n_n9361 <= n1160;
    n_n9304 <= n1165;
    n_n7651 <= n1170;
    n_n7712 <= n1175;
    n_n7735 <= n1180;
    n_n7934 <= n1185;
    n_n7811 <= n1190;
    n_n8053 <= n1195;
    n_n9015 <= n1200;
    n_n8066 <= n1205;
    n_n9518 <= n1210;
    n_n8091 <= n1215;
    n_n9257 <= n1220;
    n_n8175 <= n1225;
    n_n8491 <= n1230;
    n_n8114 <= n1235;
    n_n7951 <= n1240;
    n_n8913 <= n1245;
    n_n8035 <= n1250;
    n_n8631 <= n1255;
    n_n8243 <= n1260;
    n_n7857 <= n1265;
    ngfdn_3 <= n1270;
    n_n7791 <= n1275;
    n_n9175 <= n1280;
    n_n9588 <= n1285;
    n_n9049 <= n1290;
    n_n9483 <= n1295;
    n_n9410 <= n1300;
    n_n7691 <= n1305;
    n_n7740 <= n1310;
    n_n7602 <= n1315;
    n_n7783 <= n1320;
    n_n7948 <= n1325;
    n_n7054 <= n1330;
    n_n9343 <= n1335;
    n_n9400 <= n1340;
    nsr1_2 <= n1345;
    n_n9127 <= n1350;
    n_n8531 <= n1355;
    n_n9335 <= n1360;
    n_n7324 <= n1365;
    n_n9611 <= n1370;
    n_n8112 <= n1375;
    n_n9406 <= n1380;
    n_n9618 <= n1385;
    n_n9613 <= n1390;
    n_n9242 <= n1395;
    n_n7384 <= n1400;
    n_n8884 <= n1405;
    n_n7462 <= n1410;
    n_n7908 <= n1415;
    n_n8765 <= n1420;
    n_n7909 <= n1425;
    n_n7898 <= n1430;
    n_n9135 <= n1435;
    n_n8862 <= n1440;
    n_n8037 <= n1445;
    ndn3_18 <= n1450;
    ndn3_22 <= n1455;
    n_n8974 <= n1460;
    n_n7286 <= n1465;
    n_n9223 <= n1470;
    n_n7306 <= n1475;
    n_n9169 <= n1480;
    n_n9125 <= n1485;
    nen3_39 <= n1490;
    n_n8278 <= n1495;
    n_n9557 <= n1500;
    n_n7758 <= n1505;
    n_n9391 <= n1510;
    n_n8110 <= n1515;
    n_n9597 <= n1520;
    n_n8568 <= n1525;
    n_n7428 <= n1530;
    n_n7931 <= n1535;
    n_n7742 <= n1540;
    n_n7236 <= n1545;
    n_n8219 <= n1550;
    n_n9568 <= n1555;
    n_n9200 <= n1560;
    n_n8545 <= n1565;
    n_n7823 <= n1570;
    n_n8005 <= n1575;
    n_n8736 <= n1580;
    n_n9339 <= n1585;
    n_n8499 <= n1590;
    n_n8086 <= n1595;
    n_n7803 <= n1600;
    n_n7640 <= n1605;
    n_n9098 <= n1610;
    n_n7160 <= n1615;
    n_n7713 <= n1620;
    n_n9566 <= n1625;
    n_n7955 <= n1630;
    n_n8414 <= n1635;
    n_n8006 <= n1640;
    n_n9560 <= n1645;
    n_n8742 <= n1650;
    n_n7174 <= n1655;
    n_n8882 <= n1660;
    n_n7546 <= n1665;
    n_n8282 <= n1670;
    n_n8998 <= n1675;
    n_n7656 <= n1680;
    n_n9465 <= n1685;
    n_n9601 <= n1690;
    n_n8875 <= n1695;
    n_n7954 <= n1700;
    n_n8959 <= n1705;
    n_n8957 <= n1710;
    n_n8247 <= n1715;
    n_n8258 <= n1720;
    n_n7641 <= n1725;
    n_n8843 <= n1730;
    n_n9321 <= n1735;
    n_n7702 <= n1740;
    nsr3_23 <= n1745;
    n_n8199 <= n1750;
    n_n7983 <= n1755;
    n_n7217 <= n1760;
    n_n7821 <= n1765;
    n_n9489 <= n1770;
    n_n8348 <= n1775;
    n_n9408 <= n1780;
    n_n8445 <= n1785;
    n_n9501 <= n1790;
    n_n7831 <= n1795;
    n_n7757 <= n1800;
    n_n9174 <= n1805;
    n_n9432 <= n1810;
    n_n8678 <= n1815;
    n_n8024 <= n1820;
    n_n7806 <= n1825;
    n_n8996 <= n1830;
    n_n7918 <= n1835;
    n_n8260 <= n1840;
    n_n9341 <= n1845;
    n_n9189 <= n1850;
    n_n9096 <= n1855;
    ndn3_30 <= n1860;
    n_n7775 <= n1865;
    n_n7693 <= n1870;
    nen3_16 <= n1875;
    n_n7643 <= n1880;
    n_n8941 <= n1885;
    n_n8042 <= n1890;
    n_n8681 <= n1895;
    n_n8659 <= n1900;
    n_n9110 <= n1905;
    n_n9573 <= n1910;
    n_n8951 <= n1915;
    n_n9589 <= n1920;
    n_n9387 <= n1925;
    n_n8279 <= n1930;
    n_n7790 <= n1935;
    n_n8406 <= n1940;
    n_n8582 <= n1945;
    n_n7911 <= n1950;
    n_n7474 <= n1955;
    n_n8466 <= n1960;
    n_n6984 <= n1965;
    n_n7760 <= n1970;
    n_n7847 <= n1975;
    n_n9559 <= n1980;
    n_n7362 <= n1985;
    n_n9300 <= n1990;
    n_n9550 <= n1995;
    n_n9492 <= n2000;
    n_n8777 <= n2005;
    n_n7764 <= n2010;
    n_n7826 <= n2015;
    n_n7777 <= n2020;
    n_n7824 <= n2025;
    n_n8173 <= n2030;
    n_n7498 <= n2035;
    n_n9148 <= n2040;
    n_n8753 <= n2045;
    n_n8772 <= n2050;
    n_n8049 <= n2055;
    n_n9362 <= n2060;
    ndn1_4 <= n2065;
    n_n9561 <= n2070;
    n_n9004 <= n2075;
    n_n8203 <= n2080;
    n_n8153 <= n2085;
    n_n9263 <= n2090;
    n_n8369 <= n2095;
    n_n9331 <= n2100;
    n_n7454 <= n2105;
    ndn3_7 <= n2110;
    n_n7527 <= n2115;
    n_n9036 <= n2120;
    n_n7875 <= n2125;
    n_n8697 <= n2130;
    n_n9497 <= n2135;
    n_n7291 <= n2140;
    nsr3_13 <= n2145;
    nsr3_38 <= n2150;
    n_n8240 <= n2155;
    n_n7703 <= n2160;
    n_n9282 <= n2165;
    n_n8237 <= n2170;
    n_n8935 <= n2175;
    n_n9244 <= n2180;
    n_n8648 <= n2185;
    n_n8235 <= n2190;
    n_n8611 <= n2195;
    n_n9045 <= n2200;
    n_n9334 <= n2205;
    n_n8572 <= n2210;
    n_n9491 <= n2215;
    n_n9134 <= n2220;
    n_n9555 <= n2225;
    n_n9336 <= n2230;
    n_n7050 <= n2235;
    n_n9346 <= n2240;
    n_n7140 <= n2245;
    n_n7681 <= n2250;
    n_n6948 <= n2255;
    n_n8549 <= n2260;
    ndn3_19 <= n2265;
    ndn3_28 <= n2270;
    n_n7102 <= n2275;
    n_n8093 <= n2280;
    n_n9041 <= n2285;
    n_n8381 <= n2290;
    n_n8810 <= n2295;
    nen3_36 <= n2300;
    n_n9047 <= n2305;
    n_n9333 <= n2310;
    n_n7736 <= n2315;
    n_n7820 <= n2320;
    n_n8986 <= n2325;
    n_n8891 <= n2330;
    n_n8000 <= n2335;
    n_n7968 <= n2340;
    n_n8750 <= n2345;
    n_n9558 <= n2350;
    n_n9368 <= n2355;
    n_n8519 <= n2360;
    n_n6956 <= n2365;
    n_n8298 <= n2370;
    n_n9397 <= n2375;
    n_n7017 <= n2380;
    n_n8638 <= n2385;
    n_n9552 <= n2390;
    n_n8964 <= n2395;
    n_n8016 <= n2400;
    n_n7603 <= n2405;
    n_n7696 <= n2410;
    n_n8589 <= n2415;
    n_n9337 <= n2420;
    n_n9132 <= n2425;
    n_n8652 <= n2430;
    n_n8707 <= n2435;
    n_n9407 <= n2440;
    n_n9044 <= n2445;
    n_n8808 <= n2450;
    nsr3_30 <= n2455;
    n_n8274 <= n2460;
    n_n8615 <= n2465;
    n_n8238 <= n2470;
    n_n7854 <= n2475;
    n_n8649 <= n2480;
    n_n8236 <= n2485;
    n_n8269 <= n2490;
    n_n9592 <= n2495;
    n_n8022 <= n2500;
    n_n8744 <= n2505;
    n_n8529 <= n2510;
    n_n7967 <= n2515;
    n_n9487 <= n2520;
    n_n8685 <= n2525;
    n_n9531 <= n2530;
    n_n9510 <= n2535;
    n_n7771 <= n2540;
    n_n8480 <= n2545;
    n_n8543 <= n2550;
    n_n7789 <= n2555;
    ndn3_11 <= n2560;
    ndn3_15 <= n2565;
    ndn3_21 <= n2570;
    n_n7584 <= n2575;
    n_n8354 <= n2580;
    n_n6952 <= n2585;
    n_n8864 <= n2590;
    n_n7930 <= n2595;
    n_n7962 <= n2600;
    n_n7929 <= n2605;
    n_n9316 <= n2610;
    n_n9102 <= n2615;
    n_n7308 <= n2620;
    n_n7657 <= n2625;
    n_n9264 <= n2630;
    n_n8760 <= n2635;
    n_n6912 <= n2640;
    n_n7887 <= n2645;
    n_n8911 <= n2650;
    n_n7952 <= n2655;
    n_n8704 <= n2660;
    n_n7876 <= n2665;
    n_n9596 <= n2670;
    n_n8430 <= n2675;
    n_n9019 <= n2680;
    n_n7699 <= n2685;
    n_n7375 <= n2690;
    n_n7936 <= n2695;
    n_n8340 <= n2700;
    n_n8809 <= n2705;
    n_n6961 <= n2710;
    n_n9429 <= n2715;
    n_n7743 <= n2720;
    n_n8980 <= n2725;
    n_n7582 <= n2730;
    n_n8968 <= n2735;
    n_n9371 <= n2740;
    n_n8741 <= n2745;
    n_n9502 <= n2750;
    n_n9373 <= n2755;
    n_n9248 <= n2760;
    n_n7822 <= n2765;
    n_n9054 <= n2770;
    n_n8273 <= n2775;
    n_n6937 <= n2780;
    n_n9342 <= n2785;
    n_n9325 <= n2790;
    n_n9609 <= n2795;
    n_n9623 <= n2800;
    n_n9470 <= n2805;
    n_n7570 <= n2810;
    n_n9310 <= n2815;
    n_n9366 <= n2820;
    n_n7181 <= n2825;
    n_n8739 <= n2830;
    n_n8939 <= n2835;
    n_n7256 <= n2840;
    n_n8983 <= n2845;
    n_n7487 <= n2850;
    n_n9268 <= n2855;
    n_n8906 <= n2860;
    n_n7988 <= n2865;
    n_n9181 <= n2870;
    n_n8725 <= n2875;
    n_n8626 <= n2880;
    ndn3_27 <= n2885;
    n_n8210 <= n2890;
    n_n7415 <= n2895;
    n_n8900 <= n2900;
    nen3_19 <= n2905;
    n_n8762 <= n2910;
    n_n8512 <= n2915;
    n_n8095 <= n2920;
    n_n8982 <= n2925;
    n_n7387 <= n2930;
    n_n9494 <= n2935;
    n_n7689 <= n2940;
    n_n7835 <= n2945;
    n_n9157 <= n2950;
    n_n8552 <= n2955;
    n_n7381 <= n2960;
    n_n9446 <= n2965;
    n_n8633 <= n2970;
    n_n7684 <= n2975;
    n_n7310 <= n2980;
    n_n8402 <= n2985;
    n_n9315 <= n2990;
    n_n7950 <= n2995;
    n_n8504 <= n3000;
    n_n8456 <= n3005;
    n_n7514 <= n3010;
    n_n7315 <= n3015;
    n_n9476 <= n3020;
    n_n8276 <= n3025;
    n_n8833 <= n3030;
    n_n7923 <= n3035;
    n_n9395 <= n3040;
    n_n9512 <= n3045;
    n_n9319 <= n3050;
    nsr3_35 <= n3055;
    n_n7154 <= n3060;
    n_n9495 <= n3065;
    n_n9137 <= n3070;
    n_n8854 <= n3075;
    n_n9183 <= n3080;
    n_n9323 <= n3085;
    n_n9349 <= n3090;
    n_n7896 <= n3095;
    n_n8073 <= n3100;
    n_n8970 <= n3105;
    n_n9314 <= n3110;
    n_n8486 <= n3115;
    n_n7246 <= n3120;
    n_n7866 <= n3125;
    n_n9599 <= n3130;
    n_n7635 <= n3135;
    n_n8984 <= n3140;
    n_n7360 <= n3145;
    n_n8794 <= n3150;
    n_n9108 <= n3155;
    n_n9286 <= n3160;
    ndn3_12 <= n3165;
    ndn3_16 <= n3170;
    n_n7708 <= n3175;
    n_n7807 <= n3180;
    n_n7650 <= n3185;
    n_n7947 <= n3190;
    n_n9500 <= n3195;
    n_n7734 <= n3200;
    n_n8464 <= n3205;
    n_n7659 <= n3210;
    n_n7630 <= n3215;
    n_n7756 <= n3220;
    n_n8691 <= n3225;
    n_n9176 <= n3230;
    n_n9327 <= n3235;
    n_n7995 <= n3240;
    n_n7395 <= n3245;
    n_n7878 <= n3250;
    n_n7507 <= n3255;
    n_n7959 <= n3260;
    n_n7825 <= n3265;
    n_n8009 <= n3270;
    n_n8281 <= n3275;
    n_n7685 <= n3280;
    n_n8106 <= n3285;
    n_n7687 <= n3290;
    n_n7766 <= n3295;
    n_n7880 <= n3300;
    n_n8961 <= n3305;
    n_n8014 <= n3310;
    n_n9278 <= n3315;
    n_n9087 <= n3320;
    n_n9182 <= n3325;
    n_n7852 <= n3330;
    n_n9324 <= n3335;
    nak3_13 <= n3340;
    n_n9416 <= n3345;
    nsr3_14 <= n3350;
    n_n8603 <= n3355;
    n_n7026 <= n3360;
    n_n8856 <= n3365;
    n_n8272 <= n3370;
    n_n9312 <= n3375;
    n_n7985 <= n3380;
    n_n8312 <= n3385;
    n_n7231 <= n3390;
    n_n9396 <= n3395;
    n_n8801 <= n3400;
    n_n8683 <= n3405;
    ndn3_39 <= n3410;
    n_n8245 <= n3415;
    n_n9458 <= n3420;
    n_n9302 <= n3425;
    n_n7392 <= n3430;
    n_n6963 <= n3435;
    n_n7808 <= n3440;
    n_n7225 <= n3445;
    n_n7817 <= n3450;
    n_n8201 <= n3455;
    n_n7793 <= n3460;
    n_n8177 <= n3465;
    n_n8389 <= n3470;
    n_n9440 <= n3475;
    n_n7683 <= n3480;
    n_n7761 <= n3485;
    n_n7667 <= n3490;
    n_n7980 <= n3495;
    n_n7509 <= n3500;
    n_n7813 <= n3505;
    n_n8396 <= n3510;
    n_n9535 <= n3515;
    n_n7209 <= n3520;
    n_n7003 <= n3525;
    n_n7695 <= n3530;
    n_n7624 <= n3535;
    n_n8791 <= n3540;
    n_n7374 <= n3545;
    n_n7429 <= n3550;
    n_n7944 <= n3555;
    n_n9266 <= n3560;
    n_n8100 <= n3565;
    n_n6988 <= n3570;
    n_n6986 <= n3575;
    n_n8933 <= n3580;
    n_n7117 <= n3585;
    n_n9043 <= n3590;
    n_n8241 <= n3595;
    n_n9219 <= n3600;
    n_n8198 <= n3605;
    n_n8081 <= n3610;
    n_n8575 <= n3615;
    n_n8710 <= n3620;
    n_n7622 <= n3625;
    n_n7966 <= n3630;
    n_n7885 <= n3635;
    n_n7033 <= n3640;
    ndn3_34 <= n3645;
    n_n9186 <= n3650;
    ndn3_50 <= n3655;
    n_n7879 <= n3660;
    n_n7019 <= n3665;
    n_n9171 <= n3670;
    n_n7261 <= n3675;
    n_n8223 <= n3680;
    n_n8989 <= n3685;
    n_n7993 <= n3690;
    n_n7845 <= n3695;
    n_n8253 <= n3700;
    n_n8889 <= n3705;
    n_n7809 <= n3710;
    n_n8918 <= n3715;
    n_n8515 <= n3720;
    n_n7933 <= n3725;
    n_n8075 <= n3730;
    n_n7338 <= n3735;
    n_n8104 <= n3740;
    n_n8171 <= n3745;
    n_n9059 <= n3750;
    n_n9023 <= n3755;
    n_n7692 <= n3760;
    n_n9441 <= n3765;
    n_n6920 <= n3770;
    n_n8831 <= n3775;
    n_n8441 <= n3780;
    n_n9576 <= n3785;
    n_n9252 <= n3790;
    n_n9363 <= n3795;
    ndn3_4 <= n3800;
    n_n9247 <= n3805;
    n_n7561 <= n3810;
    n_n8923 <= n3815;
    n_n7978 <= n3820;
    n_n8978 <= n3825;
    n_n9499 <= n3830;
    n_n8713 <= n3835;
    n_n8944 <= n3840;
    n_n8239 <= n3845;
    n_n7652 <= n3850;
    n_n9042 <= n3855;
    n_n8530 <= n3860;
    n_n9271 <= n3865;
    n_n9318 <= n3870;
    n_n7706 <= n3875;
    n_n7964 <= n3880;
    n_n8222 <= n3885;
    n_n8898 <= n3890;
    n_n7976 <= n3895;
    n_n7649 <= n3900;
    n_n7604 <= n3905;
    n_n7961 <= n3910;
    n_n7424 <= n3915;
    n_n7476 <= n3920;
    n_n9259 <= n3925;
    n_n9309 <= n3930;
    n_n9161 <= n3935;
    n_n8436 <= n3940;
    n_n9121 <= n3945;
    n_n8061 <= n3950;
    n_n8004 <= n3955;
    n_n9360 <= n3960;
    n_n9205 <= n3965;
    n_n8392 <= n3970;
    n_n9034 <= n3975;
    n_n8375 <= n3980;
    n_n8328 <= n3985;
    n_n9298 <= n3990;
    n_n7598 <= n3995;
    n_n8506 <= n4000;
    pdn <= n4005;
    n_n7737 <= n4009;
    n_n7420 <= n4014;
    n_n9291 <= n4019;
    n_n7946 <= n4024;
    n_n8584 <= n4029;
    n_n9308 <= n4034;
    n_n9403 <= n4039;
    n_n7284 <= n4044;
    n_n9270 <= n4049;
    n_n7390 <= n4054;
    n_n9351 <= n4059;
    n_n6968 <= n4064;
    n_n8668 <= n4069;
    n_n9605 <= n4074;
    n_n7013 <= n4079;
    n_n9626 <= n4084;
    n_n8200 <= n4089;
    n_n9028 <= n4094;
    n_n8803 <= n4099;
    n_n9570 <= n4104;
    n_n8366 <= n4109;
    n_n9050 <= n4114;
    n_n8650 <= n4119;
    n_n8574 <= n4124;
    n_n7276 <= n4129;
    n_n9212 <= n4134;
    n_n8384 <= n4139;
    ndn3_35 <= n4144;
    n_n8449 <= n4149;
    ndn3_46 <= n4154;
    n_n7554 <= n4159;
    n_n8743 <= n4164;
    n_n8277 <= n4169;
    n_n9359 <= n4174;
    n_n8425 <= n4179;
    n_n9104 <= n4184;
    n_n9221 <= n4189;
    n_n9448 <= n4194;
    n_n9537 <= n4199;
    n_n8003 <= n4204;
    n_n7467 <= n4209;
    n_n8233 <= n4214;
    n_n7932 <= n4219;
    n_n8064 <= n4224;
    n_n9162 <= n4229;
    n_n7971 <= n4234;
    n_n8055 <= n4239;
    n_n7711 <= n4244;
    n_n8256 <= n4249;
    n_n7925 <= n4254;
    n_n7762 <= n4259;
    n_n7668 <= n4264;
    n_n7914 <= n4269;
    n_n7873 <= n4274;
    n_n7849 <= n4279;
    n_n9421 <= n4284;
    n_n7626 <= n4289;
    n_n7848 <= n4294;
    n_n8263 <= n4299;
    n_n9100 <= n4304;
    n_n9393 <= n4309;
    n_n9591 <= n4314;
    n_n7588 <= n4319;
    n_n9123 <= n4324;
    n_n9159 <= n4329;
    n_n9128 <= n4334;
    n_n8045 <= n4339;
    n_n7728 <= n4344;
    n_n8929 <= n4349;
    n_n7739 <= n4354;
    n_n9355 <= n4359;
    n_n9394 <= n4364;
    n_n8470 <= n4369;
    n_n8571 <= n4374;
    n_n8796 <= n4379;
    ndn3_36 <= n4384;
    n_n7990 <= n4389;
    n_n8781 <= n4394;
    n_n8817 <= n4399;
    n_n9160 <= n4404;
    n_n9092 <= n4409;
    n_n8513 <= n4414;
    n_n8213 <= n4419;
    n_n8581 <= n4424;
    n_n9284 <= n4429;
    n_n7837 <= n4434;
    n_n8224 <= n4439;
    n_n9203 <= n4444;
    n_n7655 <= n4449;
    n_n8946 <= n4454;
    n_n7052 <= n4459;
    n_n9615 <= n4464;
    n_n8473 <= n4469;
    n_n7741 <= n4474;
    n_n9460 <= n4479;
    n_n7912 <= n4484;
    n_n7606 <= n4489;
    n_n9021 <= n4494;
    n_n7781 <= n4499;
    n_n7810 <= n4504;
    n_n7108 <= n4509;
    n_n7697 <= n4514;
    n_n7642 <= n4519;
    n_n9595 <= n4524;
    n_n7694 <= n4529;
    n_n8221 <= n4534;
    n_n7600 <= n4539;
    n_n7935 <= n4544;
    n_n9230 <= n4549;
    n_n7701 <= n4554;
    n_n7510 <= n4559;
    n_n7627 <= n4564;
    n_n8502 <= n4569;
    n_n8516 <= n4574;
    n_n7913 <= n4579;
    n_n9320 <= n4584;
    n_n7411 <= n4589;
    n_n9129 <= n4594;
    n_n9053 <= n4599;
    n_n7069 <= n4604;
    n_n8617 <= n4609;
    n_n7242 <= n4614;
    n_n8230 <= n4619;
    n_n9294 <= n4624;
    n_n8249 <= n4629;
    n_n8972 <= n4634;
    n_n7074 <= n4639;
    n_n7493 <= n4644;
    n_n8290 <= n4649;
    n_n8821 <= n4654;
    n_n7769 <= n4659;
    n_n7491 <= n4664;
    n_n9600 <= n4669;
    n_n9317 <= n4674;
    n_n8047 <= n4679;
    n_n9629 <= n4684;
    n_n9126 <= n4689;
    n_n9508 <= n4694;
    n_n9155 <= n4699;
    n_n8528 <= n4704;
    ndn3_37 <= n4709;
    ndn3_42 <= n4714;
    n_n9358 <= n4719;
    n_n8185 <= n4724;
    nen3_28 <= n4729;
    n_n8839 <= n4734;
    n_n7903 <= n4739;
    n_n9139 <= n4744;
    n_n9075 <= n4749;
    n_n9439 <= n4754;
    n_n9353 <= n4759;
    n_n7665 <= n4764;
    n_n8798 <= n4769;
    n_n7146 <= n4774;
    n_n7890 <= n4779;
    n_n7176 <= n4784;
    n_n8477 <= n4789;
    n_n8514 <= n4794;
    n_n8636 <= n4799;
    n_n7183 <= n4804;
    n_n8657 <= n4809;
    n_n9493 <= n4814;
    n_n7969 <= n4819;
    n_n9255 <= n4824;
    n_n8535 <= n4829;
    n_n8619 <= n4834;
    n_n8909 <= n4839;
    n_n7744 <= n4844;
    n_n9119 <= n4849;
    n_n7827 <= n4854;
    n_n8916 <= n4859;
    n_n8729 <= n4864;
    n_n9011 <= n4869;
    n_n8779 <= n4874;
    n_n6980 <= n4879;
    n_n7715 <= n4884;
    n_n9067 <= n4889;
    n_n9164 <= n4894;
    n_n7402 <= n4899;
    n_n8938 <= n4904;
    n_n9046 <= n4909;
    n_n8789 <= n4914;
    n_n9390 <= n4919;
    n_n7768 <= n4924;
    n_n9136 <= n4929;
    n_n8670 <= n4934;
    n_n8644 <= n4939;
    n_n9178 <= n4944;
    n_n8188 <= n4949;
    n_n7083 <= n4954;
    n_n9344 <= n4959;
    n_n7366 <= n4964;
    n_n8361 <= n4969;
    n_n9228 <= n4974;
    n_n9402 <= n4979;
    n_n8510 <= n4984;
    n_n8881 <= n4989;
    n_n9404 <= n4994;
    n_n9424 <= n4999;
    n_n9031 <= n5004;
    nsr3_37 <= n5009;
    n_n8197 <= n5014;
    n_n8468 <= n5019;
    n_n7121 <= n5024;
    n_n7511 <= n5029;
    ndn3_44 <= n5034;
    n_n9322 <= n5039;
    n_n7682 <= n5044;
    n_n9603 <= n5049;
    nlc1_2 <= n5054;
    n_n8408 <= n5059;
    n_n8577 <= n5064;
    n_n7079 <= n5069;
    n_n8828 <= n5074;
    n_n9340 <= n5079;
    n_n8586 <= n5084;
    n_n7901 <= n5089;
    n_n8628 <= n5094;
    n_n8869 <= n5099;
    n_n7710 <= n5104;
    n_n8993 <= n5109;
    n_n9586 <= n5114;
    n_n8852 <= n5119;
    n_n8583 <= n5124;
    n_n8011 <= n5129;
    n_n7717 <= n5134;
    n_n8326 <= n5139;
    n_n9163 <= n5144;
    n_n8344 <= n5149;
    n_n8296 <= n5154;
    n_n8116 <= n5159;
    n_n8267 <= n5164;
    n_n7686 <= n5169;
    n_n9061 <= n5174;
    n_n9338 <= n5179;
    n_n7688 <= n5184;
    n_n9081 <= n5189;
    n_n6910 <= n5194;
    n_n8727 <= n5199;
    n_n7674 <= n5204;
    n_n7330 <= n5209;
    n_n8966 <= n5214;
    n_n7843 <= n5219;
    n_n8847 <= n5224;
    n_n9376 <= n5229;
    n_n7553 <= n5234;
    n_n9292 <= n5239;
    n_n7464 <= n5244;
    n_n8146 <= n5249;
    n_n8439 <= n5254;
    n_n9498 <= n5259;
    n_n8118 <= n5264;
    n_n9452 <= n5269;
    n_n9239 <= n5274;
    n_n9237 <= n5279;
    n_n9488 <= n5284;
    ndn3_2 <= n5289;
    n_n9522 <= n5294;
    n_n9313 <= n5299;
    n_n7435 <= n5304;
    n_n8665 <= n5309;
    n_n9593 <= n5314;
    n_n8303 <= n5319;
    n_n7022 <= n5324;
    n_n9173 <= n5329;
    n_n9261 <= n5334;
    n_n7150 <= n5339;
    n_n9455 <= n5344;
    n_n8371 <= n5349;
    nsr3_20 <= n5354;
    n_n8271 <= n5359;
    n_n9542 <= n5364;
    n_n7444 <= n5369;
    ndn3_40 <= n5374;
    n_n7130 <= n5379;
    n_n9347 <= n5384;
    n_n8102 <= n5389;
    n_n9225 <= n5394;
    n_n8462 <= n5399;
    n_n8088 <= n5404;
    n_n9026 <= n5409;
    n_n9289 <= n5414;
    n_n7661 <= n5419;
    n_n8108 <= n5424;
    n_n8921 <= n5429;
    n_n7859 <= n5434;
    n_n7732 <= n5439;
    n_n7956 <= n5444;
    n_n9520 <= n5449;
    n_n7666 <= n5454;
    n_n7678 <= n5459;
    n_n7846 <= n5464;
    n_n8280 <= n5469;
    n_n8841 <= n5474;
    n_n7336 <= n5479;
    n_n8226 <= n5484;
    n_n8151 <= n5489;
    n_n7644 <= n5494;
    n_n8770 <= n5499;
    n_n8423 <= n5504;
    n_n7763 <= n5509;
    n_n9525 <= n5514;
    n_n8033 <= n5519;
    n_n7881 <= n5524;
    n_n7815 <= n5529;
    n_n9232 <= n5534;
    n_n7792 <= n5539;
    n_n9563 <= n5544;
    n_n8672 <= n5549;
    n_n7346 <= n5554;
    n_n7949 <= n5559;
    n_n8756 <= n5564;
    n_n8641 <= n5569;
    n_n8192 <= n5574;
    n_n8058 <= n5579;
    n_n8561 <= n5584;
    n_n9306 <= n5589;
    n_n9165 <= n5594;
    n_n8850 <= n5599;
    n_n9210 <= n5604;
    ndn2_2 <= n5609;
    n_n7342 <= n5614;
    n_n8051 <= n5619;
    n_n7136 <= n5624;
    n_n9348 <= n5629;
    n_n9006 <= n5634;
    n_n7653 <= n5639;
    n_n7905 <= n5644;
    n_n9166 <= n5649;
    n_n7065 <= n5654;
    n_n9490 <= n5659;
    n_n7024 <= n5664;
    n_n7586 <= n5669;
    n_n8416 <= n5674;
    n_n8937 <= n5679;
    n_n8141 <= n5684;
    n_n7853 <= n5689;
    n_n8121 <= n5694;
    n_n9604 <= n5699;
    n_n9496 <= n5704;
    n_n8195 <= n5709;
    n_n9516 <= n5714;
    n_n9077 <= n5719;
    n_n9436 <= n5724;
    n_n9051 <= n5729;
    n_n7664 <= n5734;
    n_n8419 <= n5739;
    n_n7874 <= n5744;
    n_n9133 <= n5749;
    n_n9392 <= n5754;
    n_n7770 <= n5759;
    ndn3_32 <= n5764;
    n_n7601 <= n5769;
    n_n8206 <= n5774;
    n_n7927 <= n5779;
    n_n9606 <= n5784;
    n_n7111 <= n5789;
    n_n9269 <= n5794;
    ndn3_38 <= n5799;
    n_n7886 <= n5804;
    n_n9179 <= n5809;
    n_n9357 <= n5814;
    n_n9594 <= n5819;
    n_n7628 <= n5824;
    n_n8454 <= n5829;
    ndn3_20 <= n5834;
    n_n9505 <= n5839;
    nen3_34 <= n5844;
    n_n9632 <= n5849;
    n_n7076 <= n5854;
    n_n9262 <= n5859;
    n_n9048 <= n5864;
    n_n9578 <= n5869;
    n_n8135 <= n5874;
    ndn3_26 <= n5879;
    n_n7500 <= n5884;
    n_n6974 <= n5889;
    n_n8605 <= n5894;
    n_n9296 <= n5899;
    n_n7156 <= n5904;
    n_n7920 <= n5909;
    n_n8895 <= n5914;
    n_n8991 <= n5919;
    n_n8139 <= n5924;
    n_n9275 <= n5929;
    n_n7203 <= n5934;
    n_n9590 <= n5939;
    n_n7344 <= n5944;
    n_n6976 <= n5949;
    n_n7629 <= n5954;
    ndn3_14 <= n5959;
    n_n7862 <= n5964;
    n_n9013 <= n5969;
    n_n7288 <= n5974;
    n_n8078 <= n5979;
    n_n7334 <= n5984;
    n_n7704 <= n5989;
    n_n7788 <= n5994;
    n_n8526 <= n5999;
    n_n9556 <= n6004;
    n_n9345 <= n6009;
    n_n8447 <= n6014;
    n_n7485 <= n6019;
    n_n8570 <= n6024;
    n_n7453 <= n6029;
    n_n7928 <= n6034;
    n_n8646 <= n6039;
    n_n9405 <= n6044;
    n_n8948 <= n6049;
    n_n9131 <= n6054;
    n_n8216 <= n6059;
    n_n9177 <= n6064;
    n_n7844 <= n6069;
    n_n8811 <= n6074;
    n_n9145 <= n6079;
    n_n8428 <= n6084;
    n_n8858 <= n6089;
    n_n8580 <= n6094;
  end
endmodule


