*****************************
*     FPGA SPICE Netlist    *
* Description: Connection Block X-channel  [1][0] in FPGA *
*    Author: Xifan TANG     *
* Organization: EPFL/IC/LSI *
* Date: Thu Nov 15 14:26:08 2018
 *
*****************************
.subckt cbx[1][0] 
+ chanx[1][0]_midout[0] 
+ chanx[1][0]_midout[1] 
+ chanx[1][0]_midout[2] 
+ chanx[1][0]_midout[3] 
+ chanx[1][0]_midout[4] 
+ chanx[1][0]_midout[5] 
+ chanx[1][0]_midout[6] 
+ chanx[1][0]_midout[7] 
+ chanx[1][0]_midout[8] 
+ chanx[1][0]_midout[9] 
+ chanx[1][0]_midout[10] 
+ chanx[1][0]_midout[11] 
+ chanx[1][0]_midout[12] 
+ chanx[1][0]_midout[13] 
+ chanx[1][0]_midout[14] 
+ chanx[1][0]_midout[15] 
+ chanx[1][0]_midout[16] 
+ chanx[1][0]_midout[17] 
+ chanx[1][0]_midout[18] 
+ chanx[1][0]_midout[19] 
+ chanx[1][0]_midout[20] 
+ chanx[1][0]_midout[21] 
+ chanx[1][0]_midout[22] 
+ chanx[1][0]_midout[23] 
+ chanx[1][0]_midout[24] 
+ chanx[1][0]_midout[25] 
+ chanx[1][0]_midout[26] 
+ chanx[1][0]_midout[27] 
+ chanx[1][0]_midout[28] 
+ chanx[1][0]_midout[29] 
+ chanx[1][0]_midout[30] 
+ chanx[1][0]_midout[31] 
+ chanx[1][0]_midout[32] 
+ chanx[1][0]_midout[33] 
+ chanx[1][0]_midout[34] 
+ chanx[1][0]_midout[35] 
+ chanx[1][0]_midout[36] 
+ chanx[1][0]_midout[37] 
+ chanx[1][0]_midout[38] 
+ chanx[1][0]_midout[39] 
+ chanx[1][0]_midout[40] 
+ chanx[1][0]_midout[41] 
+ chanx[1][0]_midout[42] 
+ chanx[1][0]_midout[43] 
+ chanx[1][0]_midout[44] 
+ chanx[1][0]_midout[45] 
+ chanx[1][0]_midout[46] 
+ chanx[1][0]_midout[47] 
+ chanx[1][0]_midout[48] 
+ chanx[1][0]_midout[49] 
+ chanx[1][0]_midout[50] 
+ chanx[1][0]_midout[51] 
+ chanx[1][0]_midout[52] 
+ chanx[1][0]_midout[53] 
+ chanx[1][0]_midout[54] 
+ chanx[1][0]_midout[55] 
+ chanx[1][0]_midout[56] 
+ chanx[1][0]_midout[57] 
+ chanx[1][0]_midout[58] 
+ chanx[1][0]_midout[59] 
+ chanx[1][0]_midout[60] 
+ chanx[1][0]_midout[61] 
+ chanx[1][0]_midout[62] 
+ chanx[1][0]_midout[63] 
+ chanx[1][0]_midout[64] 
+ chanx[1][0]_midout[65] 
+ chanx[1][0]_midout[66] 
+ chanx[1][0]_midout[67] 
+ chanx[1][0]_midout[68] 
+ chanx[1][0]_midout[69] 
+ chanx[1][0]_midout[70] 
+ chanx[1][0]_midout[71] 
+ chanx[1][0]_midout[72] 
+ chanx[1][0]_midout[73] 
+ chanx[1][0]_midout[74] 
+ chanx[1][0]_midout[75] 
+ chanx[1][0]_midout[76] 
+ chanx[1][0]_midout[77] 
+ chanx[1][0]_midout[78] 
+ chanx[1][0]_midout[79] 
+ chanx[1][0]_midout[80] 
+ chanx[1][0]_midout[81] 
+ chanx[1][0]_midout[82] 
+ chanx[1][0]_midout[83] 
+ chanx[1][0]_midout[84] 
+ chanx[1][0]_midout[85] 
+ chanx[1][0]_midout[86] 
+ chanx[1][0]_midout[87] 
+ chanx[1][0]_midout[88] 
+ chanx[1][0]_midout[89] 
+ chanx[1][0]_midout[90] 
+ chanx[1][0]_midout[91] 
+ chanx[1][0]_midout[92] 
+ chanx[1][0]_midout[93] 
+ chanx[1][0]_midout[94] 
+ chanx[1][0]_midout[95] 
+ chanx[1][0]_midout[96] 
+ chanx[1][0]_midout[97] 
+ chanx[1][0]_midout[98] 
+ chanx[1][0]_midout[99] 
+ grid[1][1]_pin[0][2][2] 
+ grid[1][1]_pin[0][2][6] 
+ grid[1][1]_pin[0][2][10] 
+ grid[1][1]_pin[0][2][14] 
+ grid[1][1]_pin[0][2][18] 
+ grid[1][1]_pin[0][2][22] 
+ grid[1][1]_pin[0][2][26] 
+ grid[1][1]_pin[0][2][30] 
+ grid[1][1]_pin[0][2][34] 
+ grid[1][1]_pin[0][2][38] 
+ grid[1][1]_pin[0][2][50] 
+ grid[1][0]_pin[0][0][0] 
+ grid[1][0]_pin[0][0][2] 
+ grid[1][0]_pin[0][0][4] 
+ grid[1][0]_pin[0][0][6] 
+ grid[1][0]_pin[0][0][8] 
+ grid[1][0]_pin[0][0][10] 
+ grid[1][0]_pin[0][0][12] 
+ grid[1][0]_pin[0][0][14] 
+ svdd sgnd
Xmux_2level_tapbuf_size16[0] chanx[1][0]_midout[0] chanx[1][0]_midout[1] chanx[1][0]_midout[12] chanx[1][0]_midout[13] chanx[1][0]_midout[24] chanx[1][0]_midout[25] chanx[1][0]_midout[38] chanx[1][0]_midout[39] chanx[1][0]_midout[50] chanx[1][0]_midout[51] chanx[1][0]_midout[62] chanx[1][0]_midout[63] chanx[1][0]_midout[74] chanx[1][0]_midout[75] chanx[1][0]_midout[88] chanx[1][0]_midout[89] grid[1][1]_pin[0][2][2] sram[2082]->outb sram[2082]->out sram[2083]->out sram[2083]->outb sram[2084]->out sram[2084]->outb sram[2085]->out sram[2085]->outb sram[2086]->outb sram[2086]->out sram[2087]->out sram[2087]->outb sram[2088]->out sram[2088]->outb sram[2089]->out sram[2089]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[0], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2082] sram->in sram[2082]->out sram[2082]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2082]->out) 0
.nodeset V(sram[2082]->outb) vsp
Xsram[2083] sram->in sram[2083]->out sram[2083]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2083]->out) 0
.nodeset V(sram[2083]->outb) vsp
Xsram[2084] sram->in sram[2084]->out sram[2084]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2084]->out) 0
.nodeset V(sram[2084]->outb) vsp
Xsram[2085] sram->in sram[2085]->out sram[2085]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2085]->out) 0
.nodeset V(sram[2085]->outb) vsp
Xsram[2086] sram->in sram[2086]->out sram[2086]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2086]->out) 0
.nodeset V(sram[2086]->outb) vsp
Xsram[2087] sram->in sram[2087]->out sram[2087]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2087]->out) 0
.nodeset V(sram[2087]->outb) vsp
Xsram[2088] sram->in sram[2088]->out sram[2088]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2088]->out) 0
.nodeset V(sram[2088]->outb) vsp
Xsram[2089] sram->in sram[2089]->out sram[2089]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2089]->out) 0
.nodeset V(sram[2089]->outb) vsp
Xmux_2level_tapbuf_size16[1] chanx[1][0]_midout[0] chanx[1][0]_midout[1] chanx[1][0]_midout[14] chanx[1][0]_midout[15] chanx[1][0]_midout[26] chanx[1][0]_midout[27] chanx[1][0]_midout[38] chanx[1][0]_midout[39] chanx[1][0]_midout[50] chanx[1][0]_midout[51] chanx[1][0]_midout[64] chanx[1][0]_midout[65] chanx[1][0]_midout[76] chanx[1][0]_midout[77] chanx[1][0]_midout[88] chanx[1][0]_midout[89] grid[1][1]_pin[0][2][6] sram[2090]->outb sram[2090]->out sram[2091]->out sram[2091]->outb sram[2092]->out sram[2092]->outb sram[2093]->out sram[2093]->outb sram[2094]->outb sram[2094]->out sram[2095]->out sram[2095]->outb sram[2096]->out sram[2096]->outb sram[2097]->out sram[2097]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[1], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2090] sram->in sram[2090]->out sram[2090]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2090]->out) 0
.nodeset V(sram[2090]->outb) vsp
Xsram[2091] sram->in sram[2091]->out sram[2091]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2091]->out) 0
.nodeset V(sram[2091]->outb) vsp
Xsram[2092] sram->in sram[2092]->out sram[2092]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2092]->out) 0
.nodeset V(sram[2092]->outb) vsp
Xsram[2093] sram->in sram[2093]->out sram[2093]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2093]->out) 0
.nodeset V(sram[2093]->outb) vsp
Xsram[2094] sram->in sram[2094]->out sram[2094]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2094]->out) 0
.nodeset V(sram[2094]->outb) vsp
Xsram[2095] sram->in sram[2095]->out sram[2095]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2095]->out) 0
.nodeset V(sram[2095]->outb) vsp
Xsram[2096] sram->in sram[2096]->out sram[2096]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2096]->out) 0
.nodeset V(sram[2096]->outb) vsp
Xsram[2097] sram->in sram[2097]->out sram[2097]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2097]->out) 0
.nodeset V(sram[2097]->outb) vsp
Xmux_2level_tapbuf_size16[2] chanx[1][0]_midout[2] chanx[1][0]_midout[3] chanx[1][0]_midout[14] chanx[1][0]_midout[15] chanx[1][0]_midout[28] chanx[1][0]_midout[29] chanx[1][0]_midout[40] chanx[1][0]_midout[41] chanx[1][0]_midout[52] chanx[1][0]_midout[53] chanx[1][0]_midout[64] chanx[1][0]_midout[65] chanx[1][0]_midout[78] chanx[1][0]_midout[79] chanx[1][0]_midout[90] chanx[1][0]_midout[91] grid[1][1]_pin[0][2][10] sram[2098]->outb sram[2098]->out sram[2099]->out sram[2099]->outb sram[2100]->out sram[2100]->outb sram[2101]->out sram[2101]->outb sram[2102]->outb sram[2102]->out sram[2103]->out sram[2103]->outb sram[2104]->out sram[2104]->outb sram[2105]->out sram[2105]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[2], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2098] sram->in sram[2098]->out sram[2098]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2098]->out) 0
.nodeset V(sram[2098]->outb) vsp
Xsram[2099] sram->in sram[2099]->out sram[2099]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2099]->out) 0
.nodeset V(sram[2099]->outb) vsp
Xsram[2100] sram->in sram[2100]->out sram[2100]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2100]->out) 0
.nodeset V(sram[2100]->outb) vsp
Xsram[2101] sram->in sram[2101]->out sram[2101]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2101]->out) 0
.nodeset V(sram[2101]->outb) vsp
Xsram[2102] sram->in sram[2102]->out sram[2102]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2102]->out) 0
.nodeset V(sram[2102]->outb) vsp
Xsram[2103] sram->in sram[2103]->out sram[2103]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2103]->out) 0
.nodeset V(sram[2103]->outb) vsp
Xsram[2104] sram->in sram[2104]->out sram[2104]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2104]->out) 0
.nodeset V(sram[2104]->outb) vsp
Xsram[2105] sram->in sram[2105]->out sram[2105]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2105]->out) 0
.nodeset V(sram[2105]->outb) vsp
Xmux_2level_tapbuf_size16[3] chanx[1][0]_midout[4] chanx[1][0]_midout[5] chanx[1][0]_midout[16] chanx[1][0]_midout[17] chanx[1][0]_midout[28] chanx[1][0]_midout[29] chanx[1][0]_midout[40] chanx[1][0]_midout[41] chanx[1][0]_midout[54] chanx[1][0]_midout[55] chanx[1][0]_midout[66] chanx[1][0]_midout[67] chanx[1][0]_midout[78] chanx[1][0]_midout[79] chanx[1][0]_midout[90] chanx[1][0]_midout[91] grid[1][1]_pin[0][2][14] sram[2106]->outb sram[2106]->out sram[2107]->out sram[2107]->outb sram[2108]->out sram[2108]->outb sram[2109]->out sram[2109]->outb sram[2110]->outb sram[2110]->out sram[2111]->out sram[2111]->outb sram[2112]->out sram[2112]->outb sram[2113]->out sram[2113]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[3], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2106] sram->in sram[2106]->out sram[2106]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2106]->out) 0
.nodeset V(sram[2106]->outb) vsp
Xsram[2107] sram->in sram[2107]->out sram[2107]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2107]->out) 0
.nodeset V(sram[2107]->outb) vsp
Xsram[2108] sram->in sram[2108]->out sram[2108]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2108]->out) 0
.nodeset V(sram[2108]->outb) vsp
Xsram[2109] sram->in sram[2109]->out sram[2109]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2109]->out) 0
.nodeset V(sram[2109]->outb) vsp
Xsram[2110] sram->in sram[2110]->out sram[2110]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2110]->out) 0
.nodeset V(sram[2110]->outb) vsp
Xsram[2111] sram->in sram[2111]->out sram[2111]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2111]->out) 0
.nodeset V(sram[2111]->outb) vsp
Xsram[2112] sram->in sram[2112]->out sram[2112]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2112]->out) 0
.nodeset V(sram[2112]->outb) vsp
Xsram[2113] sram->in sram[2113]->out sram[2113]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2113]->out) 0
.nodeset V(sram[2113]->outb) vsp
Xmux_2level_tapbuf_size16[4] chanx[1][0]_midout[4] chanx[1][0]_midout[5] chanx[1][0]_midout[18] chanx[1][0]_midout[19] chanx[1][0]_midout[30] chanx[1][0]_midout[31] chanx[1][0]_midout[42] chanx[1][0]_midout[43] chanx[1][0]_midout[54] chanx[1][0]_midout[55] chanx[1][0]_midout[68] chanx[1][0]_midout[69] chanx[1][0]_midout[80] chanx[1][0]_midout[81] chanx[1][0]_midout[92] chanx[1][0]_midout[93] grid[1][1]_pin[0][2][18] sram[2114]->outb sram[2114]->out sram[2115]->out sram[2115]->outb sram[2116]->out sram[2116]->outb sram[2117]->out sram[2117]->outb sram[2118]->outb sram[2118]->out sram[2119]->out sram[2119]->outb sram[2120]->out sram[2120]->outb sram[2121]->out sram[2121]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[4], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2114] sram->in sram[2114]->out sram[2114]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2114]->out) 0
.nodeset V(sram[2114]->outb) vsp
Xsram[2115] sram->in sram[2115]->out sram[2115]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2115]->out) 0
.nodeset V(sram[2115]->outb) vsp
Xsram[2116] sram->in sram[2116]->out sram[2116]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2116]->out) 0
.nodeset V(sram[2116]->outb) vsp
Xsram[2117] sram->in sram[2117]->out sram[2117]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2117]->out) 0
.nodeset V(sram[2117]->outb) vsp
Xsram[2118] sram->in sram[2118]->out sram[2118]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2118]->out) 0
.nodeset V(sram[2118]->outb) vsp
Xsram[2119] sram->in sram[2119]->out sram[2119]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2119]->out) 0
.nodeset V(sram[2119]->outb) vsp
Xsram[2120] sram->in sram[2120]->out sram[2120]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2120]->out) 0
.nodeset V(sram[2120]->outb) vsp
Xsram[2121] sram->in sram[2121]->out sram[2121]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2121]->out) 0
.nodeset V(sram[2121]->outb) vsp
Xmux_2level_tapbuf_size16[5] chanx[1][0]_midout[6] chanx[1][0]_midout[7] chanx[1][0]_midout[18] chanx[1][0]_midout[19] chanx[1][0]_midout[30] chanx[1][0]_midout[31] chanx[1][0]_midout[44] chanx[1][0]_midout[45] chanx[1][0]_midout[56] chanx[1][0]_midout[57] chanx[1][0]_midout[68] chanx[1][0]_midout[69] chanx[1][0]_midout[80] chanx[1][0]_midout[81] chanx[1][0]_midout[94] chanx[1][0]_midout[95] grid[1][1]_pin[0][2][22] sram[2122]->outb sram[2122]->out sram[2123]->out sram[2123]->outb sram[2124]->out sram[2124]->outb sram[2125]->out sram[2125]->outb sram[2126]->out sram[2126]->outb sram[2127]->out sram[2127]->outb sram[2128]->out sram[2128]->outb sram[2129]->outb sram[2129]->out svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[5], level=2, select_path_id=3. *****
*****10000001*****
Xsram[2122] sram->in sram[2122]->out sram[2122]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2122]->out) 0
.nodeset V(sram[2122]->outb) vsp
Xsram[2123] sram->in sram[2123]->out sram[2123]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2123]->out) 0
.nodeset V(sram[2123]->outb) vsp
Xsram[2124] sram->in sram[2124]->out sram[2124]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2124]->out) 0
.nodeset V(sram[2124]->outb) vsp
Xsram[2125] sram->in sram[2125]->out sram[2125]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2125]->out) 0
.nodeset V(sram[2125]->outb) vsp
Xsram[2126] sram->in sram[2126]->out sram[2126]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2126]->out) 0
.nodeset V(sram[2126]->outb) vsp
Xsram[2127] sram->in sram[2127]->out sram[2127]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2127]->out) 0
.nodeset V(sram[2127]->outb) vsp
Xsram[2128] sram->in sram[2128]->out sram[2128]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2128]->out) 0
.nodeset V(sram[2128]->outb) vsp
Xsram[2129] sram->in sram[2129]->out sram[2129]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2129]->out) 0
.nodeset V(sram[2129]->outb) vsp
Xmux_2level_tapbuf_size16[6] chanx[1][0]_midout[8] chanx[1][0]_midout[9] chanx[1][0]_midout[20] chanx[1][0]_midout[21] chanx[1][0]_midout[32] chanx[1][0]_midout[33] chanx[1][0]_midout[44] chanx[1][0]_midout[45] chanx[1][0]_midout[58] chanx[1][0]_midout[59] chanx[1][0]_midout[70] chanx[1][0]_midout[71] chanx[1][0]_midout[82] chanx[1][0]_midout[83] chanx[1][0]_midout[94] chanx[1][0]_midout[95] grid[1][1]_pin[0][2][26] sram[2130]->outb sram[2130]->out sram[2131]->out sram[2131]->outb sram[2132]->out sram[2132]->outb sram[2133]->out sram[2133]->outb sram[2134]->outb sram[2134]->out sram[2135]->out sram[2135]->outb sram[2136]->out sram[2136]->outb sram[2137]->out sram[2137]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[6], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2130] sram->in sram[2130]->out sram[2130]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2130]->out) 0
.nodeset V(sram[2130]->outb) vsp
Xsram[2131] sram->in sram[2131]->out sram[2131]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2131]->out) 0
.nodeset V(sram[2131]->outb) vsp
Xsram[2132] sram->in sram[2132]->out sram[2132]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2132]->out) 0
.nodeset V(sram[2132]->outb) vsp
Xsram[2133] sram->in sram[2133]->out sram[2133]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2133]->out) 0
.nodeset V(sram[2133]->outb) vsp
Xsram[2134] sram->in sram[2134]->out sram[2134]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2134]->out) 0
.nodeset V(sram[2134]->outb) vsp
Xsram[2135] sram->in sram[2135]->out sram[2135]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2135]->out) 0
.nodeset V(sram[2135]->outb) vsp
Xsram[2136] sram->in sram[2136]->out sram[2136]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2136]->out) 0
.nodeset V(sram[2136]->outb) vsp
Xsram[2137] sram->in sram[2137]->out sram[2137]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2137]->out) 0
.nodeset V(sram[2137]->outb) vsp
Xmux_2level_tapbuf_size16[7] chanx[1][0]_midout[8] chanx[1][0]_midout[9] chanx[1][0]_midout[20] chanx[1][0]_midout[21] chanx[1][0]_midout[34] chanx[1][0]_midout[35] chanx[1][0]_midout[46] chanx[1][0]_midout[47] chanx[1][0]_midout[58] chanx[1][0]_midout[59] chanx[1][0]_midout[70] chanx[1][0]_midout[71] chanx[1][0]_midout[84] chanx[1][0]_midout[85] chanx[1][0]_midout[96] chanx[1][0]_midout[97] grid[1][1]_pin[0][2][30] sram[2138]->outb sram[2138]->out sram[2139]->out sram[2139]->outb sram[2140]->out sram[2140]->outb sram[2141]->out sram[2141]->outb sram[2142]->outb sram[2142]->out sram[2143]->out sram[2143]->outb sram[2144]->out sram[2144]->outb sram[2145]->out sram[2145]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[7], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2138] sram->in sram[2138]->out sram[2138]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2138]->out) 0
.nodeset V(sram[2138]->outb) vsp
Xsram[2139] sram->in sram[2139]->out sram[2139]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2139]->out) 0
.nodeset V(sram[2139]->outb) vsp
Xsram[2140] sram->in sram[2140]->out sram[2140]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2140]->out) 0
.nodeset V(sram[2140]->outb) vsp
Xsram[2141] sram->in sram[2141]->out sram[2141]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2141]->out) 0
.nodeset V(sram[2141]->outb) vsp
Xsram[2142] sram->in sram[2142]->out sram[2142]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2142]->out) 0
.nodeset V(sram[2142]->outb) vsp
Xsram[2143] sram->in sram[2143]->out sram[2143]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2143]->out) 0
.nodeset V(sram[2143]->outb) vsp
Xsram[2144] sram->in sram[2144]->out sram[2144]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2144]->out) 0
.nodeset V(sram[2144]->outb) vsp
Xsram[2145] sram->in sram[2145]->out sram[2145]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2145]->out) 0
.nodeset V(sram[2145]->outb) vsp
Xmux_2level_tapbuf_size16[8] chanx[1][0]_midout[10] chanx[1][0]_midout[11] chanx[1][0]_midout[22] chanx[1][0]_midout[23] chanx[1][0]_midout[34] chanx[1][0]_midout[35] chanx[1][0]_midout[48] chanx[1][0]_midout[49] chanx[1][0]_midout[60] chanx[1][0]_midout[61] chanx[1][0]_midout[72] chanx[1][0]_midout[73] chanx[1][0]_midout[84] chanx[1][0]_midout[85] chanx[1][0]_midout[98] chanx[1][0]_midout[99] grid[1][1]_pin[0][2][34] sram[2146]->outb sram[2146]->out sram[2147]->out sram[2147]->outb sram[2148]->out sram[2148]->outb sram[2149]->out sram[2149]->outb sram[2150]->outb sram[2150]->out sram[2151]->out sram[2151]->outb sram[2152]->out sram[2152]->outb sram[2153]->out sram[2153]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[8], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2146] sram->in sram[2146]->out sram[2146]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2146]->out) 0
.nodeset V(sram[2146]->outb) vsp
Xsram[2147] sram->in sram[2147]->out sram[2147]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2147]->out) 0
.nodeset V(sram[2147]->outb) vsp
Xsram[2148] sram->in sram[2148]->out sram[2148]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2148]->out) 0
.nodeset V(sram[2148]->outb) vsp
Xsram[2149] sram->in sram[2149]->out sram[2149]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2149]->out) 0
.nodeset V(sram[2149]->outb) vsp
Xsram[2150] sram->in sram[2150]->out sram[2150]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2150]->out) 0
.nodeset V(sram[2150]->outb) vsp
Xsram[2151] sram->in sram[2151]->out sram[2151]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2151]->out) 0
.nodeset V(sram[2151]->outb) vsp
Xsram[2152] sram->in sram[2152]->out sram[2152]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2152]->out) 0
.nodeset V(sram[2152]->outb) vsp
Xsram[2153] sram->in sram[2153]->out sram[2153]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2153]->out) 0
.nodeset V(sram[2153]->outb) vsp
Xmux_2level_tapbuf_size16[9] chanx[1][0]_midout[10] chanx[1][0]_midout[11] chanx[1][0]_midout[24] chanx[1][0]_midout[25] chanx[1][0]_midout[36] chanx[1][0]_midout[37] chanx[1][0]_midout[48] chanx[1][0]_midout[49] chanx[1][0]_midout[60] chanx[1][0]_midout[61] chanx[1][0]_midout[74] chanx[1][0]_midout[75] chanx[1][0]_midout[86] chanx[1][0]_midout[87] chanx[1][0]_midout[98] chanx[1][0]_midout[99] grid[1][1]_pin[0][2][38] sram[2154]->outb sram[2154]->out sram[2155]->out sram[2155]->outb sram[2156]->out sram[2156]->outb sram[2157]->out sram[2157]->outb sram[2158]->outb sram[2158]->out sram[2159]->out sram[2159]->outb sram[2160]->out sram[2160]->outb sram[2161]->out sram[2161]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[9], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2154] sram->in sram[2154]->out sram[2154]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2154]->out) 0
.nodeset V(sram[2154]->outb) vsp
Xsram[2155] sram->in sram[2155]->out sram[2155]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2155]->out) 0
.nodeset V(sram[2155]->outb) vsp
Xsram[2156] sram->in sram[2156]->out sram[2156]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2156]->out) 0
.nodeset V(sram[2156]->outb) vsp
Xsram[2157] sram->in sram[2157]->out sram[2157]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2157]->out) 0
.nodeset V(sram[2157]->outb) vsp
Xsram[2158] sram->in sram[2158]->out sram[2158]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2158]->out) 0
.nodeset V(sram[2158]->outb) vsp
Xsram[2159] sram->in sram[2159]->out sram[2159]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2159]->out) 0
.nodeset V(sram[2159]->outb) vsp
Xsram[2160] sram->in sram[2160]->out sram[2160]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2160]->out) 0
.nodeset V(sram[2160]->outb) vsp
Xsram[2161] sram->in sram[2161]->out sram[2161]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2161]->out) 0
.nodeset V(sram[2161]->outb) vsp
Xmux_2level_tapbuf_size16[10] chanx[1][0]_midout[0] chanx[1][0]_midout[1] chanx[1][0]_midout[12] chanx[1][0]_midout[13] chanx[1][0]_midout[24] chanx[1][0]_midout[25] chanx[1][0]_midout[36] chanx[1][0]_midout[37] chanx[1][0]_midout[50] chanx[1][0]_midout[51] chanx[1][0]_midout[62] chanx[1][0]_midout[63] chanx[1][0]_midout[74] chanx[1][0]_midout[75] chanx[1][0]_midout[86] chanx[1][0]_midout[87] grid[1][0]_pin[0][0][0] sram[2162]->outb sram[2162]->out sram[2163]->out sram[2163]->outb sram[2164]->out sram[2164]->outb sram[2165]->out sram[2165]->outb sram[2166]->outb sram[2166]->out sram[2167]->out sram[2167]->outb sram[2168]->out sram[2168]->outb sram[2169]->out sram[2169]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[10], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2162] sram->in sram[2162]->out sram[2162]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2162]->out) 0
.nodeset V(sram[2162]->outb) vsp
Xsram[2163] sram->in sram[2163]->out sram[2163]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2163]->out) 0
.nodeset V(sram[2163]->outb) vsp
Xsram[2164] sram->in sram[2164]->out sram[2164]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2164]->out) 0
.nodeset V(sram[2164]->outb) vsp
Xsram[2165] sram->in sram[2165]->out sram[2165]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2165]->out) 0
.nodeset V(sram[2165]->outb) vsp
Xsram[2166] sram->in sram[2166]->out sram[2166]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2166]->out) 0
.nodeset V(sram[2166]->outb) vsp
Xsram[2167] sram->in sram[2167]->out sram[2167]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2167]->out) 0
.nodeset V(sram[2167]->outb) vsp
Xsram[2168] sram->in sram[2168]->out sram[2168]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2168]->out) 0
.nodeset V(sram[2168]->outb) vsp
Xsram[2169] sram->in sram[2169]->out sram[2169]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2169]->out) 0
.nodeset V(sram[2169]->outb) vsp
Xmux_2level_tapbuf_size16[11] chanx[1][0]_midout[0] chanx[1][0]_midout[1] chanx[1][0]_midout[14] chanx[1][0]_midout[15] chanx[1][0]_midout[26] chanx[1][0]_midout[27] chanx[1][0]_midout[38] chanx[1][0]_midout[39] chanx[1][0]_midout[50] chanx[1][0]_midout[51] chanx[1][0]_midout[64] chanx[1][0]_midout[65] chanx[1][0]_midout[76] chanx[1][0]_midout[77] chanx[1][0]_midout[88] chanx[1][0]_midout[89] grid[1][0]_pin[0][0][2] sram[2170]->outb sram[2170]->out sram[2171]->out sram[2171]->outb sram[2172]->out sram[2172]->outb sram[2173]->out sram[2173]->outb sram[2174]->outb sram[2174]->out sram[2175]->out sram[2175]->outb sram[2176]->out sram[2176]->outb sram[2177]->out sram[2177]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[11], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2170] sram->in sram[2170]->out sram[2170]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2170]->out) 0
.nodeset V(sram[2170]->outb) vsp
Xsram[2171] sram->in sram[2171]->out sram[2171]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2171]->out) 0
.nodeset V(sram[2171]->outb) vsp
Xsram[2172] sram->in sram[2172]->out sram[2172]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2172]->out) 0
.nodeset V(sram[2172]->outb) vsp
Xsram[2173] sram->in sram[2173]->out sram[2173]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2173]->out) 0
.nodeset V(sram[2173]->outb) vsp
Xsram[2174] sram->in sram[2174]->out sram[2174]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2174]->out) 0
.nodeset V(sram[2174]->outb) vsp
Xsram[2175] sram->in sram[2175]->out sram[2175]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2175]->out) 0
.nodeset V(sram[2175]->outb) vsp
Xsram[2176] sram->in sram[2176]->out sram[2176]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2176]->out) 0
.nodeset V(sram[2176]->outb) vsp
Xsram[2177] sram->in sram[2177]->out sram[2177]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2177]->out) 0
.nodeset V(sram[2177]->outb) vsp
Xmux_2level_tapbuf_size16[12] chanx[1][0]_midout[2] chanx[1][0]_midout[3] chanx[1][0]_midout[14] chanx[1][0]_midout[15] chanx[1][0]_midout[28] chanx[1][0]_midout[29] chanx[1][0]_midout[40] chanx[1][0]_midout[41] chanx[1][0]_midout[52] chanx[1][0]_midout[53] chanx[1][0]_midout[64] chanx[1][0]_midout[65] chanx[1][0]_midout[78] chanx[1][0]_midout[79] chanx[1][0]_midout[90] chanx[1][0]_midout[91] grid[1][0]_pin[0][0][4] sram[2178]->outb sram[2178]->out sram[2179]->out sram[2179]->outb sram[2180]->out sram[2180]->outb sram[2181]->out sram[2181]->outb sram[2182]->outb sram[2182]->out sram[2183]->out sram[2183]->outb sram[2184]->out sram[2184]->outb sram[2185]->out sram[2185]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[12], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2178] sram->in sram[2178]->out sram[2178]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2178]->out) 0
.nodeset V(sram[2178]->outb) vsp
Xsram[2179] sram->in sram[2179]->out sram[2179]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2179]->out) 0
.nodeset V(sram[2179]->outb) vsp
Xsram[2180] sram->in sram[2180]->out sram[2180]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2180]->out) 0
.nodeset V(sram[2180]->outb) vsp
Xsram[2181] sram->in sram[2181]->out sram[2181]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2181]->out) 0
.nodeset V(sram[2181]->outb) vsp
Xsram[2182] sram->in sram[2182]->out sram[2182]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2182]->out) 0
.nodeset V(sram[2182]->outb) vsp
Xsram[2183] sram->in sram[2183]->out sram[2183]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2183]->out) 0
.nodeset V(sram[2183]->outb) vsp
Xsram[2184] sram->in sram[2184]->out sram[2184]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2184]->out) 0
.nodeset V(sram[2184]->outb) vsp
Xsram[2185] sram->in sram[2185]->out sram[2185]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2185]->out) 0
.nodeset V(sram[2185]->outb) vsp
Xmux_2level_tapbuf_size16[13] chanx[1][0]_midout[4] chanx[1][0]_midout[5] chanx[1][0]_midout[16] chanx[1][0]_midout[17] chanx[1][0]_midout[28] chanx[1][0]_midout[29] chanx[1][0]_midout[42] chanx[1][0]_midout[43] chanx[1][0]_midout[54] chanx[1][0]_midout[55] chanx[1][0]_midout[66] chanx[1][0]_midout[67] chanx[1][0]_midout[78] chanx[1][0]_midout[79] chanx[1][0]_midout[92] chanx[1][0]_midout[93] grid[1][0]_pin[0][0][6] sram[2186]->outb sram[2186]->out sram[2187]->out sram[2187]->outb sram[2188]->out sram[2188]->outb sram[2189]->out sram[2189]->outb sram[2190]->outb sram[2190]->out sram[2191]->out sram[2191]->outb sram[2192]->out sram[2192]->outb sram[2193]->out sram[2193]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[13], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2186] sram->in sram[2186]->out sram[2186]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2186]->out) 0
.nodeset V(sram[2186]->outb) vsp
Xsram[2187] sram->in sram[2187]->out sram[2187]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2187]->out) 0
.nodeset V(sram[2187]->outb) vsp
Xsram[2188] sram->in sram[2188]->out sram[2188]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2188]->out) 0
.nodeset V(sram[2188]->outb) vsp
Xsram[2189] sram->in sram[2189]->out sram[2189]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2189]->out) 0
.nodeset V(sram[2189]->outb) vsp
Xsram[2190] sram->in sram[2190]->out sram[2190]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2190]->out) 0
.nodeset V(sram[2190]->outb) vsp
Xsram[2191] sram->in sram[2191]->out sram[2191]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2191]->out) 0
.nodeset V(sram[2191]->outb) vsp
Xsram[2192] sram->in sram[2192]->out sram[2192]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2192]->out) 0
.nodeset V(sram[2192]->outb) vsp
Xsram[2193] sram->in sram[2193]->out sram[2193]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2193]->out) 0
.nodeset V(sram[2193]->outb) vsp
Xmux_2level_tapbuf_size16[14] chanx[1][0]_midout[6] chanx[1][0]_midout[7] chanx[1][0]_midout[18] chanx[1][0]_midout[19] chanx[1][0]_midout[30] chanx[1][0]_midout[31] chanx[1][0]_midout[42] chanx[1][0]_midout[43] chanx[1][0]_midout[56] chanx[1][0]_midout[57] chanx[1][0]_midout[68] chanx[1][0]_midout[69] chanx[1][0]_midout[80] chanx[1][0]_midout[81] chanx[1][0]_midout[92] chanx[1][0]_midout[93] grid[1][0]_pin[0][0][8] sram[2194]->outb sram[2194]->out sram[2195]->out sram[2195]->outb sram[2196]->out sram[2196]->outb sram[2197]->out sram[2197]->outb sram[2198]->outb sram[2198]->out sram[2199]->out sram[2199]->outb sram[2200]->out sram[2200]->outb sram[2201]->out sram[2201]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[14], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2194] sram->in sram[2194]->out sram[2194]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2194]->out) 0
.nodeset V(sram[2194]->outb) vsp
Xsram[2195] sram->in sram[2195]->out sram[2195]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2195]->out) 0
.nodeset V(sram[2195]->outb) vsp
Xsram[2196] sram->in sram[2196]->out sram[2196]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2196]->out) 0
.nodeset V(sram[2196]->outb) vsp
Xsram[2197] sram->in sram[2197]->out sram[2197]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2197]->out) 0
.nodeset V(sram[2197]->outb) vsp
Xsram[2198] sram->in sram[2198]->out sram[2198]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2198]->out) 0
.nodeset V(sram[2198]->outb) vsp
Xsram[2199] sram->in sram[2199]->out sram[2199]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2199]->out) 0
.nodeset V(sram[2199]->outb) vsp
Xsram[2200] sram->in sram[2200]->out sram[2200]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2200]->out) 0
.nodeset V(sram[2200]->outb) vsp
Xsram[2201] sram->in sram[2201]->out sram[2201]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2201]->out) 0
.nodeset V(sram[2201]->outb) vsp
Xmux_2level_tapbuf_size16[15] chanx[1][0]_midout[6] chanx[1][0]_midout[7] chanx[1][0]_midout[20] chanx[1][0]_midout[21] chanx[1][0]_midout[32] chanx[1][0]_midout[33] chanx[1][0]_midout[44] chanx[1][0]_midout[45] chanx[1][0]_midout[56] chanx[1][0]_midout[57] chanx[1][0]_midout[70] chanx[1][0]_midout[71] chanx[1][0]_midout[82] chanx[1][0]_midout[83] chanx[1][0]_midout[94] chanx[1][0]_midout[95] grid[1][0]_pin[0][0][10] sram[2202]->outb sram[2202]->out sram[2203]->out sram[2203]->outb sram[2204]->out sram[2204]->outb sram[2205]->out sram[2205]->outb sram[2206]->outb sram[2206]->out sram[2207]->out sram[2207]->outb sram[2208]->out sram[2208]->outb sram[2209]->out sram[2209]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[15], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2202] sram->in sram[2202]->out sram[2202]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2202]->out) 0
.nodeset V(sram[2202]->outb) vsp
Xsram[2203] sram->in sram[2203]->out sram[2203]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2203]->out) 0
.nodeset V(sram[2203]->outb) vsp
Xsram[2204] sram->in sram[2204]->out sram[2204]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2204]->out) 0
.nodeset V(sram[2204]->outb) vsp
Xsram[2205] sram->in sram[2205]->out sram[2205]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2205]->out) 0
.nodeset V(sram[2205]->outb) vsp
Xsram[2206] sram->in sram[2206]->out sram[2206]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2206]->out) 0
.nodeset V(sram[2206]->outb) vsp
Xsram[2207] sram->in sram[2207]->out sram[2207]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2207]->out) 0
.nodeset V(sram[2207]->outb) vsp
Xsram[2208] sram->in sram[2208]->out sram[2208]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2208]->out) 0
.nodeset V(sram[2208]->outb) vsp
Xsram[2209] sram->in sram[2209]->out sram[2209]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2209]->out) 0
.nodeset V(sram[2209]->outb) vsp
Xmux_2level_tapbuf_size16[16] chanx[1][0]_midout[8] chanx[1][0]_midout[9] chanx[1][0]_midout[20] chanx[1][0]_midout[21] chanx[1][0]_midout[34] chanx[1][0]_midout[35] chanx[1][0]_midout[46] chanx[1][0]_midout[47] chanx[1][0]_midout[58] chanx[1][0]_midout[59] chanx[1][0]_midout[70] chanx[1][0]_midout[71] chanx[1][0]_midout[84] chanx[1][0]_midout[85] chanx[1][0]_midout[96] chanx[1][0]_midout[97] grid[1][0]_pin[0][0][12] sram[2210]->outb sram[2210]->out sram[2211]->out sram[2211]->outb sram[2212]->out sram[2212]->outb sram[2213]->out sram[2213]->outb sram[2214]->outb sram[2214]->out sram[2215]->out sram[2215]->outb sram[2216]->out sram[2216]->outb sram[2217]->out sram[2217]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[16], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2210] sram->in sram[2210]->out sram[2210]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2210]->out) 0
.nodeset V(sram[2210]->outb) vsp
Xsram[2211] sram->in sram[2211]->out sram[2211]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2211]->out) 0
.nodeset V(sram[2211]->outb) vsp
Xsram[2212] sram->in sram[2212]->out sram[2212]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2212]->out) 0
.nodeset V(sram[2212]->outb) vsp
Xsram[2213] sram->in sram[2213]->out sram[2213]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2213]->out) 0
.nodeset V(sram[2213]->outb) vsp
Xsram[2214] sram->in sram[2214]->out sram[2214]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2214]->out) 0
.nodeset V(sram[2214]->outb) vsp
Xsram[2215] sram->in sram[2215]->out sram[2215]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2215]->out) 0
.nodeset V(sram[2215]->outb) vsp
Xsram[2216] sram->in sram[2216]->out sram[2216]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2216]->out) 0
.nodeset V(sram[2216]->outb) vsp
Xsram[2217] sram->in sram[2217]->out sram[2217]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2217]->out) 0
.nodeset V(sram[2217]->outb) vsp
Xmux_2level_tapbuf_size16[17] chanx[1][0]_midout[10] chanx[1][0]_midout[11] chanx[1][0]_midout[22] chanx[1][0]_midout[23] chanx[1][0]_midout[34] chanx[1][0]_midout[35] chanx[1][0]_midout[48] chanx[1][0]_midout[49] chanx[1][0]_midout[60] chanx[1][0]_midout[61] chanx[1][0]_midout[72] chanx[1][0]_midout[73] chanx[1][0]_midout[84] chanx[1][0]_midout[85] chanx[1][0]_midout[98] chanx[1][0]_midout[99] grid[1][0]_pin[0][0][14] sram[2218]->outb sram[2218]->out sram[2219]->out sram[2219]->outb sram[2220]->out sram[2220]->outb sram[2221]->out sram[2221]->outb sram[2222]->outb sram[2222]->out sram[2223]->out sram[2223]->outb sram[2224]->out sram[2224]->outb sram[2225]->out sram[2225]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[17], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2218] sram->in sram[2218]->out sram[2218]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2218]->out) 0
.nodeset V(sram[2218]->outb) vsp
Xsram[2219] sram->in sram[2219]->out sram[2219]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2219]->out) 0
.nodeset V(sram[2219]->outb) vsp
Xsram[2220] sram->in sram[2220]->out sram[2220]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2220]->out) 0
.nodeset V(sram[2220]->outb) vsp
Xsram[2221] sram->in sram[2221]->out sram[2221]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2221]->out) 0
.nodeset V(sram[2221]->outb) vsp
Xsram[2222] sram->in sram[2222]->out sram[2222]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2222]->out) 0
.nodeset V(sram[2222]->outb) vsp
Xsram[2223] sram->in sram[2223]->out sram[2223]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2223]->out) 0
.nodeset V(sram[2223]->outb) vsp
Xsram[2224] sram->in sram[2224]->out sram[2224]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2224]->out) 0
.nodeset V(sram[2224]->outb) vsp
Xsram[2225] sram->in sram[2225]->out sram[2225]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2225]->out) 0
.nodeset V(sram[2225]->outb) vsp
.eom
