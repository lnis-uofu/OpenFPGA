// Benchmark "TOP" written by ABC on Mon Feb  4 17:25:42 2019

module apex4 ( 
    i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_,
    o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_,
    o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_  );
  input  i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;
  output o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_,
    o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_;
  wire n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
    n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
    n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
    n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
    n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
    n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
    n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
    n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
    n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
    n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
    n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
    n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
    n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
    n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
    n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
    n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
    n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
    n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
    n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
    n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
    n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
    n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
    n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
    n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
    n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
    n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
    n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749;
  assign o_0_ = 1'b0;
  assign o_1_ = ~n134;
  assign o_2_ = ~n492;
  assign o_3_ = ~n129;
  assign o_4_ = ~n128;
  assign o_5_ = ~n119;
  assign o_6_ = ~n110;
  assign o_7_ = ~n101;
  assign o_8_ = ~n313;
  assign o_9_ = ~n100;
  assign o_10_ = ~n526;
  assign o_11_ = ~n91;
  assign o_12_ = ~n87;
  assign o_13_ = ~n80;
  assign o_14_ = ~n72;
  assign o_15_ = ~n64;
  assign o_16_ = ~n63;
  assign o_17_ = ~n61;
  assign o_18_ = ~n53;
  assign n47 = n440 | n512;
  assign n48 = n539 | n454;
  assign n49 = n425 | n540;
  assign n50 = n305 | n557;
  assign n51 = n643 & n644 & n409 & n616 & n645 & n646 & n642 & n647;
  assign n52 = n65 & (n515 | n514);
  assign n53 = n47 & n48 & n49 & n50 & n51 & n52;
  assign n54 = n641 & n501 & n624 & n620 & n586;
  assign n55 = n314 | n591;
  assign n56 = n528 | n208;
  assign n57 = n425 | n558;
  assign n58 = n236 | n576;
  assign n59 = n545 | ~i_6_ | n531;
  assign n60 = n49 & n742;
  assign n61 = n48 & n54 & n55 & n56 & n57 & n58 & n59 & n60;
  assign n62 = n651 & n652 & n653 & n654 & n650 & n259 & n604 & n655;
  assign n63 = n54 & n62 & n50 & n47;
  assign n64 = n51 & n62 & n58 & n56;
  assign n65 = n190 | n543 | n514;
  assign n66 = n229 | n548;
  assign n67 = n443 | ~i_0_ | n419;
  assign n68 = n190 | n562;
  assign n69 = n656 & n247 & n657 & n621 & n658 & n599 & n659;
  assign n70 = n437 & n456 & n513 & n660 & n661 & n516 & n662 & n663;
  assign n71 = n504 & n505 & n506 & n507 & n508 & n509 & n510 & n511;
  assign n72 = n65 & n66 & n67 & n68 & n69 & n70 & n71;
  assign n73 = n664 & n597 & n556 & n264 & n358 & n391 & n434 & ~n522;
  assign n74 = n360 & n517 & n399 & n518 & n519 & n520 & n521;
  assign n75 = n515 | n245;
  assign n76 = n440 | n558;
  assign n77 = ~i_0_ | n190 | n250 | n252;
  assign n78 = n430 | n419;
  assign n79 = ~n332 | n345;
  assign n80 = n73 & n74 & n75 & n70 & n76 & n77 & n78 & n79;
  assign n81 = n634 & n596 & n350 & n468 & n130 & n665 & n666 & n667;
  assign n82 = n440 | n144;
  assign n83 = i_3_ | n373 | n419;
  assign n84 = n190 | n575;
  assign n85 = n342 | n559;
  assign n86 = n182 | n575;
  assign n87 = n74 & n81 & n82 & n69 & n83 & n84 & n85 & n86;
  assign n88 = n560 | n575;
  assign n89 = ~i_3_ | i_5_ | n440 | ~n461;
  assign n90 = n345 | ~i_0_ | n250;
  assign n91 = n88 & n89 & n59 & n90 & n71 & n73 & n81;
  assign n92 = n570 & n193 & n202 & n199 & n588 & n589;
  assign n93 = n178 & n184 & n183 & n185 & n186 & n187 & n188 & n189;
  assign n94 = n141 & n155 & n160 & n164 & n172 & n122 & n173 & n174;
  assign n95 = n221 & n222 & (n223 | n224);
  assign n96 = n213 & n214 & n215 & n216 & n217 & n218 & n219 & n220;
  assign n97 = n210 & n206 & n583 & n212 & n584 & n585 & n586 & n587;
  assign n98 = n582 & n580 & ~n255 & n123 & n238 & n249 & ~n254;
  assign n99 = n660 & n685 & n615 & n686 & n687 & n325 & n253 & n684;
  assign n100 = n92 & n93 & n94 & n95 & n96 & n97 & n98 & n99;
  assign n101 = n102 & n348 & n349 & n347 & n350 & n351 & n352 & n353;
  assign n102 = n325 & n326 & n152 & n327 & n328 & n329 & n330 & n331;
  assign n103 = n371 & (i_5_ | n372);
  assign n104 = n369 & (n190 | n223 | n370);
  assign n105 = n630 & n366 & n368 & n149 & n216 & n631;
  assign n106 = n151 & n358 & n359 & n360 & n361 & n362 & n363 & n364;
  assign n107 = n580 & n379 & n210 & n267 & n285 & ~n377;
  assign n108 = n90 & n417 & n712 & n148 & n568 & n713;
  assign n109 = n646 & n66 & n75 & n86 & n374 & ~n376;
  assign n110 = n102 & n103 & n104 & n105 & n106 & n107 & n108 & n109;
  assign n111 = n414 & (n415 | n416);
  assign n112 = n281 & n413 & (n224 | ~n332);
  assign n113 = n407 & n79 & n408 & n409 & n49 & n410 & n411 & n412;
  assign n114 = n399 & n400 & n401 & n402 & n403 & n404 & n405 & n406;
  assign n115 = n391 & n392 & n393 & n394 & n395 & n396 & n397 & n398;
  assign n116 = n349 & n424 & n420 & n431 & n94 & n307;
  assign n117 = n638 & n656 & n713 & n694 & n57 & n651;
  assign n118 = n427 & n428 & n429 & n614 & n86 & n696;
  assign n119 = n111 & n112 & n113 & n114 & n115 & n116 & n117 & n118;
  assign n120 = n262 & n266 & n267 & n268 & n269 & n270 & n271 & n272;
  assign n121 = n315 & n202 & n613 & n614;
  assign n122 = n168 & n169 & (n170 | n171);
  assign n123 = n88 & n231 & (n232 | n233);
  assign n124 = n240 | n415 | i_0_ | ~i_2_;
  assign n125 = n443 | n190 | n444;
  assign n126 = n500 & n719 & n720;
  assign n127 = n435 & n457 & n442 & n437 & n386 & n111 & n348 & n106;
  assign n128 = n120 & n121 & n122 & n123 & n124 & n125 & n126 & n127;
  assign n129 = n447 & n456 & n455 & n457 & n115 & n347 & n458 & n459;
  assign n130 = n382 & n496 & (n145 | n335);
  assign n131 = n640 & n494 & n495 & n505 & n504 & n619;
  assign n132 = n661 & n657 & n497;
  assign n133 = n603 & n48 & n68 & n720 & n279 & n187 & n602 & n741;
  assign n134 = ~n499 & n97 & n112 & n130 & n131 & n132 & n133 & ~n498;
  assign n135 = n339 | n542;
  assign n136 = n440 | n416;
  assign n137 = n166 | n541;
  assign n138 = n236 | n538;
  assign n139 = (n440 | n237) & (n305 | n224);
  assign n140 = n679 & (n301 | n226 | n515);
  assign n141 = n135 & n136 & n137 & n138 & n139 & n140;
  assign n142 = n301 | n354 | n474;
  assign n143 = n166 | n341;
  assign n144 = n430 | n158;
  assign n145 = i_6_ | i_7_;
  assign n146 = n142 & n143 & (n144 | n145);
  assign n147 = n422 | n467;
  assign n148 = n170 | n544;
  assign n149 = n342 | n367;
  assign n150 = n440 | n436;
  assign n151 = n166 | n365;
  assign n152 = ~i_6_ | ~i_8_ | n453;
  assign n153 = n422 | n546;
  assign n154 = n146 & (n440 | n232 | n430);
  assign n155 = n147 & n148 & n149 & n150 & n151 & n152 & n153 & n154;
  assign n156 = n425 | n448;
  assign n157 = n229 | n252 | n226;
  assign n158 = i_5_ | n533;
  assign n159 = n182 | ~n332;
  assign n160 = n156 & n157 & (n158 | n159);
  assign n161 = n529 | n548;
  assign n162 = n425 | n546;
  assign n163 = (n440 | n534) & (n423 | n454);
  assign n164 = n161 & n162 & n163;
  assign n165 = n182 | n430;
  assign n166 = i_5_ | n240;
  assign n167 = n165 | n166;
  assign n168 = n240 | n223 | n208;
  assign n169 = n342 | n337;
  assign n170 = ~i_5_ | n533;
  assign n171 = n425 | n430;
  assign n172 = n553 & n554 & n167 & n286 & n555 & n556;
  assign n173 = n683 & n477 & (n425 | n195);
  assign n174 = n633 & n482 & n637 & n609 & n681 & n682 & n621 & n680;
  assign n175 = n454 | n463;
  assign n176 = n236 | n209;
  assign n177 = (n166 | n559) & (n158 | n341);
  assign n178 = n175 & n176 & n177;
  assign n179 = n560 | n441;
  assign n180 = n531 | n224;
  assign n181 = n166 | n305;
  assign n182 = ~i_6_ | n529;
  assign n183 = n179 & n180 & (n181 | n182);
  assign n184 = n295 & n294 & n563;
  assign n185 = n166 | n367;
  assign n186 = n529 | n531 | n472;
  assign n187 = n225 | n301 | ~n332;
  assign n188 = n678 & (~i_8_ | n562);
  assign n189 = n675 & n676 & n269 & n76 & n362 & n624 & n677 & n50;
  assign n190 = i_7_ | i_8_;
  assign n191 = ~i_6_ | n543;
  assign n192 = ~i_0_ | ~n469;
  assign n193 = n85 & (n190 | n191 | n192);
  assign n194 = i_6_ | ~i_7_;
  assign n195 = n166 | n223;
  assign n196 = n194 | n195;
  assign n197 = n416 | n454;
  assign n198 = n232 | n223;
  assign n199 = n197 & (n198 | n145);
  assign n200 = n166 | n566;
  assign n201 = n339 | n274;
  assign n202 = n200 & n201 & (n182 | n144);
  assign n203 = n166 | n337;
  assign n204 = n425 | n209;
  assign n205 = (n158 | n233) & (n198 | n454);
  assign n206 = n203 & n204 & n205;
  assign n207 = n145 | n170 | ~n461;
  assign n208 = ~i_6_ | n229;
  assign n209 = n241 | n545;
  assign n210 = n207 & (n208 | n209);
  assign n211 = n223 | n339;
  assign n212 = n211 | n208;
  assign n213 = n440 | n209;
  assign n214 = n158 | n274;
  assign n215 = n236 | n572;
  assign n216 = n182 | n572;
  assign n217 = n415 | n211;
  assign n218 = n301 | n191 | n488;
  assign n219 = n182 | n211;
  assign n220 = (n166 | n573) & (n532 | n145);
  assign n221 = n531 | n229 | n545;
  assign n222 = n59 & (n232 | ~n332 | n574);
  assign n223 = ~i_2_ | n321;
  assign n224 = n425 | n339;
  assign n225 = i_6_ | n487;
  assign n226 = ~i_1_ | n443;
  assign n227 = n226 | ~i_7_ | n225;
  assign n228 = i_0_ | n191 | ~n469;
  assign n229 = ~i_7_ | ~i_8_;
  assign n230 = n228 | n229;
  assign n231 = n422 | n195;
  assign n232 = ~i_5_ | n240;
  assign n233 = n182 | ~n461;
  assign n234 = n190 | n515 | n488;
  assign n235 = n342 | n372;
  assign n236 = i_6_ | n529;
  assign n237 = n531 | n158;
  assign n238 = n234 & n235 & (n236 | n237);
  assign n239 = n321 | n577;
  assign n240 = ~i_3_ | i_4_;
  assign n241 = ~i_2_ | n373;
  assign n242 = ~i_6_ | i_8_;
  assign n243 = n239 & (n240 | n241 | n242);
  assign n244 = i_6_ | n323;
  assign n245 = n190 | ~n461;
  assign n246 = n244 | n245;
  assign n247 = n339 | n573;
  assign n248 = i_3_ | i_4_ | i_6_;
  assign n249 = n247 & (n229 | n248 | ~n332);
  assign n250 = i_2_ | ~i_3_;
  assign n251 = n250 | ~i_0_ | n225;
  assign n252 = i_6_ | ~i_4_ | i_5_;
  assign n253 = ~i_1_ | ~i_7_ | n250 | n252;
  assign n254 = i_8_ & (~n251 | (~n430 & ~n472));
  assign n255 = ~i_5_ & (~n591 | (~n422 & ~n561));
  assign n256 = n425 | n436;
  assign n257 = n378 | ~n461;
  assign n258 = n170 | n367;
  assign n259 = n208 | n558;
  assign n260 = n327 & (n166 | n229 | ~n461);
  assign n261 = n301 | n144;
  assign n262 = n256 & n257 & n258 & n259 & n260 & n261;
  assign n263 = n415 | n538;
  assign n264 = n181 | n208;
  assign n265 = n578 & (n301 | n241 | n444);
  assign n266 = n78 & n263 & n264 & n265;
  assign n267 = n592 & n593;
  assign n268 = n238 & n700 & (n537 | n191);
  assign n269 = n339 | n440 | ~n461;
  assign n270 = n342 | n365;
  assign n271 = n232 | n241 | n242;
  assign n272 = n669 & n699 & n656 & n410;
  assign n273 = ~n415 & (~n237 | (~n305 & ~n533));
  assign n274 = n208 | ~n332;
  assign n275 = n274 | n170;
  assign n276 = n444 | n565;
  assign n277 = n365 | ~i_4_ | i_5_;
  assign n278 = n276 & n277 & (n225 | n245);
  assign n279 = n232 | n372;
  assign n280 = n529 | n571;
  assign n281 = n342 | n159;
  assign n282 = n182 | n539;
  assign n283 = n691 & (n527 | n544);
  assign n284 = n689 & n466 & n690 & n658 & n452 & n648 & n138 & n402;
  assign n285 = n279 & n280 & n281 & n282 & n183 & n146 & n283 & n284;
  assign n286 = n545 | n274;
  assign n287 = n158 | n542;
  assign n288 = n532 | n425;
  assign n289 = n425 | n453;
  assign n290 = n170 | n302 | n430;
  assign n291 = n182 | n423;
  assign n292 = (n532 | n454) & (n528 | n145);
  assign n293 = n286 & n136 & n287 & n288 & n289 & n290 & n291 & n292;
  assign n294 = n208 | n546;
  assign n295 = n440 | n493;
  assign n296 = n236 | n564;
  assign n297 = n158 | n591;
  assign n298 = n688 & (n158 | n236 | ~n332);
  assign n299 = n305 | n229 | n354;
  assign n300 = n294 & n295 & n296 & n297 & n298 & n299;
  assign n301 = ~i_7_ | i_8_;
  assign n302 = i_6_ | ~i_8_;
  assign n303 = n531 | n339;
  assign n304 = (n301 | n228) & (n302 | n303);
  assign n305 = i_2_ | n321;
  assign n306 = i_3_ | i_5_;
  assign n307 = n239 & (n305 | n236 | n306);
  assign n308 = n602 & n603 & n604 & n519;
  assign n309 = n702 & (~i_1_ | n182 | n342);
  assign n310 = n351 & n285 & n120 & n300 & n304 & n293;
  assign n311 = n673 & n84 & n640 & n675 & n701 & n67;
  assign n312 = n76 & n404 & n219 & n636 & n649 & n79;
  assign n313 = n308 & n95 & n307 & n309 & n160 & n310 & n311 & n312;
  assign n314 = i_3_ | n487;
  assign n315 = n159 | n314;
  assign n316 = n165 | n232;
  assign n317 = n440 | n423;
  assign n318 = n190 | n248 | ~n332;
  assign n319 = (n236 | n536) & (n415 | n575);
  assign n320 = n317 & n318 & n319;
  assign n321 = i_0_ | ~i_1_;
  assign n322 = n191 | n301 | n321 | i_3_;
  assign n323 = i_3_ | ~i_5_;
  assign n324 = n208 | n223 | n323;
  assign n325 = n537 | n252;
  assign n326 = n415 | n467;
  assign n327 = n342 | n573;
  assign n328 = n706 & (i_0_ | n443 | n419);
  assign n329 = i_3_ | n566;
  assign n330 = n320 & n478 & n300 & n172 & n121 & n612 & n617;
  assign n331 = n705 & n218 & n403 & n257 & n150 & n187 & n583 & n704;
  assign n332 = ~i_2_ & ~n426;
  assign n333 = ~n170 & (~n233 | (~n301 & n332));
  assign n334 = ~n430 & (~n224 | (~n314 & ~n529));
  assign n335 = n342 | n241;
  assign n336 = n335 | n190;
  assign n337 = ~n332 | n422;
  assign n338 = n337 | n232;
  assign n339 = i_5_ | n527;
  assign n340 = n242 | n339 | ~n461;
  assign n341 = n415 | ~n461;
  assign n342 = ~i_5_ | n527;
  assign n343 = n341 | n342;
  assign n344 = n681 & n563 & n703;
  assign n345 = n229 | n444;
  assign n346 = i_1_ | ~n469;
  assign n347 = n243 & n344 & (n345 | n346);
  assign n348 = n621 & n622 & n623 & n624 & n496 & n625 & n626 & n627;
  assign n349 = n340 & n343 & n58 & n620;
  assign n350 = n618 & n405 & n619;
  assign n351 = n605 & n178 & n606 & n607 & n278 & n596 & n601 & n608;
  assign n352 = n582 & n193 & n266;
  assign n353 = n399 & n258 & n695 & n708 & n506 & n186 & n654 & n707;
  assign n354 = ~i_6_ | n487;
  assign n355 = n301 | n354 | ~n461;
  assign n356 = ~i_4_ | ~i_5_;
  assign n357 = n356 | n165;
  assign n358 = n182 | n448;
  assign n359 = n241 | n224;
  assign n360 = n232 | n182 | n241;
  assign n361 = n166 | n159;
  assign n362 = n170 | n341;
  assign n363 = n47 & n501 & n147;
  assign n364 = n408 & n396 & n676 & n197 & n710 & n388 & n711 & n709;
  assign n365 = n430 | n208;
  assign n366 = n365 | n232;
  assign n367 = ~n332 | n425;
  assign n368 = n367 | n158;
  assign n369 = n531 | n208 | n547;
  assign n370 = i_6_ | n547;
  assign n371 = n534 | n449;
  assign n372 = n425 | ~n461;
  assign n373 = ~i_0_ | ~i_1_;
  assign n374 = n373 | n301 | n339;
  assign n375 = (i_1_ & (~i_5_ | ~n426)) | (i_5_ & ~n426);
  assign n376 = ~n454 & ~i_4_ & n375;
  assign n377 = ~n195 & (~n425 | ~n449);
  assign n378 = n232 | n236;
  assign n379 = ~n332 | n378;
  assign n380 = n241 | n557;
  assign n381 = n423 | n208;
  assign n382 = n166 | n590;
  assign n383 = n232 | n542;
  assign n384 = (n170 | n541) & (n422 | n453);
  assign n385 = n716 & (~i_1_ | i_2_ | n577);
  assign n386 = n380 & n381 & n382 & n383 & n384 & n385;
  assign n387 = n422 | n549;
  assign n388 = n355 & n357 & n628 & n629;
  assign n389 = n529 | n515;
  assign n390 = n387 & n388 & (n389 | n346);
  assign n391 = n236 | n549;
  assign n392 = n170 | n590;
  assign n393 = n415 | n441;
  assign n394 = n182 | n564;
  assign n395 = n425 | n538;
  assign n396 = n208 | n441;
  assign n397 = n425 | n441;
  assign n398 = n390 & n320 & n386 & n308 & n278 & n718;
  assign n399 = n166 | n430 | n454;
  assign n400 = n170 | n159;
  assign n401 = n314 | n559;
  assign n402 = n425 | n564;
  assign n403 = n144 | n454;
  assign n404 = n314 | n274;
  assign n405 = n538 | n208;
  assign n406 = n326 & n607 & n282 & n697 & n714 & n715;
  assign n407 = n474 | n438;
  assign n408 = n314 | n449 | ~n461;
  assign n409 = n449 | n564;
  assign n410 = n182 | n467;
  assign n411 = n708 & n625 & (n537 | n248);
  assign n412 = n613 & n698 & n710;
  assign n413 = n594 & n693 & n90;
  assign n414 = n301 | n430 | n252;
  assign n415 = i_6_ | n301;
  assign n416 = n305 | n170;
  assign n417 = n415 | n453;
  assign n418 = n425 | n576;
  assign n419 = n225 | n229;
  assign n420 = n417 & n418 & (n192 | n419);
  assign n421 = n574 | ~n332 | n545;
  assign n422 = ~i_6_ | n301;
  assign n423 = n166 | n241;
  assign n424 = n421 & (n422 | n423);
  assign n425 = ~i_6_ | n190;
  assign n426 = ~i_0_ | i_1_;
  assign n427 = n425 | n240 | n426;
  assign n428 = n354 | i_7_ | n192;
  assign n429 = n229 | n241 | n244;
  assign n430 = i_2_ | n373;
  assign n431 = n224 | n430;
  assign n432 = ~n454 & ((~n223 & ~n306) | ~n534);
  assign n433 = n372 | n158;
  assign n434 = n415 | n546;
  assign n435 = n434 & (n229 | ~n332 | n370);
  assign n436 = n223 | n545;
  assign n437 = n401 & (n236 | n436);
  assign n438 = n229 | n515;
  assign n439 = ~i_0_ | ~i_2_;
  assign n440 = i_6_ | n190;
  assign n441 = n223 | n170;
  assign n442 = (n438 | n439) & (n440 | n441);
  assign n443 = ~i_2_ | i_3_;
  assign n444 = i_6_ | n356;
  assign n445 = n208 | n493;
  assign n446 = (n422 | n575) & (n529 | n441);
  assign n447 = n445 & n361 & n446;
  assign n448 = n430 | n545;
  assign n449 = ~i_6_ | ~i_7_;
  assign n450 = n448 | n449;
  assign n451 = n232 | n367;
  assign n452 = n305 | n422 | n533;
  assign n453 = n342 | n223;
  assign n454 = i_6_ | n229;
  assign n455 = n451 & n452 & (n453 | n454);
  assign n456 = n636 & n450 & n622 & n579;
  assign n457 = n635 & n634 & n633 & n632 & n553 & n552 & ~n432 & n433;
  assign n458 = n601 & n249 & n617;
  assign n459 = n294 & n297 & n701 & n721 & n206 & n199 & n722 & n155;
  assign n460 = ~n252 & ~n529;
  assign n461 = i_2_ & ~n426;
  assign n462 = n461 & ((~n194 & ~n314) | n460);
  assign n463 = n305 | n339;
  assign n464 = n463 | n415;
  assign n465 = n182 | n534;
  assign n466 = n314 | n365;
  assign n467 = n241 | n158;
  assign n468 = n465 & n466 & (n236 | n467);
  assign n469 = i_3_ & i_2_;
  assign n470 = n469 & ((~n229 & ~n252) | ~n389);
  assign n471 = ~n470 & (i_2_ | n306 | n440);
  assign n472 = ~i_6_ | n527;
  assign n473 = (n229 | n472) & (i_7_ | n370);
  assign n474 = i_3_ | n426;
  assign n475 = (n321 | n158) & (i_4_ | n474);
  assign n476 = n639 & n638 & n637 & n464 & n148 & ~n462;
  assign n477 = n550 & n551 & n552;
  assign n478 = n291 & n322 & n324;
  assign n479 = n732 & n734 & (~i_1_ | n471);
  assign n480 = n554 & n701 & n731 & n730 & n396 & n161 & n688 & n727;
  assign n481 = n468 & n420 & n476 & n96 & n477 & n478 & n479 & n480;
  assign n482 = n440 | n540;
  assign n483 = n482 & (n198 | n415);
  assign n484 = n302 | n158;
  assign n485 = n166 | n236;
  assign n486 = n484 & n485 & (~i_5_ | n440);
  assign n487 = i_4_ | ~i_5_;
  assign n488 = i_3_ | ~i_0_ | i_2_;
  assign n489 = (n487 | n488) & (n373 | n170);
  assign n490 = n262 & n92 & n612 & n738 & n739 & n737;
  assign n491 = n621 & n649 & n644 & n643 & n289 & n162 & n393 & n736;
  assign n492 = n483 & n447 & n481 & n114 & n103 & n442 & n490 & n491;
  assign n493 = n241 | n314;
  assign n494 = n493 | n422;
  assign n495 = n209 | n182;
  assign n496 = n425 | n493;
  assign n497 = n356 | n182 | n346;
  assign n498 = ~n170 & ~n449 & (~n430 | n461);
  assign n499 = n332 & (~n378 | ~n485 | ~n740);
  assign n500 = n545 | n145 | ~n332;
  assign n501 = n531 | n557;
  assign n502 = (n342 | n171) & (n449 | n335);
  assign n503 = n500 & n501 & n502;
  assign n504 = n166 | n274;
  assign n505 = n158 | n566;
  assign n506 = n422 | n576;
  assign n507 = n719 & (n190 | n354 | n561);
  assign n508 = n430 | n345;
  assign n509 = n476 & n455 & n503 & n293 & n570 & n424;
  assign n510 = n611 & n383 & n203 & n213 & n682 & n361;
  assign n511 = n317 & n176 & n175 & n643 & n641 & n318;
  assign n512 = n166 | n531;
  assign n513 = n270 & (n425 | n512);
  assign n514 = i_3_ | n530;
  assign n515 = i_6_ | n543;
  assign n516 = n514 | n515;
  assign n517 = n145 | n575;
  assign n518 = n166 | n233;
  assign n519 = n170 | n566;
  assign n520 = n669 & n387 & n217 & n693 & n200;
  assign n521 = n404 & n692 & n359 & n744 & n650 & n642 & n483 & n105;
  assign n522 = ~n232 & (~n544 | ~n591);
  assign n523 = n390 & n104 & n113 & n93 & n141 & n304;
  assign n524 = n745 & n746 & n747 & n77 & n381 & n605;
  assign n525 = n689 & n271 & n705 & n360 & n47 & n618;
  assign n526 = n481 & n435 & n131 & n513 & n503 & n523 & n524 & n525;
  assign n527 = i_3_ | ~i_4_;
  assign n528 = n305 | n342;
  assign n529 = i_7_ | ~i_8_;
  assign n530 = i_1_ | i_0_;
  assign n531 = ~i_2_ | n530;
  assign n532 = n342 | n531;
  assign n533 = ~i_3_ | ~i_4_;
  assign n534 = n170 | n241;
  assign n535 = i_0_ | n443 | n225;
  assign n536 = n339 | n430;
  assign n537 = n223 | n229;
  assign n538 = n531 | n170;
  assign n539 = n305 | n158;
  assign n540 = n305 | n314;
  assign n541 = n422 | n430;
  assign n542 = n208 | ~n461;
  assign n543 = i_4_ | i_5_;
  assign n544 = n415 | n430;
  assign n545 = i_4_ | n306;
  assign n546 = n305 | n545;
  assign n547 = ~i_3_ | ~i_5_;
  assign n548 = n430 | n370;
  assign n549 = n223 | n158;
  assign n550 = n232 | n341;
  assign n551 = n170 | n372;
  assign n552 = n208 | n540;
  assign n553 = n182 | n549;
  assign n554 = n208 | n463;
  assign n555 = n540 | n454;
  assign n556 = n425 | n467;
  assign n557 = n422 | n339;
  assign n558 = n531 | n314;
  assign n559 = ~n332 | n454;
  assign n560 = ~i_6_ | i_7_;
  assign n561 = i_1_ | n443;
  assign n562 = n426 | ~i_3_ | n252;
  assign n563 = n236 | n211;
  assign n564 = n305 | n232;
  assign n565 = n529 | n474;
  assign n566 = n422 | ~n461;
  assign n567 = n236 | n463;
  assign n568 = n536 | n560;
  assign n569 = n339 | n341;
  assign n570 = n567 & n196 & n568 & n569;
  assign n571 = n223 | n314;
  assign n572 = n241 | n339;
  assign n573 = ~n332 | n415;
  assign n574 = i_6_ | i_8_;
  assign n575 = ~n461 | n545;
  assign n576 = n232 | n531;
  assign n577 = i_3_ | n190 | n444;
  assign n578 = n49 & n394 & n421 & n387 & n445;
  assign n579 = n440 | n564;
  assign n580 = n246 & n578 & n243 & n410 & n579 & n418;
  assign n581 = ~n461 | n485;
  assign n582 = n227 & n230 & n451 & n581;
  assign n583 = n422 | n441;
  assign n584 = n422 | n571;
  assign n585 = n182 | n546;
  assign n586 = n425 | n416;
  assign n587 = n182 | n436;
  assign n588 = n672 & n673 & n606 & n674;
  assign n589 = n668 & n626 & n669 & n670 & n671 & n287 & n645 & n296;
  assign n590 = ~n332 | n440;
  assign n591 = n182 | n531;
  assign n592 = n407 & n135 & n692 & n392 & n137 & n693 & n694 & n55;
  assign n593 = n695 & n696 & n685 & n687 & n585 & n697 & n698 & n681;
  assign n594 = n339 | n559;
  assign n595 = n181 | n425;
  assign n596 = n418 & n393 & n594 & n595 & n550;
  assign n597 = ~n332 | n557;
  assign n598 = n425 | n144;
  assign n599 = n440 | n571;
  assign n600 = n314 | n541;
  assign n601 = n600 & n599 & n598 & n597 & n518 & ~n273 & n275;
  assign n602 = n182 | n493;
  assign n603 = n232 | n274;
  assign n604 = n422 | n558;
  assign n605 = n170 | n236 | ~n461;
  assign n606 = n430 | n485;
  assign n607 = n208 | n416;
  assign n608 = n551 & n686 & n639 & n637 & n671 & n569 & n57 & n653;
  assign n609 = n339 | n159;
  assign n610 = n422 | n237;
  assign n611 = n237 | n454;
  assign n612 = n609 & n395 & n316 & n610 & n611 & n391;
  assign n613 = n236 | n416;
  assign n614 = n539 | n242;
  assign n615 = n181 | n302;
  assign n616 = n454 | n564;
  assign n617 = n615 & n256 & n269 & n234 & n214 & n270 & n50 & n616;
  assign n618 = n529 | n535;
  assign n619 = n223 | n557;
  assign n620 = n532 | n208;
  assign n621 = n422 | n538;
  assign n622 = n182 | n571;
  assign n623 = n181 | n440;
  assign n624 = n182 | n463;
  assign n625 = n182 | n195;
  assign n626 = n565 | n191;
  assign n627 = n397 & n338 & n336 & ~n334 & n82 & ~n333;
  assign n628 = n425 | n571;
  assign n629 = n342 | n274;
  assign n630 = n236 | n342 | ~n461;
  assign n631 = n534 | n415;
  assign n632 = n232 | n171;
  assign n633 = n236 | n539;
  assign n634 = n342 | n233;
  assign n635 = n672 & (n252 | ~n332 | n529);
  assign n636 = n546 | n454;
  assign n637 = n232 | n159;
  assign n638 = n182 | n416;
  assign n639 = n430 | n557;
  assign n640 = n422 | n540;
  assign n641 = i_2_ | n530;
  assign n642 = n402 & n623 & n641 & n394;
  assign n643 = n425 | n237;
  assign n644 = n237 | n208;
  assign n645 = n415 | n564;
  assign n646 = n415 | n576;
  assign n647 = n138 & n263 & n694 & n610 & n501 & n677 & n297;
  assign n648 = n440 | n576;
  assign n649 = n440 | n303;
  assign n650 = n59 & n57 & n648 & n649 & n587;
  assign n651 = n339 | n591;
  assign n652 = i_5_ | n236 | n514;
  assign n653 = n528 | n422;
  assign n654 = n303 | n194;
  assign n655 = n742 & n55 & n180;
  assign n656 = n181 | n454;
  assign n657 = n236 | n448;
  assign n658 = n198 | n182;
  assign n659 = n214 & n235 & n671 & n58 & n652 & n137;
  assign n660 = n528 | n425;
  assign n661 = n440 | n572;
  assign n662 = n725 & n632 & n581 & n231 & n400 & n699 & n584;
  assign n663 = n147 & n143 & n644 & n410 & n296 & n201 & n362 & n743;
  assign n664 = n651 & n445 & n628;
  assign n665 = n670 & n713 & n668 & n633 & n598 & n600;
  assign n666 = n180 & n257 & n151 & n49 & n694 & n742;
  assign n667 = n403 & n219 & n555 & n392 & n371 & n629;
  assign n668 = n415 | n448;
  assign n669 = n208 | n549;
  assign n670 = n454 | n441;
  assign n671 = n440 | n467;
  assign n672 = n440 | n195;
  assign n673 = n422 | n209;
  assign n674 = n236 | n453;
  assign n675 = n198 | n425;
  assign n676 = n236 | n493;
  assign n677 = n440 | n538;
  assign n678 = n301 | n561 | n444;
  assign n679 = n208 | n303;
  assign n680 = n263 & n610 & n56;
  assign n681 = n208 | n467;
  assign n682 = n539 | n449;
  assign n683 = ~n461 | ~i_3_ | n454;
  assign n684 = n658 & n288 & n623 & n653 & n631 & n630 & n595;
  assign n685 = n301 | n423;
  assign n686 = n301 | n535;
  assign n687 = n536 | n229;
  assign n688 = n208 | n575;
  assign n689 = n422 | n531 | n356;
  assign n690 = n241 | n378;
  assign n691 = n301 | n241 | n472;
  assign n692 = n538 | n454;
  assign n693 = n314 | n544;
  assign n694 = n440 | n539;
  assign n695 = n190 | n548;
  assign n696 = n192 | n389;
  assign n697 = n208 | n448;
  assign n698 = n236 | n335;
  assign n699 = n342 | n590;
  assign n700 = n153 & (n440 | n223 | n306);
  assign n701 = n440 | n549;
  assign n702 = n305 | ~i_7_ | n244;
  assign n703 = n527 | n182 | n373;
  assign n704 = n638 & n235 & n136 & n677 & n669 & n567 & n217;
  assign n705 = n540 | n574;
  assign n706 = n425 | n241 | n547;
  assign n707 = n164 & (n321 | n415 | n543);
  assign n708 = n181 | n301;
  assign n709 = n674 & (~i_7_ | n223 | n248);
  assign n710 = n342 | n541;
  assign n711 = n158 | n337;
  assign n712 = ~i_3_ | i_5_ | n305 | n415;
  assign n713 = n422 | n198;
  assign n714 = n712 & (n354 | ~n461 | n529);
  assign n715 = n171 | n323;
  assign n716 = i_7_ | n244 | ~n461;
  assign n717 = n301 | n225 | n226;
  assign n718 = n717 & (n419 | n346);
  assign n719 = n182 | n453;
  assign n720 = n529 | n225 | n488;
  assign n721 = n679 & (n226 | n438);
  assign n722 = (n449 | n195) & (n223 | n224);
  assign n723 = (n527 | n194) & (n301 | n232);
  assign n724 = (n529 | n444) & (n190 | n166);
  assign n725 = n339 | n233;
  assign n726 = n549 | n194;
  assign n727 = n517 & n149 & n725 & n726;
  assign n728 = i_8_ | n252 | n488;
  assign n729 = n728 & (n240 | n373 | n415);
  assign n730 = n729 & (i_3_ | n454 | ~n461);
  assign n731 = n533 | n236 | ~n332;
  assign n732 = (n475 | n425) & (n473 | n241);
  assign n733 = (n194 | n512) & (n529 | n540);
  assign n734 = n733 & (n430 | (n724 & n723));
  assign n735 = ~i_0_ | ~i_2_ | ~i_7_ | n342;
  assign n736 = n280 & n89 & n735 & n380 & n169 & n83;
  assign n737 = (~n332 | n486) & (n232 | n591);
  assign n738 = n489 | n190;
  assign n739 = n373 | n208 | n547;
  assign n740 = (n533 | n415) & (n422 | n232);
  assign n741 = n383 & n295 & n675;
  assign n742 = i_4_ | i_6_ | n514;
  assign n743 = n215 & n204 & n690 & n162 & n726 & n258;
  assign n744 = n184 & (n534 | n236);
  assign n745 = ~i_2_ | ~i_5_ | n748 | n749;
  assign n746 = i_3_ | n430 | n574;
  assign n747 = n487 | n565;
  assign n748 = i_1_ & (i_4_ | n229);
  assign n749 = ~i_1_ & (~i_4_ | n208);
endmodule


