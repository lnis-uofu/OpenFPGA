`ifndef STIMULI_IF
`define STIMULI_IF

//`timescale 1ns / 1ps
// Not using this interface, instead connecting directly to bs_if
interface stimuli_if();

// insert signals

endinterface


`endif
