// Benchmark "TOP" written by ABC on Tue Mar  5 09:56:39 2019

module diffeq ( clk, 
    PRESET, Pdxport_0_0_, Pdxport_1_1_, Pdxport_2_2_, Pdxport_3_3_,
    Pdxport_4_4_, Pdxport_5_5_, Pdxport_6_6_, Pdxport_7_7_, Pdxport_8_8_,
    Pdxport_9_9_, Pdxport_10_10_, Pdxport_11_11_, Paport_0_0_, Paport_1_1_,
    Paport_2_2_, Paport_3_3_, Paport_4_4_, Paport_5_5_, Paport_6_6_,
    Paport_7_7_, Paport_8_8_, Paport_9_9_, Paport_10_10_, Paport_11_11_,
    Preset_0_0_, Pready_0_0_,
    PDN, Pnext_0_0_, Pover_0_0_  );
  input  clk, PRESET, Pdxport_0_0_, Pdxport_1_1_, Pdxport_2_2_,
    Pdxport_3_3_, Pdxport_4_4_, Pdxport_5_5_, Pdxport_6_6_, Pdxport_7_7_,
    Pdxport_8_8_, Pdxport_9_9_, Pdxport_10_10_, Pdxport_11_11_,
    Paport_0_0_, Paport_1_1_, Paport_2_2_, Paport_3_3_, Paport_4_4_,
    Paport_5_5_, Paport_6_6_, Paport_7_7_, Paport_8_8_, Paport_9_9_,
    Paport_10_10_, Paport_11_11_, Preset_0_0_, Pready_0_0_;
  output PDN, Pnext_0_0_, Pover_0_0_;
  reg N_N4054, N_N3745, N_N4119, N_N3826, N_N3818, N_N3345, N_N3924,
    N_N3815, N_N3691, N_N3157, N_N3872, N_N3788, N_N3375, N_N3143, N_N4197,
    N_N3843, N_N3426, N_N4118, N_N3580, N_N3175, N_N3071, N_N3808, N_N3923,
    N_N3250, N_N4221, N_N3069, N_N3464, N_N3535, N_N3871, N_N3248, N_N4180,
    N_N3311, N_N3442, N_N3981, N_N3842, N_N3105, N_N4133, N_N4117, N_N3420,
    N_N3761, N_N3062, N_N4071, N_N4227, N_N3807, N_N4145, N_N3922, N_N3516,
    N_N3489, N_N4030, N_N3540, N_N3513, N_N4083, N_N3841, N_N4018, N_N3971,
    N_N4232, N_N4246, N_N3806, N_N3992, N_N4086, N_N4230, N_N4212,
    Pnext_0_0_, N_N3626, N_N3965, N_N3890, NDN3_11, NDN5_10, N_N3786,
    N_N4171, NDN5_16, N_N3799, N_N3844, N_N3196, N_N4126, N_N3681, N_N3679,
    N_N3340, N_N4116, N_N3810, N_N3235, N_N3283, N_N3716, N_N3701, N_N3921,
    N_N3625, N_N3751, N_N3736, N_N3870, N_N4024, N_N3876, N_N3840, N_N4021,
    N_N3932, NLC1_2, N_N3805, N_N3700, N_N3735, NLak3_2, NLak3_9, N_N3906,
    N_N3388, N_N4057, N_N3011, N_N3346, N_N3677, N_N4165, N_N4080, N_N3373,
    N_N3709, N_N4206, N_N3324, N_N3575, N_N4159, NAK5_2, N_N3916, N_N3743,
    N_N4242, N_N3312, N_N3733, N_N3774, N_N4214, N_N3294, N_N3796, N_N3574,
    N_N3791, N_N3480, N_N4243, N_N3940, N_N3509, N_N4015, N_N2989, N_N3919,
    N_N3578, N_N3529, N_N4222, N_N3910, N_N3868, N_N3947, N_N4181, N_N3793,
    N_N3822, N_N3813, N_N4114, N_N4134, N_N3866, N_N4218, N_N3939, N_N3776,
    N_N3387, N_N4194, N_N3821, N_N3882, N_N4167, N_N3800, N_N4237, N_N3417,
    N_N3918, N_N4158, N_N3630, N_N3344, N_N4072, N_N3274, N_N3473, N_N4205,
    N_N4111, N_N3680, N_N3838, N_N3262, N_N4099, N_N3607, N_N3323, N_N3612,
    N_N4079, PDN, N_N3457, N_N3445, N_N3794, N_N3663, N_N3715, N_N4039,
    N_N3280, N_N4239, N_N3988, N_N3433, N_N4075, N_N3468, N_N4045, N_N3482,
    N_N3832, N_N3304, N_N3750, N_N3634, N_N3293, N_N3659, N_N4252, N_N3912,
    N_N3862, N_N3221, N_N3875, N_N3949, N_N3908, N_N3711, N_N3931, N_N3469,
    N_N3436, N_N3974, N_N3905, N_N3741, N_N3369, N_N3164, N_N3500, N_N3996,
    N_N3356, N_N4093, Pover_0_0_, N_N4224, N_N4027, NDN1_4, N_N3384,
    N_N4036, N_N3968, N_N4183, NGFDN_3, N_N4090, N_N4004, N_N3205, N_N4136,
    N_N3303, N_N3533, N_N3336, N_N3961, N_N3331, N_N3203, N_N4236, N_N3884,
    N_N3367, N_N4140, NDN2_2, N_N4106, N_N3100, N_N4193, N_N3470, N_N3424,
    N_N3959, N_N3393, N_N4042, N_N3188, N_N4095, N_N3957, N_N3517, N_N4047,
    N_N3081, N_N3541, N_N4177, NDN3_3, N_N4176, N_N3585, NDN3_8, N_N4209,
    N_N3824, N_N4208, N_N4120, N_N3708, N_N4220, N_N3999, N_N4223, N_N3179,
    N_N4179, N_N3475, N_N4132, N_N4182, N_N3797, N_N3214, N_N4070, N_N4135,
    NLD3_9, NDN5_2, NDN5_3, N_N3778, NDN5_4, N_N3212, NDN5_5, NDN5_6,
    NDN5_7, NDN5_8, N_N4073, NDN5_9, NEN5_9, N_N3684, N_N4056, N_N3713,
    N_N3829, N_N4060, NSr3_2, NSr5_2, NSr5_3, N_N3462, N_N3460, NSr5_4,
    NSr3_9, NSr5_5, NSr5_7, NSr5_8, N_N3998;
  wire n946, n947, n949, n951, n953, n955, n957, n959, n961, n963, n965,
    n967, n969, n971, n973, n975, n977, n979, n981, n983, n985, n987, n989,
    n991, n993, n995, n997, n999, n1001, n1003, n1005, n1007, n1009,
    n1011_1, n1013, n1015, n1017, n1019, n1021_1, n1023, n1025, n1027,
    n1030, n1032, n1034, n1036_1, n1038, n1040, n1042, n1044, n1046_1,
    n1048, n1050, n1052, n1054, n1056_1, n1058, n1060, n1062, n1065, n1067,
    n1069, n1071_1, n1073, n1076_1, n1078, n1081, n1083, n1085, n1087,
    n1089, n1091, n1093, n1095, n1097, n1099, n1101_1, n1104, n1106_1,
    n1107, n1110, n1112, n1114, n1116, n1118, n1120, n1122, n1124, n1126_1,
    n1128, n1130, n1132, n1134, n1136_1, n1138, n1140_1, n1142, n1145_1,
    n1147, n1149, n1151, n1153, n1155_1, n1157, n1159, n1161, n1163,
    n1165_1, n1167, n1169, n1171, n1173, n1176, n1178, n1180, n1182, n1184,
    n1186, n1189, n1192, n1194, n1196, n1198, n1200, n1202, n1204, n1206,
    n1211, n1213, n1215_1, n1217, n1220_1, n1223, n1225_1, n1227, n1229,
    n1231, n1233, n1235, n1237, n1239, n1241, n1244, n1248, n1250, n1252,
    n1254, n1256, n1258, n1260_1, n1262, n1264, n1266, n1268, n1270_1,
    n1272, n1274, n1276, n1278, n1280_1, n1282, n1284, n1286, n1288, n1291,
    n1293, n1295, n1297, n1299, n1301, n1303, n1305_1, n1307, n1309, n1311,
    n1313, n1315_1, n1317, n1319, n1321, n1323, n1325_1, n1330_1, n1332,
    n1334, n1336, n1338, n1340_1, n1342, n1344, n1346, n1348, n1350_1,
    n1352, n1355_1, n1357, n1359, n1361, n1363, n1365_1, n1367, n1369,
    n1371, n1373, n1375_1, n1377, n1380_1, n1382, n1384, n1387, n1389,
    n1391, n1393, n1395_1, n1397, n1399, n1401, n1404, n1407, n1409, n1411,
    n1413, n1416, n1418, n1420_1, n1422, n1424, n1426, n1428, n1430_1,
    n1432, n1434, n1437, n1439, n1441, n1443, n1445_1, n1447, n1449, n1451,
    n1453, n1455_1, n1457, n1459, n1461, n1463, n1465_1, n1469, n1471,
    n1473, n1475_1, n1479, n1481, n1483, n1485_1, n1487, n1489, n1491,
    n1493, n1495_1, n1497, n1499, n1501, n1503, n1505_1, n1507, n1509,
    n1510_1, n1511, n1512, n1513, n1514, n1515_1, n1516, n1517, n1518,
    n1519, n1520_1, n1521, n1522, n1523, n1524, n1525_1, n1526, n1527,
    n1528, n1529, n1530_1, n1531, n1532, n1533, n1534, n1535_1, n1536,
    n1537, n1538, n1539, n1540_1, n1541, n1542, n1543, n1544, n1545_1,
    n1546, n1547, n1548, n1549, n1550_1, n1551, n1552, n1553, n1554,
    n1555_1, n1556, n1557, n1558, n1559, n1560_1, n1561, n1562, n1564,
    n1565_1, n1566, n1567, n1568, n1569, n1570_1, n1571, n1572, n1573,
    n1574, n1575_1, n1576, n1577, n1578, n1579, n1580_1, n1581, n1582,
    n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
    n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
    n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
    n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
    n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
    n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
    n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
    n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
    n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
    n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
    n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
    n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
    n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
    n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
    n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
    n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
    n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
    n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
    n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
    n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
    n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
    n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
    n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
    n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
    n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
    n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
    n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
    n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
    n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
    n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
    n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
    n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
    n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
    n1913, n1914, n1915, n1916, n1918, n1920, n1923, n1924, n1925, n1926,
    n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
    n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
    n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
    n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
    n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1975, n1976, n1979,
    n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
    n1990, n1991, n1992, n1993, n63_1, n68_1, n73_1, n78_1, n83_1, n88,
    n93_1, n98_1, n103, n108_1, n113_1, n118_1, n123_1, n128, n133, n138_1,
    n143_1, n148_1, n153_1, n158_1, n163_1, n168_1, n173_1, n178_1, n183_1,
    n188_1, n193_1, n198_1, n203_1, n208_1, n213_1, n218_1, n223_1, n228_1,
    n233, n238, n243_1, n248_1, n253_1, n258_1, n263_1, n268, n273, n278_1,
    n283, n288_1, n293, n298, n303_1, n308_1, n313_1, n318_1, n323_1,
    n328_1, n333_1, n338_1, n343_1, n348_1, n353_1, n358_1, n363_1, n368,
    n373, n377, n382_1, n387_1, n392_1, n397_1, n402_1, n407, n412_1,
    n417_1, n422_1, n427, n432_1, n437_1, n442, n447, n452_1, n457, n462,
    n467, n472, n477, n482, n487_1, n492, n497, n502_1, n507, n512, n517_1,
    n522_1, n527, n532, n537_1, n542_1, n547, n552, n557_1, n562, n567_1,
    n572, n577_1, n582, n587, n592, n597_1, n602_1, n607_1, n612, n617,
    n622, n627, n632, n637_1, n642_1, n647, n652, n657, n662_1, n667, n672,
    n677, n682_1, n687_1, n692, n697, n702_1, n707, n712_1, n717, n722_1,
    n727_1, n732, n737, n742_1, n747, n752_1, n757, n762, n767_1, n772,
    n777, n782, n787, n792, n797, n802_1, n807_1, n812_1, n817, n822_1,
    n827_1, n832_1, n837, n842_1, n847_1, n852_1, n857_1, n862, n867_1,
    n872_1, n877, n882_1, n887_1, n892_1, n897_1, n902, n907, n912, n917,
    n922, n927_1, n932_1, n936, n941, n946_1, n951_1, n956_1, n961_1,
    n966_1, n971_1, n976, n981_1, n986, n991_1, n996, n1001_1, n1006_1,
    n1011, n1016_1, n1021, n1026, n1031_1, n1036, n1041_1, n1046, n1051_1,
    n1056, n1061_1, n1066_1, n1071, n1076, n1081_1, n1086_1, n1091_1,
    n1096, n1101, n1106, n1111, n1116_1, n1121, n1126, n1131, n1136, n1140,
    n1145, n1150, n1155, n1160, n1165, n1170, n1175, n1180_1, n1185_1,
    n1190, n1195_1, n1200_1, n1205_1, n1210_1, n1215, n1220, n1225,
    n1230_1, n1235_1, n1240, n1245_1, n1250_1, n1255, n1260, n1265, n1270,
    n1275_1, n1280, n1285_1, n1290_1, n1295_1, n1300, n1305, n1310, n1315,
    n1320, n1325, n1330, n1335, n1340, n1345, n1350, n1355, n1360, n1365,
    n1370, n1375, n1380, n1385, n1390, n1395, n1400, n1405, n1410, n1415,
    n1420, n1425, n1430, n1435, n1440, n1445, n1450, n1455, n1460, n1465,
    n1470, n1475, n1480, n1485, n1490, n1495, n1500, n1505, n1510, n1515,
    n1520, n1525, n1530, n1535, n1540, n1545, n1550, n1555, n1560, n1565,
    n1570, n1575, n1580;
  assign n946 = ~PRESET & n1558;
  assign n947 = N_N3460 & ~n1556 & n1557;
  assign n1385 = n946 & (n947 | N_N3999);
  assign n949 = (n1585 | ~N_N4239) & (PRESET | n1584);
  assign n971_1 = ~n949;
  assign n951 = n1586 | ~N_N4232;
  assign n338_1 = ~n951;
  assign n953 = n1586 | ~N_N4230;
  assign n363_1 = ~n953;
  assign n955 = n1586 | ~N_N4218;
  assign n792 = ~n955;
  assign n957 = ~PRESET & n1961;
  assign n737 = N_N4222 & n957;
  assign n959 = (n1644 | ~n1934) & (~n1962 | ~N_N4167);
  assign n827_1 = ~n959;
  assign n961 = (n1585 | ~N_N4140) & (PRESET | n1646);
  assign n1245_1 = ~n961;
  assign n963 = (n1648 | ~n1934) & (n1647 | ~N_N4114);
  assign n777 = ~n963;
  assign n965 = (n1653 | n1654) & (n1652 | ~N_N4111);
  assign n887_1 = ~n965;
  assign n967 = n1586 | ~N_N4106;
  assign n1255 = ~n967;
  assign n969 = (n1585 | ~N_N4099) & (PRESET | n1656);
  assign n907 = ~n969;
  assign n971 = (n1585 | ~N_N4095) & (PRESET | n1658);
  assign n1300 = ~n971;
  assign n973 = n1586 | ~N_N4090;
  assign n1180_1 = ~n973;
  assign n975 = (n1585 | ~N_N4086) & (PRESET | n1660);
  assign n358_1 = ~n975;
  assign n977 = (n1662 | n1663) & (n1661 | ~N_N4075);
  assign n986 = ~n977;
  assign n979 = (n1586 | ~N_N4056) & (~Paport_5_5_ | n1587);
  assign n1510 = ~n979;
  assign n981 = (n1586 | ~N_N4054) & (~Paport_7_7_ | n1587);
  assign n63_1 = ~n981;
  assign n983 = (n1665 | n1666) & (n1664 | ~N_N4047);
  assign n1315 = ~n983;
  assign n985 = (n1664 | ~N_N4045) & (n1663 | n1665);
  assign n996 = ~n985;
  assign n987 = (n1668 | n1669) & (n1667 | ~N_N4042);
  assign n1290_1 = ~n987;
  assign n989 = (n1668 | n1670) & (n1667 | ~N_N4039);
  assign n961_1 = ~n989;
  assign n991 = (n1648 | n1709) & (n1647 | ~N_N4079);
  assign n927_1 = ~n991;
  assign n993 = (n1711 | n1712) & (n1710 | ~N_N4030);
  assign n303_1 = ~n993;
  assign n995 = (n1713 | ~N_N4236) & (n1670 | n1714);
  assign n1230_1 = ~n995;
  assign n997 = (n1662 | n1715) & (n1661 | ~N_N4024);
  assign n507 = ~n997;
  assign n999 = (n1662 | n1716) & (n1661 | ~N_N4021);
  assign n522_1 = ~n999;
  assign n1001 = (n1586 | ~N_N4057) & (~Pdxport_2_2_ | n1587);
  assign n572 = ~n1001;
  assign n1003 = (n1738 | n1739) & (n1737 | ~N_N3988);
  assign n976 = ~n1003;
  assign n1005 = (n1654 | n1740) & (n1652 | ~N_N3981);
  assign n228_1 = ~n1005;
  assign n1007 = (n1665 | n1741) & (n1664 | ~N_N4116);
  assign n452_1 = ~n1007;
  assign n1009 = (n1668 | n1741) & (n1667 | ~N_N3968);
  assign n1165 = ~n1009;
  assign n1011_1 = (n1586 | ~N_N4179) & (~Pdxport_5_5_ | n1587);
  assign n1400 = ~n1011_1;
  assign n1013 = (n1662 | n1741) & (n1661 | ~N_N3959);
  assign n1280 = ~n1013;
  assign n1015 = (n1662 | n1742) & (n1661 | ~N_N3957);
  assign n1305 = ~n1015;
  assign n1017 = (n1644 | n1743) & (~n1962 | ~N_N3947);
  assign n752_1 = ~n1017;
  assign n1019 = (n1586 | ~N_N4220) & (~Pdxport_3_3_ | n1587);
  assign n1380 = ~n1019;
  assign n1021_1 = (n1586 | ~N_N3916) & (~Paport_0_0_ | n1587);
  assign n637_1 = ~n1021_1;
  assign n1023 = (n1586 | ~N_N4243) & (~Paport_6_6_ | n1587);
  assign n697 = ~n1023;
  assign n1025 = (n1586 | ~N_N4015) & (~Paport_8_8_ | n1587);
  assign n712_1 = ~n1025;
  assign n1027 = (n1714 | n1744) & (n1713 | ~N_N3910);
  assign n742_1 = ~n1027;
  assign n1096 = N_N3905 & n957;
  assign n1030 = (n1586 | ~N_N4120) & (~Pdxport_1_1_ | n1587);
  assign n1370 = ~n1030;
  assign n1032 = (n1808 | ~N_N4197) & (n1806 | n1807);
  assign n133 = ~n1032;
  assign n1034 = (n1644 | n1809) & (~n1962 | ~N_N3829);
  assign n1520 = ~n1034;
  assign n1036_1 = (n1644 | n1810) & (~n1962 | ~N_N3826);
  assign n78_1 = ~n1036_1;
  assign n1038 = (n1662 | n1669) & (n1661 | ~N_N3824);
  assign n1360 = ~n1038;
  assign n1040 = (n1586 | ~N_N3818) & (~Paport_9_9_ | n1587);
  assign n83_1 = ~n1040;
  assign n1042 = (n1644 | n1811) & (~n1962 | ~N_N3815);
  assign n98_1 = ~n1042;
  assign n1044 = n1586 | ~N_N3876;
  assign n512 = ~n1044;
  assign n1046_1 = (n1585 | ~N_N3971) & (PRESET | n1813);
  assign n333_1 = ~n1046_1;
  assign n1048 = (n1668 | n1715) & (n1667 | ~N_N3799);
  assign n417_1 = ~n1048;
  assign n1050 = (n1644 | n1814) & (~n1962 | ~N_N3796);
  assign n677 = ~n1050;
  assign n1052 = (n1644 | n1815) & (~n1962 | ~N_N3788);
  assign n118_1 = ~n1052;
  assign n1054 = n1586 | ~N_N3786;
  assign n402_1 = ~n1054;
  assign n1056_1 = (n1665 | n1712) & (n1664 | ~N_N3870);
  assign n502_1 = ~n1056_1;
  assign n1058 = ~PRESET & ~NGFDN_3;
  assign n1350 = n1058 & (NDN3_8 | NDN3_3);
  assign n1060 = n1816 & (PRESET | ~N_N3745);
  assign n68_1 = ~n1060;
  assign n1062 = n1586 | ~N_N3741;
  assign n1101 = ~n1062;
  assign n1460 = ~PRESET & ~NSr5_4;
  assign n1065 = (n1808 | ~N_N3992) & (n1807 | n1817);
  assign n353_1 = ~n1065;
  assign n1067 = (n1713 | ~N_N4193) & (n1663 | n1714);
  assign n1265 = ~n1067;
  assign n1069 = (n1808 | ~N_N4018) & (n1807 | n1818);
  assign n328_1 = ~n1069;
  assign n1071_1 = (n1648 | n1819) & (n1647 | ~N_N3713);
  assign n1515 = ~n1071_1;
  assign n1073 = (n1711 | n1716) & (n1710 | ~N_N3711);
  assign n1071 = ~n1073;
  assign n1375 = N_N3708 & n957;
  assign n1076_1 = (n1586 | ~N_N3882) & (~Paport_10_10_ | n1587);
  assign n822_1 = ~n1076_1;
  assign n1078 = (n1714 | n1715) & (n1713 | ~N_N3793);
  assign n762 = ~n1078;
  assign n103 = N_N3691 & n957;
  assign n1081 = (n1644 | n1820) & (~n1962 | ~N_N3684);
  assign n1505 = ~n1081;
  assign n1083 = (n1585 | ~N_N4252) & (PRESET | n1822);
  assign n1036 = ~n1083;
  assign n1085 = (n1585 | ~N_N3843) & (PRESET | n1824);
  assign n138_1 = ~n1085;
  assign n1087 = (n1648 | n1825) & (n1647 | ~N_N3743);
  assign n642_1 = ~n1087;
  assign n1089 = (n1648 | n1826) & (n1647 | ~N_N3774);
  assign n662_1 = ~n1089;
  assign n1091 = (n1737 | ~N_N3663) & (n1670 | n1738);
  assign n951_1 = ~n1091;
  assign n1093 = (n1711 | n1741) & (n1710 | ~N_N4117);
  assign n248_1 = ~n1093;
  assign n1095 = (n1665 | n1670) & (n1664 | ~N_N3659);
  assign n1031_1 = ~n1095;
  assign n1097 = (n1648 | n1827) & (n1647 | ~N_N3791);
  assign n687_1 = ~n1097;
  assign n1099 = (n1711 | n1742) & (n1710 | ~N_N3922);
  assign n288_1 = ~n1099;
  assign n1101_1 = (n1654 | n1828) & (n1652 | ~N_N3761);
  assign n258_1 = ~n1101_1;
  assign n632 = ~PRESET & ~n1558;
  assign n1104 = n1586 | ~N_N3634;
  assign n1021 = ~n1104;
  assign n1106_1 = (n1735 | n1736) & (N_N3336 | ~N_N4205);
  assign n1107 = NLD3_9 & (n1106_1 | (N_N3336 & ~N_N4205));
  assign n532 = ~PRESET & ~PDN;
  assign n932_1 = n532 & (NGFDN_3 | ~n1169);
  assign n1110 = (n1829 | ~NEN5_9) & (NLD3_9 | n1830);
  assign n1500 = ~n1110;
  assign n1112 = (n1648 | n1831) & (n1647 | ~N_N3709);
  assign n607_1 = ~n1112;
  assign n1114 = (n1737 | ~N_N4071) & (n1669 | n1738);
  assign n268 = ~n1114;
  assign n1116 = (n1714 | n1716) & (n1713 | ~N_N3776);
  assign n802_1 = ~n1116;
  assign n1118 = (n1662 | n1670) & (n1661 | ~N_N3612);
  assign n922 = ~n1118;
  assign n1120 = (n1808 | ~N_N3949) & (n1807 | n1832);
  assign n1061_1 = ~n1120;
  assign n1122 = (n1836 | ~N_N4212) & (PRESET | n1835);
  assign n368 = ~n1122;
  assign n1124 = (n1836 | ~N_N4171) & (PRESET | n1838);
  assign n407 = ~n1124;
  assign n1126_1 = (n1586 | ~N_N3733) & (~Paport_2_2_ | n1587);
  assign n657 = ~n1126_1;
  assign n1128 = (n1585 | ~N_N3918) & (PRESET | n1840);
  assign n847_1 = ~n1128;
  assign n1130 = (n1585 | ~N_N3939) & (PRESET | n1842);
  assign n797 = ~n1130;
  assign n1132 = (n1585 | ~N_N4224) & (PRESET | n1844);
  assign n1140 = ~n1132;
  assign n1134 = (n1662 | n1845) & (n1661 | ~N_N3585);
  assign n1345 = ~n1134;
  assign n1136_1 = n1586 | ~N_N3580;
  assign n153_1 = ~n1136_1;
  assign n1138 = n1846 & (n1847 | ~N_N3751);
  assign n387_1 = ~n1138;
  assign n1140_1 = (n1654 | n1831) & (n1652 | ~N_N3794);
  assign n946_1 = ~n1140_1;
  assign n1142 = (n1662 | n1744) & (n1661 | ~N_N3625);
  assign n487_1 = ~n1142;
  assign n1335 = n1058 & (NDN3_3 | ~NSr3_2);
  assign n1145_1 = (n1665 | n1742) & (n1664 | ~N_N3921);
  assign n482 = ~n1145_1;
  assign n1147 = (n1586 | ~N_N3574) & (~Paport_4_4_ | n1587);
  assign n682_1 = ~n1147;
  assign n1149 = (n1586 | ~N_N4205) & (~Paport_11_11_ | n1587);
  assign n882_1 = ~n1149;
  assign n1151 = (n1585 | ~N_N4118) & (PRESET | n1849);
  assign n148_1 = ~n1151;
  assign n1153 = (n1585 | ~N_N4209) & (PRESET | n1851);
  assign n1355 = ~n1153;
  assign n1155_1 = (n1585 | ~N_N3500) & (PRESET | n1853);
  assign n1116_1 = ~n1155_1;
  assign n1157 = (n1654 | n1854) & (n1652 | ~N_N3489);
  assign n298 = ~n1157;
  assign n1159 = (n1654 | n1819) & (n1652 | ~N_N3513);
  assign n313_1 = ~n1159;
  assign n1161 = (n1738 | n1742) & (n1737 | ~N_N4221);
  assign n183_1 = ~n1161;
  assign n1163 = (n1586 | ~N_N4206) & (~Pdxport_6_6_ | n1587);
  assign n612 = ~n1163;
  assign n1165_1 = (n1667 | ~N_N3482) & (n1663 | n1668);
  assign n1001_1 = ~n1165_1;
  assign n1167 = n1855 & (n1847 | ~N_N4080);
  assign n1340 = ~n1167;
  assign n1169 = ~Preset_0_0_ | PDN | NLC1_2;
  assign n1250_1 = ~PRESET & n1169 & NDN2_2;
  assign n1171 = (n1648 | n1740) & (n1647 | ~N_N3475);
  assign n1405 = ~n1171;
  assign n1173 = (n1737 | ~N_N3473) & (n1663 | n1738);
  assign n877 = ~n1173;
  assign n557_1 = ~PRESET & n1107;
  assign n1176 = ~n1440 & (n1829 | ~NEN5_9);
  assign n1495 = ~n1176;
  assign n1178 = (n1667 | ~N_N3736) & (n1666 | n1668);
  assign n497 = ~n1178;
  assign n1180 = (n1654 | n1856) & (n1652 | ~N_N3535);
  assign n198_1 = ~n1180;
  assign n1182 = (n1808 | ~N_N3912) & (n1807 | n1857);
  assign n1041_1 = ~n1182;
  assign n1184 = (n1648 | n1862) & (n1647 | ~N_N4158);
  assign n852_1 = ~n1184;
  assign n1186 = (n1711 | n1739) & (n1710 | ~N_N3436);
  assign n1086_1 = ~n1186;
  assign n897_1 = ~PRESET & (n947 | N_N3838);
  assign n1189 = (n1711 | n1845) & (n1710 | ~N_N3841);
  assign n323_1 = ~n1189;
  assign n143_1 = N_N3426 & n957;
  assign n1192 = (n1665 | n1716) & (n1664 | ~N_N3424);
  assign n1275_1 = ~n1192;
  assign n1194 = n1586 | ~N_N3417;
  assign n842_1 = ~n1194;
  assign n1196 = (n1585 | ~N_N3842) & (PRESET | n1864);
  assign n233 = ~n1196;
  assign n1198 = (n1585 | ~N_N3924) & (PRESET | n1866);
  assign n93_1 = ~n1198;
  assign n1200 = (n1585 | ~N_N4119) & (PRESET | n1868);
  assign n73_1 = ~n1200;
  assign n1202 = n1586 | ~N_N3517;
  assign n1310 = ~n1202;
  assign n1204 = n1586 | ~N_N3681;
  assign n437_1 = ~n1204;
  assign n1206 = n1586 | ~N_N3716;
  assign n472 = ~n1206;
  assign n757 = N_N4181 & n957;
  assign n727_1 = N_N3578 & n946;
  assign n123_1 = N_N3375 & n957;
  assign n1211 = n1586 | ~N_N3373;
  assign n602_1 = ~n1211;
  assign n1213 = (n1665 | n1715) & (n1664 | ~N_N3367);
  assign n1240 = ~n1213;
  assign n1215_1 = n1586 | ~N_N3533;
  assign n1205_1 = ~n1215_1;
  assign n1217 = (n1585 | ~N_N3808) & (PRESET | n1870);
  assign n168_1 = ~n1217;
  assign n1470 = ~PRESET & ~NSr5_5;
  assign n1220_1 = (n1836 | ~N_N3340) & (PRESET | n1873);
  assign n447 = ~n1220_1;
  assign n1490 = N_N4073 & n957;
  assign n1223 = (~N_N3336 | n1652) & (n1654 | n1862);
  assign n1210_1 = ~n1223;
  assign n1225_1 = (n1737 | ~N_N4180) & (n1712 | n1738);
  assign n213_1 = ~n1225_1;
  assign n1227 = ~PRESET & (n1955 | (~n1229 & N_N4214));
  assign n667 = n1227 & N_N3462;
  assign n1229 = n1581 & ~N_N4060 & n1577 & n1579 & ~n1803 & n1872 & n1907 & n1956;
  assign n622 = ~PRESET & n1229;
  assign n1231 = (n1654 | n1827) & (n1652 | ~N_N3908);
  assign n1066_1 = ~n1231;
  assign n1233 = (n1654 | n1709) & (n1652 | ~N_N3884);
  assign n1235_1 = ~n1233;
  assign n1235 = (n1737 | ~N_N3323) & (n1716 | n1738);
  assign n917 = ~n1235;
  assign n1237 = n1586 | ~N_N3393;
  assign n1285_1 = ~n1237;
  assign n1239 = n1874 & (n1847 | ~N_N3932);
  assign n457 = ~n1239;
  assign n1241 = n1875 & (n1847 | ~N_N3876);
  assign n422_1 = ~n1241;
  assign n1390 = N_N4223 & n957;
  assign n1244 = (n1713 | ~N_N3311) & (n1669 | n1714);
  assign n218_1 = ~n1244;
  assign n1150 = NDN1_4 & n532;
  assign n392_1 = NDN3_11 & n1058;
  assign n1248 = (n1586 | ~N_N3778) & (~Paport_3_3_ | n1587);
  assign n1455 = ~n1248;
  assign n1250 = n1876 & (n1577 | n1807);
  assign n432_1 = ~n1250;
  assign n1252 = n1877 & (n1573 | n1807);
  assign n343_1 = ~n1252;
  assign n1254 = (n1644 | n1878) & (~n1962 | ~N_N3274);
  assign n872_1 = ~n1254;
  assign n1256 = (n1644 | n1879) & (~n1962 | ~N_N3480);
  assign n692 = ~n1256;
  assign n1258 = (n1585 | ~N_N3940) & (PRESET | n1881);
  assign n702_1 = ~n1258;
  assign n1260_1 = (n1662 | n1739) & (n1661 | ~N_N3700);
  assign n542_1 = ~n1260_1;
  assign n1262 = n1586 | ~N_N3250;
  assign n178_1 = ~n1262;
  assign n1264 = n1586 | ~N_N3248;
  assign n208_1 = ~n1264;
  assign n1266 = (n1648 | n1743) & (n1647 | ~N_N3931);
  assign n1076 = ~n1266;
  assign n1268 = (n1644 | n1882) & (~n1962 | ~N_N3509);
  assign n707 = ~n1268;
  assign n1270_1 = (n1644 | n1883) & (~n1962 | ~N_N3529);
  assign n732 = ~n1270_1;
  assign n1272 = (n1829 | ~NDN5_10) & (NLD3_9 | n1884);
  assign n397_1 = ~n1272;
  assign n1274 = (n1585 | ~N_N3923) & (PRESET | n1886);
  assign n173_1 = ~n1274;
  assign n1276 = (n1808 | ~N_N4145) & (n1807 | n1887);
  assign n283 = ~n1276;
  assign n1278 = (n1648 | n1820) & (n1647 | ~N_N3464);
  assign n193_1 = ~n1278;
  assign n1280_1 = (n1648 | n1809) & (n1647 | ~N_N3442);
  assign n223_1 = ~n1280_1;
  assign n1282 = (n1648 | n1828) & (n1647 | ~N_N3214);
  assign n1425 = ~n1282;
  assign n1284 = (n1648 | n1854) & (n1647 | ~N_N3212);
  assign n1465 = ~n1284;
  assign n1286 = (n1711 | n1744) & (n1710 | ~N_N3304);
  assign n1011 = ~n1286;
  assign n1288 = (n1711 | n1715) & (n1710 | ~N_N3221);
  assign n1051_1 = ~n1288;
  assign n867_1 = N_N4072 & n957;
  assign n1291 = (n1668 | n1742) & (n1667 | ~N_N3205);
  assign n1190 = ~n1291;
  assign n1293 = (n1668 | n1712) & (n1667 | ~N_N3203);
  assign n1225 = ~n1293;
  assign n1295 = n1888 & (n1847 | ~N_N3634);
  assign n832_1 = ~n1295;
  assign n1297 = (n1808 | ~N_N3996) & (n1807 | n1889);
  assign n1121 = ~n1297;
  assign n1299 = (n1586 | ~N_N4132) & (~Pdxport_7_7_ | n1587);
  assign n1410 = ~n1299;
  assign n1301 = (n1586 | ~N_N4070) & (~Pdxport_9_9_ | n1587);
  assign n1430 = ~n1301;
  assign n1303 = (n1586 | ~N_N4237) & (~Pdxport_11_11_ | n1587);
  assign n837 = ~n1303;
  assign n1305_1 = n1890 & (n1847 | ~N_N3517);
  assign n1195_1 = ~n1305_1;
  assign n1307 = n1891 & (n1847 | ~N_N3393);
  assign n1170 = ~n1307;
  assign n1309 = n1586 | ~N_N3932;
  assign n527 = ~n1309;
  assign n1311 = (n1648 | n1856) & (n1647 | ~N_N3179);
  assign n1395 = ~n1311;
  assign n1313 = (n1737 | ~N_N3293) & (n1666 | n1738);
  assign n1026 = ~n1313;
  assign n1315_1 = (n1738 | n1741) & (n1737 | ~N_N3175);
  assign n158_1 = ~n1315_1;
  assign n1317 = (n1710 | ~N_N3806) & (n1669 | n1711);
  assign n348_1 = ~n1317;
  assign n1319 = (n1710 | ~N_N3433) & (n1670 | n1711);
  assign n981_1 = ~n1319;
  assign n1321 = (n1836 | ~N_N3369) & (PRESET | n1893);
  assign n1106 = ~n1321;
  assign n1323 = (n1586 | ~N_N3797) & (~Paport_1_1_ | n1587);
  assign n1420 = ~n1323;
  assign n1325_1 = (n1668 | n1744) & (n1667 | ~N_N3626);
  assign n377 = ~n1325_1;
  assign n1445 = ~PRESET & ~NSr5_2;
  assign n782 = N_N4134 & n957;
  assign n941 = N_N3445 & n957;
  assign n1330_1 = n1894 & (n1847 | ~N_N3280);
  assign n772 = ~n1330_1;
  assign n1332 = n1586 | ~N_N3196;
  assign n427 = ~n1332;
  assign n1334 = (n1836 | ~N_N4093) & (PRESET | n1896);
  assign n1131 = ~n1334;
  assign n1336 = (n1586 | ~N_N4165) & (~Pdxport_4_4_ | n1587);
  assign n592 = ~n1336;
  assign n1338 = (n1738 | n1744) & (n1737 | ~N_N3387);
  assign n807_1 = ~n1338;
  assign n1340_1 = (n1710 | ~N_N3164) & (n1666 | n1711);
  assign n1111 = ~n1340_1;
  assign n1342 = (n1714 | n1742) & (n1713 | ~N_N3143);
  assign n128 = ~n1342;
  assign n1344 = (n1665 | n1845) & (n1664 | ~N_N3840);
  assign n517_1 = ~n1344;
  assign n1346 = (n1665 | n1669) & (n1664 | ~N_N3805);
  assign n537_1 = ~n1346;
  assign n1348 = n1897 & (n1847 | ~N_N4159);
  assign n1365 = ~n1348;
  assign n1350_1 = n1898 & (n1847 | ~N_N3235);
  assign n278_1 = ~n1350_1;
  assign n1352 = (n1585 | ~N_N3872) & (PRESET | n1900);
  assign n113_1 = ~n1352;
  assign n617 = N_N3324 & n957;
  assign n1355_1 = (n1654 | n1826) & (n1652 | ~N_N3862);
  assign n1046 = ~n1355_1;
  assign n1357 = n1586 | ~N_N3751;
  assign n492 = ~n1357;
  assign n1359 = (n1648 | n1883) & (n1647 | ~N_N3875);
  assign n1056 = ~n1359;
  assign n1361 = (n1808 | ~N_N3965) & (n1807 | n1901);
  assign n382_1 = ~n1361;
  assign n1363 = n1586 | ~N_N3105;
  assign n238 = ~n1363;
  assign n1365_1 = (n1737 | ~N_N3344) & (n1715 | n1738);
  assign n862 = ~n1365_1;
  assign n1367 = (n1710 | ~N_N3457) & (n1663 | n1711);
  assign n936 = ~n1367;
  assign n1369 = (n1665 | n1744) & (n1664 | ~N_N3303);
  assign n1200_1 = ~n1369;
  assign n1371 = n1902 & (n1579 | n1807);
  assign n1160 = ~n1371;
  assign n1373 = n1903 & (n1581 | n1807);
  assign n1185_1 = ~n1373;
  assign n1375_1 = (n1585 | ~N_N4177) & (PRESET | n1905);
  assign n1330 = ~n1375_1;
  assign n1377 = (n1654 | n1825) & (n1652 | ~N_N3832);
  assign n1006_1 = ~n1377;
  assign n88 = N_N3345 & n957;
  assign n1380_1 = (n1665 | n1739) & (n1664 | ~N_N3188);
  assign n1295_1 = ~n1380_1;
  assign n1382 = (n1713 | ~N_N3071) & (n1712 | n1714);
  assign n163_1 = ~n1382;
  assign n1384 = (n1714 | n1845) & (n1713 | ~N_N3069);
  assign n188_1 = ~n1384;
  assign n412_1 = NDN5_16 & ~n1829;
  assign n1387 = n1586 | ~N_N4159;
  assign n627 = ~n1387;
  assign n1389 = n1586 | ~N_N3331;
  assign n1220 = ~n1389;
  assign n1391 = (n1836 | ~N_N3283) & (PRESET | n1908);
  assign n467 = ~n1391;
  assign n1393 = (n1586 | ~N_N4242) & (~Pdxport_8_8_ | n1587);
  assign n647 = ~n1393;
  assign n1395_1 = (n1586 | ~N_N4194) & (~Pdxport_10_10_ | n1587);
  assign n812_1 = ~n1395_1;
  assign n1397 = (n1648 | n1815) & (n1647 | ~N_N3540);
  assign n308_1 = ~n1397;
  assign n1399 = (n1668 | n1716) & (n1667 | ~N_N3679);
  assign n442 = ~n1399;
  assign n1401 = (n1668 | n1739) & (n1667 | ~N_N3701);
  assign n477 = ~n1401;
  assign n1450 = ~PRESET & ~NSr5_3;
  assign n1404 = (n1648 | n1882) & (n1647 | ~N_N3750);
  assign n1016_1 = ~n1404;
  assign n991_1 = N_N3468 & n957;
  assign n1407 = n1816 & (PRESET | ~N_N3346);
  assign n582 = ~n1407;
  assign n1409 = n1909 & (n1847 | ~N_N3822);
  assign n1270 = ~n1409;
  assign n1411 = (n1668 | n1845) & (n1667 | ~N_N3100);
  assign n1260 = ~n1411;
  assign n1413 = (n1808 | ~N_N3974) & (n1807 | n1910);
  assign n1091_1 = ~n1413;
  assign n1475 = (NDN5_6 | ~n1514) & ~n1829;
  assign n1416 = (n1662 | n1666) & (n1661 | ~N_N3735);
  assign n547 = ~n1416;
  assign n1418 = (n1648 | n1878) & (n1647 | ~N_N3821);
  assign n817 = ~n1418;
  assign n1420_1 = n1586 | ~N_N4080;
  assign n597_1 = ~n1420_1;
  assign n1422 = n1586 | ~N_N3062;
  assign n263_1 = ~n1422;
  assign n1424 = (n1648 | n1814) & (n1647 | ~N_N3680);
  assign n892_1 = ~n1424;
  assign n1426 = (n1648 | n1879) & (n1647 | ~N_N3715);
  assign n956_1 = ~n1426;
  assign n1428 = n1586 | ~N_N3822;
  assign n767_1 = ~n1428;
  assign n1430_1 = (n1586 | ~N_N3906) & (~Pdxport_0_0_ | n1587);
  assign n562 = ~n1430_1;
  assign n1432 = (n1648 | n1653) & (n1647 | ~N_N3677);
  assign n587 = ~n1432;
  assign n1434 = (n1738 | n1845) & (n1737 | ~N_N4133);
  assign n243_1 = ~n1434;
  assign n1081_1 = N_N3469 & n957;
  assign n1437 = (n1648 | n1811) & (n1647 | ~N_N3516);
  assign n293 = ~n1437;
  assign n1439 = n1816 & (PRESET | ~N_N2989);
  assign n717 = ~n1439;
  assign n1441 = Pready_0_0_ & ~PDN & n1959 & ~NLak3_2;
  assign n552 = ~PRESET & NSr3_2 & n1441;
  assign n1443 = n1586 | ~N_N3262;
  assign n902 = ~n1443;
  assign n1445_1 = n1586 | ~N_N3280;
  assign n966_1 = ~n1445_1;
  assign n1447 = (n1808 | ~N_N4027) & (n1807 | n1911);
  assign n1145 = ~n1447;
  assign n1449 = n1586 | ~N_N3356;
  assign n1126 = ~n1449;
  assign n1451 = n1586 | ~N_N3384;
  assign n1155 = ~n1451;
  assign n1453 = (n1662 | n1712) & (n1661 | ~N_N3081);
  assign n1320 = ~n1453;
  assign n1455_1 = (n1714 | n1739) & (n1713 | ~N_N3630);
  assign n857_1 = ~n1455_1;
  assign n1457 = (n1713 | ~N_N3607) & (n1666 | n1714);
  assign n912 = ~n1457;
  assign n1459 = n1586 | ~N_N3235;
  assign n462 = ~n1459;
  assign n1461 = (n1648 | n1810) & (n1647 | ~N_N3420);
  assign n253_1 = ~n1461;
  assign n1463 = (n1714 | n1741) & (n1713 | ~N_N3157);
  assign n108_1 = ~n1463;
  assign n1465_1 = n1586 | ~N_N3011;
  assign n577_1 = ~n1465_1;
  assign n652 = N_N3312 & n957;
  assign n672 = N_N3294 & n957;
  assign n1469 = n1912 & (n1567 | n1807);
  assign n1215 = ~n1469;
  assign n1471 = (n1808 | ~N_N4083) & (n1807 | n1913);
  assign n318_1 = ~n1471;
  assign n1473 = n1586 | ~N_N3541;
  assign n1325 = ~n1473;
  assign n1475_1 = n1586 | ~N_N3866;
  assign n787 = ~n1475_1;
  assign n1415 = N_N4182 & n957;
  assign n1435 = N_N4135 & n957;
  assign n1479 = n1914 & (n1847 | ~N_N3262);
  assign n747 = ~n1479;
  assign n1481 = n1915 & (n1847 | ~N_N3417);
  assign n722_1 = ~n1481;
  assign n1483 = n1816 & (PRESET | ~N_N3388);
  assign n567_1 = ~n1483;
  assign n1485_1 = n1916 & (n1847 | ~N_N3786);
  assign n203_1 = ~n1485_1;
  assign n1487 = n532 & (~NSr3_2 | n1441);
  assign n1530 = ~n1487;
  assign n1489 = ~n1829 & ((~n1514 & NAK5_2) | ~NSr5_2);
  assign n1535 = ~n1489;
  assign n1491 = ~n1829 & (~NSr5_3 | (NAK5_2 & ~NSr5_2));
  assign n1540 = ~n1491;
  assign n1493 = n946 & (~N_N3462 | n1229);
  assign n1545 = ~n1493;
  assign n1495_1 = n946 & ~n1556 & (~N_N3462 | n1229);
  assign n1550 = ~n1495_1;
  assign n1497 = ~n1829 & (~NSr5_4 | (NAK5_2 & ~NSr5_3));
  assign n1555 = ~n1497;
  assign n1499 = n532 & (~NSr3_9 | (NDN3_8 & n1107));
  assign n1560 = ~n1499;
  assign n1501 = ~n1829 & ((~NSr5_4 & NAK5_2) | ~NSr5_5);
  assign n1565 = ~n1501;
  assign n1503 = ~n1829 & (~NSr5_7 | (NAK5_2 & ~NSr5_5));
  assign n1570 = ~n1503;
  assign n1505_1 = ~n1829 & (~NSr5_8 | (NAK5_2 & ~NSr5_7));
  assign n1575 = ~n1505_1;
  assign n1507 = ~PRESET & ~n1993 & (n1833 | ~N_N3998);
  assign n1580 = ~n1507;
  assign n1509 = ~n1958 & n1959;
  assign n1510_1 = ~NLD3_9 & n1583 & n1958;
  assign n1511 = ~PRESET & (n1509 | n1510_1);
  assign n1512 = n1559 & ~n1802;
  assign n1513 = ~PRESET & (n1512 | ~n1970);
  assign n1514 = NLak3_9 | ~NDN3_8 | ~NSr3_9;
  assign n1515_1 = (n1514 | ~NSr5_2) & (NSr5_4 | ~NSr5_5);
  assign n1516 = (n1528 | ~N_N3303) & (n1515_1 | ~N_N3906);
  assign n1517 = (n1542 | ~N_N3940) & (n1538 | ~N_N3939);
  assign n1518 = ~NSr5_7 | NSr5_5;
  assign n1519 = n1516 & n1517 & (n1518 | ~N_N3304);
  assign n1520_1 = (n1528 | ~N_N3188) & (n1515_1 | ~N_N4206);
  assign n1521 = (n1542 | ~N_N3813) & (n1538 | ~N_N4239);
  assign n1522 = n1520_1 & n1521 & (n1518 | ~N_N3436);
  assign n1523 = (n1528 | ~N_N3424) & (n1515_1 | ~N_N4165);
  assign n1524 = (n1542 | ~N_N3868) & (n1538 | ~N_N4099);
  assign n1525_1 = n1523 & n1524 & (n1518 | ~N_N3711);
  assign n1526 = (n1518 | ~N_N3221) & (n1515_1 | ~N_N4057);
  assign n1527 = (n1542 | ~N_N3919) & (n1538 | ~N_N3918);
  assign n1528 = NSr5_7 | ~NSr5_8;
  assign n1529 = n1526 & n1527 & (n1528 | ~N_N3367);
  assign n1530_1 = (n1528 | ~N_N4116) & (n1515_1 | ~N_N4120);
  assign n1531 = (n1542 | ~N_N4119) & (n1538 | ~N_N4118);
  assign n1532 = n1530_1 & n1531 & (n1518 | ~N_N4117);
  assign n1533 = (n1528 | ~N_N3921) & (n1515_1 | ~N_N4220);
  assign n1534 = (n1542 | ~N_N3924) & (n1538 | ~N_N3923);
  assign n1535_1 = n1533 & n1534 & (n1518 | ~N_N3922);
  assign n1536 = (n1528 | ~N_N3870) & (n1515_1 | ~N_N4179);
  assign n1537 = (n1542 | ~N_N3872) & (n1518 | ~N_N4030);
  assign n1538 = ~NSr5_4 | NSr5_3;
  assign n1539 = n1536 & n1537 & (n1538 | ~N_N3871);
  assign n1540_1 = (n1518 | ~N_N3164) & (n1515_1 | ~N_N4242);
  assign n1541 = (n1538 | ~N_N4252) & (n1528 | ~N_N4047);
  assign n1542 = ~NSr5_3 | NSr5_2;
  assign n1543 = n1540_1 & n1541 & (n1542 | ~N_N3800);
  assign n1544 = (n1528 | ~N_N3805) & (n1515_1 | ~N_N4070);
  assign n1545_1 = (n1542 | ~N_N3808) & (n1538 | ~N_N3807);
  assign n1546 = n1544 & n1545_1 & (n1518 | ~N_N3806);
  assign n1547 = (n1528 | ~N_N3840) & (n1515_1 | ~N_N4132);
  assign n1548 = (n1542 | ~N_N3843) & (n1538 | ~N_N3842);
  assign n1549 = n1547 & n1548 & (n1518 | ~N_N3841);
  assign n1550_1 = (n1518 | ~N_N3433) & (n1515_1 | ~N_N4237);
  assign n1551 = (n1542 | ~N_N4209) & (n1538 | ~N_N4208);
  assign n1552 = n1550_1 & n1551 & (n1528 | ~N_N3659);
  assign n1553 = (n1518 | ~N_N3457) & (n1515_1 | ~N_N4194);
  assign n1554 = (n1542 | ~N_N4177) & (n1538 | ~N_N4176);
  assign n1555_1 = n1553 & n1554 & (n1528 | ~N_N4045);
  assign n1556 = n1515_1 & n1528 & n1518 & n1542 & n1538;
  assign n1557 = (~N_N3999 | N_N3838) & ~n1992;
  assign n1558 = N_N3460 & (n1556 | n1557);
  assign n1559 = N_N3578 | n1558;
  assign n1560_1 = ~n1955 & (n1557 | n1559);
  assign n1561 = (~n1513 & (~N_N4060 | n1807)) | (N_N4060 & n1807);
  assign n1562 = PRESET | n1560_1;
  assign n1525 = n1561 & (n1519 | n1562);
  assign n1564 = N_N3369 | n1572;
  assign n1565_1 = n1564 & (~n1572 | ~N_N3369);
  assign n1566 = ~N_N4060 | N_N3961;
  assign n1567 = n1566 & (N_N4060 | ~N_N3961);
  assign n1568 = N_N4093 | n1570_1;
  assign n1569 = n1568 & (~n1570_1 | ~N_N4093);
  assign n1570_1 = N_N4212 | n1578;
  assign n1571 = n1570_1 & (~n1578 | ~N_N4212);
  assign n1572 = N_N4246 | n1568;
  assign n1573 = n1572 & (~n1568 | ~N_N4246);
  assign n1574 = N_N4171 | n1580_1;
  assign n1575_1 = n1574 & (~n1580_1 | ~N_N4171);
  assign n1576 = N_N4126 | n1566;
  assign n1577 = n1576 & (~n1566 | ~N_N4126);
  assign n1578 = N_N4036 | n1574;
  assign n1579 = n1578 & (~n1574 | ~N_N4036);
  assign n1580_1 = N_N4004 | n1576;
  assign n1581 = n1580_1 & (~n1576 | ~N_N4004);
  assign n1582 = (~n1509 | ~N_N4239) & (~NLD3_9 | ~N_N3774);
  assign n1583 = NDN3_8 | ~NDN3_3;
  assign n1584 = n1582 & (n1583 | ~N_N4090);
  assign n1585 = PRESET | ~n1510_1;
  assign n1586 = n1960 | PRESET;
  assign n1587 = PRESET | ~n1960;
  assign n1588 = NDN5_9 | ~NEN5_9;
  assign n1589 = NDN5_10 | NSr5_7;
  assign n1590 = (n1589 | ~N_N4039) & (n1588 | ~N_N3612);
  assign n1591 = (n1589 | ~N_N3482) & (n1588 | ~N_N4075);
  assign n1592 = (n1589 | ~N_N3736) & (n1588 | ~N_N3735);
  assign n1593 = (n1589 | ~N_N3701) & (n1588 | ~N_N3700);
  assign n1594 = (n1589 | ~N_N3679) & (n1588 | ~N_N4021);
  assign n1595 = (n1589 | ~N_N3626) & (n1588 | ~N_N3625);
  assign n1596 = (n1589 | ~N_N3799) & (n1588 | ~N_N4024);
  assign n1597 = (n1589 | ~N_N3968) & (n1588 | ~N_N3959);
  assign n1598 = (n1589 | ~N_N3205) & (n1588 | ~N_N3957);
  assign n1599 = (n1589 | ~N_N3203) & (n1588 | ~N_N3081);
  assign n1600 = (n1589 | ~N_N3100) & (n1588 | ~N_N3585);
  assign n1601 = (n1589 | ~N_N4042) & (n1588 | ~N_N3824);
  assign n1602 = (n1589 | ~N_N3470) & (n1588 | ~N_N3274);
  assign n1603 = (n1589 | ~N_N3810) & (n1588 | ~N_N3947);
  assign n1604 = n1627 & n1599 & n1593;
  assign n1605 = n1604 & n1600;
  assign n1606 = (n1589 | ~N_N4224) & (n1588 | ~N_N3829);
  assign n1607 = (n1589 | ~N_N3971) & (n1588 | ~N_N3796);
  assign n1608 = (n1589 | ~N_N3500) & (n1588 | ~N_N3684);
  assign n1609 = ~n1595 & ~n1607 & (~n1608 | ~n1610);
  assign n1610 = n1595 ^ ~n1597;
  assign n1611 = ~n1609 & (n1608 | n1610);
  assign n1612 = n1595 & n1597;
  assign n1613 = (n1589 | ~N_N4086) & (n1588 | ~N_N3480);
  assign n1614 = n1613 & ~n1924;
  assign n1615 = (n1613 | ~n1924) & (n1611 | n1614);
  assign n1616 = n1606 & n1615;
  assign n1617 = (n1616 | ~n1925) & (n1606 | n1615);
  assign n1618 = (n1589 | ~N_N3890) & (n1588 | ~N_N3509);
  assign n1619 = n1595 & n1597 & n1596;
  assign n1620 = n1619 & n1598;
  assign n1621 = n1618 & ~n1926;
  assign n1622 = (n1618 | ~n1926) & (n1617 | n1621);
  assign n1623 = (n1589 | ~N_N4183) & (n1588 | ~N_N3826);
  assign n1624 = n1623 & ~n1927;
  assign n1625 = (n1623 | ~n1927) & (n1622 | n1624);
  assign n1626 = (n1589 | ~N_N3844) & (n1588 | ~N_N3529);
  assign n1627 = n1619 & n1598 & n1594;
  assign n1628 = n1627 & n1599;
  assign n1629 = n1626 & ~n1928;
  assign n1630 = (n1626 | ~n1928) & (n1625 | n1629);
  assign n1631 = (n1589 | ~N_N4136) & (n1588 | ~N_N3815);
  assign n1632 = n1631 & ~n1929;
  assign n1633 = (n1631 | ~n1929) & (n1630 | n1632);
  assign n1634 = n1592 ^ ~n1605;
  assign n1635 = n1633 & n1634;
  assign n1636 = (n1603 | n1635) & (n1633 | n1634);
  assign n1637 = (n1589 | ~N_N4140) & (n1588 | ~N_N3788);
  assign n1638 = n1636 & n1637;
  assign n1639 = (n1638 | ~n1931) & (n1636 | n1637);
  assign n1640 = n1602 & n1639;
  assign n1641 = n1591 ^ ~n1963;
  assign n1642 = (n1640 | n1641) & (n1602 | n1639);
  assign n1643 = (n1589 | ~N_N4095) & (n1588 | ~N_N4167);
  assign n1644 = PRESET | n1589;
  assign n1645 = (~n1509 | ~N_N4140) & (~NLD3_9 | ~N_N3540);
  assign n1646 = n1645 & (n1583 | ~N_N3541);
  assign n1647 = PRESET | ~n1588;
  assign n1648 = PRESET | n1588;
  assign n1649 = NDN5_6 | n1514;
  assign n1650 = (n1649 | ~N_N3906) & (n1588 | ~N_N3910);
  assign n1651 = (n1649 | ~N_N3940) & (n1588 | ~N_N3939);
  assign n1652 = PRESET | ~n1649;
  assign n1653 = n1650 ^ ~n1651;
  assign n1654 = PRESET | n1649;
  assign n1655 = (n1583 | ~N_N3384) & (~n1509 | ~N_N4099);
  assign n1656 = n1655 & (~NLD3_9 | ~N_N3743);
  assign n1657 = (n1583 | ~N_N3866) & (~n1509 | ~N_N4095);
  assign n1658 = n1657 & (~NLD3_9 | ~N_N4114);
  assign n1659 = (~n1509 | ~N_N4086) & (~NLD3_9 | ~N_N3715);
  assign n1660 = n1659 & (n1583 | ~N_N3716);
  assign n1661 = PRESET | ~n1964;
  assign n1662 = PRESET | n1964;
  assign n1663 = ~n1557 | ~N_N4197;
  assign n1664 = PRESET | ~n1965;
  assign n1665 = PRESET | n1965;
  assign n1666 = ~n1557 | ~N_N4145;
  assign n1667 = PRESET | ~n1966;
  assign n1668 = PRESET | n1966;
  assign n1669 = ~n1557 | ~N_N3912;
  assign n1670 = ~n1557 | ~N_N4227;
  assign n1671 = (n1649 | ~N_N4194) & (n1588 | ~N_N4193);
  assign n1672 = (n1649 | ~N_N4177) & (n1588 | ~N_N4176);
  assign n1673 = (n1649 | ~N_N3800) & (n1588 | ~N_N4252);
  assign n1674 = (n1649 | ~N_N4242) & (n1588 | ~N_N3607);
  assign n1675 = (n1649 | ~N_N4220) & (n1588 | ~N_N3143);
  assign n1676 = (n1649 | ~N_N3924) & (n1588 | ~N_N3923);
  assign n1677 = (n1649 | ~N_N3919) & (n1588 | ~N_N3918);
  assign n1678 = (n1649 | ~N_N4057) & (n1588 | ~N_N3793);
  assign n1679 = (n1649 | ~N_N4119) & (n1588 | ~N_N4118);
  assign n1680 = (n1649 | ~N_N4120) & (n1588 | ~N_N3157);
  assign n1681 = ~n1650 & ~n1651 & (~n1679 | ~n1680);
  assign n1682 = ~n1681 & (n1679 | n1680);
  assign n1683 = n1678 & n1682;
  assign n1684 = (n1677 | n1683) & (n1678 | n1682);
  assign n1685 = n1676 & n1684;
  assign n1686 = (n1675 | n1685) & (n1676 | n1684);
  assign n1687 = (n1649 | ~N_N3868) & (n1588 | ~N_N4099);
  assign n1688 = (n1649 | ~N_N4165) & (n1588 | ~N_N3776);
  assign n1689 = n1687 & n1688;
  assign n1690 = (n1686 | n1689) & (n1687 | n1688);
  assign n1691 = (n1649 | ~N_N3872) & (n1588 | ~N_N3871);
  assign n1692 = (n1649 | ~N_N4179) & (n1588 | ~N_N3071);
  assign n1693 = n1691 & n1692;
  assign n1694 = (n1690 | n1693) & (n1691 | n1692);
  assign n1695 = (n1649 | ~N_N3813) & (n1588 | ~N_N4239);
  assign n1696 = (n1649 | ~N_N4206) & (n1588 | ~N_N3630);
  assign n1697 = n1695 & n1696;
  assign n1698 = (n1694 | n1697) & (n1695 | n1696);
  assign n1699 = (n1649 | ~N_N3843) & (n1588 | ~N_N3842);
  assign n1700 = (n1649 | ~N_N4132) & (n1588 | ~N_N3069);
  assign n1701 = n1699 & n1700;
  assign n1702 = (n1698 | n1701) & (n1699 | n1700);
  assign n1703 = n1674 & n1702;
  assign n1704 = (n1673 | n1703) & (n1674 | n1702);
  assign n1705 = (n1649 | ~N_N3808) & (n1588 | ~N_N3807);
  assign n1706 = (n1649 | ~N_N4070) & (n1588 | ~N_N3311);
  assign n1707 = n1705 & n1706;
  assign n1708 = (n1704 | n1707) & (n1705 | n1706);
  assign n1709 = n1708 ^ n1981;
  assign n1710 = PRESET | ~n1967;
  assign n1711 = PRESET | n1967;
  assign n1712 = ~n1557 | ~N_N3974;
  assign n1713 = PRESET | ~n1968;
  assign n1714 = PRESET | n1968;
  assign n1715 = ~n1557 | ~N_N3992;
  assign n1716 = ~n1557 | ~N_N4018;
  assign n1717 = N_N3916 & ~N_N4111 & (N_N3797 | ~N_N3535);
  assign n1718 = ~n1717 & (~N_N3797 | N_N3535);
  assign n1719 = n1718 & ~N_N3733;
  assign n1720 = (n1719 | N_N3794) & (n1718 | ~N_N3733);
  assign n1721 = n1720 & ~N_N3778;
  assign n1722 = (n1721 | N_N3981) & (n1720 | ~N_N3778);
  assign n1723 = ~n1722 & N_N3574;
  assign n1724 = (~n1722 | N_N3574) & (n1723 | ~N_N3832);
  assign n1725 = n1724 & ~N_N3761;
  assign n1726 = (n1725 | N_N4056) & (n1724 | ~N_N3761);
  assign n1727 = ~n1726 & N_N3862;
  assign n1728 = (~n1726 | N_N3862) & (n1727 | ~N_N4243);
  assign n1729 = n1728 & N_N3489;
  assign n1730 = (n1729 | ~N_N4054) & (n1728 | N_N3489);
  assign n1731 = ~n1730 & ~N_N3908;
  assign n1732 = (n1731 | N_N4015) & (~n1730 | ~N_N3908);
  assign n1733 = n1732 & ~N_N3513;
  assign n1734 = (n1733 | N_N3818) & (n1732 | ~N_N3513);
  assign n1735 = N_N3884 & (~n1734 | ~N_N3882);
  assign n1736 = ~n1734 & ~N_N3882;
  assign n1737 = PRESET | ~n1969;
  assign n1738 = PRESET | n1969;
  assign n1739 = ~n1557 | ~N_N4083;
  assign n1740 = n1684 ^ n1982;
  assign n1741 = ~n1557 | ~N_N4027;
  assign n1742 = ~n1557 | ~N_N3996;
  assign n1743 = n1634 ^ n1935;
  assign n1744 = ~n1557 | ~N_N3965;
  assign n1745 = (n1515_1 | ~N_N4095) & (~N_N3445 | n1538);
  assign n1746 = (n1528 | ~N_N4237) & (~N_N3905 | n1542);
  assign n1747 = n1745 & n1746 & (n1518 | ~N_N3663);
  assign n1748 = (n1515_1 | ~N_N3470) & (~N_N3468 | n1538);
  assign n1749 = (n1528 | ~N_N4194) & (n1518 | ~N_N3473);
  assign n1750 = n1748 & (~N_N3469 | n1542) & n1749;
  assign n1751 = (n1528 | ~N_N4070) & (n1515_1 | ~N_N4140);
  assign n1752 = (~N_N4072 | n1538) & (~N_N4073 | n1542);
  assign n1753 = n1751 & n1752 & (n1518 | ~N_N4071);
  assign n1754 = (n1518 | ~N_N3293) & (n1515_1 | ~N_N3810);
  assign n1755 = (n1528 | ~N_N4242) & (~N_N3426 | n1538);
  assign n1756 = n1754 & (~N_N3294 | n1542) & n1755;
  assign n1757 = (n1528 | ~N_N4132) & (n1515_1 | ~N_N4136);
  assign n1758 = (~N_N4134 | n1538) & (~N_N4135 | n1542);
  assign n1759 = n1757 & n1758 & (n1518 | ~N_N4133);
  assign n1760 = (n1515_1 | ~N_N3844) & (~N_N3312 | n1542);
  assign n1761 = (n1528 | ~N_N4206) & (n1518 | ~N_N3988);
  assign n1762 = n1760 & (~N_N3375 | n1538) & n1761;
  assign n1763 = (n1528 | ~N_N4179) & (n1515_1 | ~N_N4183);
  assign n1764 = (~N_N4181 | n1538) & (~N_N4182 | n1542);
  assign n1765 = n1763 & n1764 & (n1518 | ~N_N4180);
  assign n1766 = (n1518 | ~N_N3323) & (n1515_1 | ~N_N3890);
  assign n1767 = (n1528 | ~N_N4165) & (~N_N3691 | n1538);
  assign n1768 = n1766 & (~N_N3324 | n1542) & n1767;
  assign n1769 = (n1528 | ~N_N4220) & (n1515_1 | ~N_N4224);
  assign n1770 = (~N_N4222 | n1538) & (~N_N4223 | n1542);
  assign n1771 = n1769 & n1770 & (n1518 | ~N_N4221);
  assign n1772 = (n1518 | ~N_N3344) & (n1515_1 | ~N_N4086);
  assign n1773 = (n1542 | ~N_N3346) & (n1528 | ~N_N4057);
  assign n1774 = n1772 & (~N_N3345 | n1538) & n1773;
  assign n1775 = (n1538 | ~N_N2989) & (n1515_1 | ~N_N3500);
  assign n1776 = (n1528 | ~N_N4120) & (~N_N3708 | n1542);
  assign n1777 = n1775 & n1776 & (n1518 | ~N_N3175);
  assign n1778 = (n1518 | ~N_N3387) & (n1515_1 | ~N_N3971);
  assign n1779 = (n1538 | ~N_N3745) & (n1528 | ~N_N3906);
  assign n1780 = n1778 & n1779 & (n1542 | ~N_N3388);
  assign n1781 = n1780 | ~N_N3965;
  assign n1782 = n1777 & n1781;
  assign n1783 = (n1782 | ~N_N4027) & (n1777 | n1781);
  assign n1784 = n1783 & ~N_N3992;
  assign n1785 = (n1783 | ~N_N3992) & (n1774 | n1784);
  assign n1786 = n1785 & ~N_N3996;
  assign n1787 = (n1785 | ~N_N3996) & (n1771 | n1786);
  assign n1788 = n1787 & ~N_N4018;
  assign n1789 = (n1787 | ~N_N4018) & (n1768 | n1788);
  assign n1790 = n1789 & ~N_N3974;
  assign n1791 = (n1789 | ~N_N3974) & (n1765 | n1790);
  assign n1792 = n1791 & ~N_N4083;
  assign n1793 = (n1791 | ~N_N4083) & (n1762 | n1792);
  assign n1794 = n1793 & ~N_N3949;
  assign n1795 = (n1793 | ~N_N3949) & (n1759 | n1794);
  assign n1796 = n1795 & ~N_N4145;
  assign n1797 = (n1795 | ~N_N4145) & (n1756 | n1796);
  assign n1798 = n1797 & ~N_N3912;
  assign n1799 = (n1797 | ~N_N3912) & (n1753 | n1798);
  assign n1800 = n1799 & ~N_N4197;
  assign n1801 = (n1799 | ~N_N4197) & (n1750 | n1800);
  assign n1802 = ~n1803 | n1955;
  assign n1803 = ~N_N3462 | N_N3575 | ~N_N4214;
  assign n1804 = n1801 ^ n1747;
  assign n1805 = n1802 & (n1803 | n1804);
  assign n1806 = n1799 ^ n1936;
  assign n1807 = PRESET | n1803;
  assign n1808 = PRESET | n1802;
  assign n1809 = n1925 ^ ~n1937;
  assign n1810 = n1927 ^ ~n1938;
  assign n1811 = n1929 ^ ~n1939;
  assign n1812 = (~n1509 | ~N_N3971) & (~NLD3_9 | ~N_N3680);
  assign n1813 = n1812 & (n1583 | ~N_N3681);
  assign n1814 = n1595 ^ ~n1607;
  assign n1815 = n1931 ^ ~n1940;
  assign n1816 = PRESET | n1961;
  assign n1817 = n1783 ^ n1941;
  assign n1818 = n1787 ^ n1942;
  assign n1819 = n1706 ^ n1983;
  assign n1820 = n1610 ^ n1984;
  assign n1821 = (n1583 | ~N_N3533) & (~n1509 | ~N_N4252);
  assign n1822 = n1821 & (~NLD3_9 | ~N_N3791);
  assign n1823 = (n1583 | ~N_N3105) & (~n1509 | ~N_N3843);
  assign n1824 = n1823 & (~NLD3_9 | ~N_N3489);
  assign n1825 = n1688 ^ n1985;
  assign n1826 = n1696 ^ n1986;
  assign n1827 = n1702 ^ n1987;
  assign n1828 = n1692 ^ n1988;
  assign n1829 = PRESET | NLD3_9;
  assign n1830 = NSr5_8 | PRESET;
  assign n1831 = n1682 ^ n1989;
  assign n1832 = n1793 ^ n1943;
  assign n1833 = ~PDN & ~NLC1_2;
  assign n1834 = (n1522 | n1560_1) & (~N_N4212 | n1970);
  assign n1835 = n1834 & (n1571 | n1803);
  assign n1836 = PRESET | ~n1512;
  assign n1837 = (n1525_1 | n1560_1) & (~N_N4171 | n1970);
  assign n1838 = n1837 & (n1575_1 | n1803);
  assign n1839 = (n1583 | ~N_N3356) & (~n1509 | ~N_N3918);
  assign n1840 = n1839 & (~NLD3_9 | ~N_N3709);
  assign n1841 = (~n1509 | ~N_N3939) & (~NLD3_9 | ~N_N3677);
  assign n1842 = n1841 & (n1583 | ~N_N3741);
  assign n1843 = (~n1509 | ~N_N4224) & (~NLD3_9 | ~N_N3442);
  assign n1844 = n1843 & (n1583 | ~N_N4106);
  assign n1845 = ~n1557 | ~N_N3949;
  assign n1846 = (n1971 | ~N_N3750) & (~n1511 | ~N_N3890);
  assign n1847 = PRESET | n1583;
  assign n1848 = (~n1509 | ~N_N4118) & (~NLD3_9 | ~N_N3179);
  assign n1849 = n1848 & (n1583 | ~N_N4232);
  assign n1850 = (~NLD3_9 | ~N_N3336) & (~n1509 | ~N_N4209);
  assign n1851 = n1850 & (n1583 | ~N_N3373);
  assign n1852 = (n1583 | ~N_N3331) & (~n1509 | ~N_N3500);
  assign n1853 = n1852 & (~NLD3_9 | ~N_N3464);
  assign n1854 = n1700 ^ n1990;
  assign n1855 = (~n1511 | ~N_N4176) & (~N_N4079 | n1971);
  assign n1856 = n1944 ^ n1945;
  assign n1857 = n1797 ^ n1946;
  assign n1858 = (n1649 | ~N_N4237) & (n1588 | ~N_N4236);
  assign n1859 = (n1649 | ~N_N4209) & (n1588 | ~N_N4208);
  assign n1860 = n1708 & n1672;
  assign n1861 = (n1671 | n1860) & (n1672 | n1708);
  assign n1862 = n1861 ^ n1991;
  assign n1863 = (n1583 | ~N_N3196) & (~n1509 | ~N_N3842);
  assign n1864 = n1863 & (~NLD3_9 | ~N_N3212);
  assign n1865 = (n1583 | ~N_N3250) & (~n1509 | ~N_N3924);
  assign n1866 = n1865 & (~NLD3_9 | ~N_N3981);
  assign n1867 = (~NLD3_9 | ~N_N3535) & (~n1509 | ~N_N4119);
  assign n1868 = n1867 & (n1583 | ~N_N3580);
  assign n1869 = (n1583 | ~N_N3062) & (~n1509 | ~N_N3808);
  assign n1870 = n1869 & (~NLD3_9 | ~N_N3513);
  assign n1871 = (n1552 | n1560_1) & (~N_N3340 | n1970);
  assign n1872 = N_N3340 ^ n1923;
  assign n1873 = n1871 & (n1872 | n1803);
  assign n1874 = (~n1511 | ~N_N3810) & (~N_N3931 | n1971);
  assign n1875 = (~n1511 | ~N_N3844) & (~N_N3875 | n1971);
  assign n1876 = (n1529 | n1562) & (~n1513 | ~N_N4126);
  assign n1877 = (n1543 | n1562) & (~n1513 | ~N_N4246);
  assign n1878 = n1641 ^ n1947;
  assign n1879 = n1924 ^ ~n1948;
  assign n1880 = (~n1509 | ~N_N3940) & (~NLD3_9 | ~N_N4111);
  assign n1881 = n1880 & (n1583 | ~N_N4218);
  assign n1882 = n1926 ^ ~n1949;
  assign n1883 = n1928 ^ ~n1950;
  assign n1884 = NSr5_7 | PRESET;
  assign n1885 = (~n1509 | ~N_N3923) & (~NLD3_9 | ~N_N3475);
  assign n1886 = n1885 & (n1583 | ~N_N4230);
  assign n1887 = n1795 ^ n1951;
  assign n1888 = (~n1511 | ~N_N3800) & (~N_N3908 | n1971);
  assign n1889 = n1785 ^ n1952;
  assign n1890 = (n1971 | ~N_N3516) & (~n1511 | ~N_N4136);
  assign n1891 = (n1971 | ~N_N3420) & (~n1511 | ~N_N4183);
  assign n1892 = (n1546 | n1560_1) & (~N_N3369 | n1970);
  assign n1893 = n1892 & (n1565_1 | n1803);
  assign n1894 = (~N_N3862 | n1971) & (~n1511 | ~N_N3813);
  assign n1895 = (n1549 | n1560_1) & (~N_N4093 | n1970);
  assign n1896 = n1895 & (n1569 | n1803);
  assign n1897 = (~n1511 | ~N_N4208) & (~N_N4158 | n1971);
  assign n1898 = (~n1511 | ~N_N3807) & (~N_N3713 | n1971);
  assign n1899 = (n1583 | ~N_N3248) & (~n1509 | ~N_N3872);
  assign n1900 = n1899 & (~NLD3_9 | ~N_N3761);
  assign n1901 = N_N3965 ^ n1780;
  assign n1902 = (n1539 | n1562) & (~n1513 | ~N_N4036);
  assign n1903 = (n1535_1 | n1562) & (~n1513 | ~N_N4004);
  assign n1904 = (n1583 | ~N_N3011) & (~n1509 | ~N_N4177);
  assign n1905 = n1904 & (~NLD3_9 | ~N_N3884);
  assign n1906 = (n1555_1 | n1560_1) & (~N_N3283 | n1970);
  assign n1907 = N_N3283 ^ n1564;
  assign n1908 = n1906 & (n1907 | n1803);
  assign n1909 = (~n1511 | ~N_N3470) & (~N_N3821 | n1971);
  assign n1910 = n1789 ^ n1953;
  assign n1911 = n1777 ^ n1972;
  assign n1912 = (n1532 | n1562) & (~n1513 | ~N_N3961);
  assign n1913 = n1791 ^ n1954;
  assign n1914 = (~n1511 | ~N_N3868) & (~N_N3832 | n1971);
  assign n1915 = (~N_N3794 | n1971) & (~n1511 | ~N_N3919);
  assign n1916 = (~n1511 | ~N_N3871) & (~N_N3214 | n1971);
  assign n1175 = n1058 & ~NSr3_9;
  assign n1918 = ~PRESET & Pover_0_0_ & (~NGFDN_3 | NDN3_11);
  assign n1136 = n1175 | n1918;
  assign n1920 = ~PRESET & Pnext_0_0_ & (~NLD3_9 | NDN5_16);
  assign n1440 = ~PRESET & n1957;
  assign n373 = n1920 | n1440;
  assign n1923 = N_N3283 | n1564;
  assign n1924 = n1612 ^ n1596;
  assign n1925 = n1619 ^ n1598;
  assign n1926 = n1620 ^ n1594;
  assign n1927 = n1627 ^ n1599;
  assign n1928 = n1628 ^ n1593;
  assign n1929 = n1604 ^ n1600;
  assign n1930 = n1604 & n1600 & n1592;
  assign n1931 = n1930 ^ n1601;
  assign n1932 = n1642 ^ n1643;
  assign n1933 = n1590 ^ n1979;
  assign n1934 = n1932 ^ n1933;
  assign n1935 = n1633 ^ n1603;
  assign n1936 = n1750 ^ ~N_N4197;
  assign n1937 = n1615 ^ n1606;
  assign n1938 = n1622 ^ n1623;
  assign n1939 = n1630 ^ n1631;
  assign n1940 = n1636 ^ n1637;
  assign n1941 = n1774 ^ ~N_N3992;
  assign n1942 = n1768 ^ ~N_N4018;
  assign n1943 = n1759 ^ ~N_N3949;
  assign n1944 = n1679 ^ n1680;
  assign n1945 = n1651 | n1650;
  assign n1946 = n1753 ^ ~N_N3912;
  assign n1947 = n1639 ^ n1602;
  assign n1948 = n1611 ^ n1613;
  assign n1949 = n1617 ^ n1618;
  assign n1950 = n1625 ^ n1626;
  assign n1951 = n1756 ^ ~N_N4145;
  assign n1952 = n1771 ^ ~N_N3996;
  assign n1953 = n1765 ^ ~N_N3974;
  assign n1954 = n1762 ^ ~N_N4083;
  assign n1955 = n947 & ~N_N4214;
  assign n1956 = n1571 & n1573 & n1575_1 & n1565_1 & n1569 & n1567;
  assign n1957 = ~NLD3_9 & NDN5_9;
  assign n1958 = ~PDN | NDN1_4;
  assign n1959 = (~Preset_0_0_ & (~NLC1_2 | N_N3998)) | (NLC1_2 & N_N3998);
  assign n1960 = ~NDN3_3 & ~NSr3_2;
  assign n1961 = NDN2_2 | n1169;
  assign n1962 = ~PRESET & n1589;
  assign n1963 = n1601 & n1930;
  assign n1964 = NSr5_8 | NDN5_8;
  assign n1965 = NSr5_4 | NDN5_4;
  assign n1966 = NSr5_7 | NDN5_7;
  assign n1967 = NSr5_3 | NDN5_3;
  assign n1968 = NSr5_5 | NDN5_5;
  assign n1969 = NSr5_2 | NDN5_2;
  assign n1970 = ~n1557 | n1559;
  assign n1971 = PRESET | ~NLD3_9;
  assign n1972 = n1781 ^ ~N_N4027;
  assign n1973 = n1976 & (PRESET | n1805 | ~N_N4227);
  assign n273 = ~n1973;
  assign n1975 = n1532 & n1535_1 & n1539 & n1522 & n1529 & n1525_1;
  assign n1976 = ~n1804 | n1807 | N_N4227;
  assign n1480 = ~n1884;
  assign n1485 = ~n1830;
  assign n1979 = n1963 & n1591;
  assign n1980 = n1595 | n1607;
  assign n1981 = n1671 ^ n1672;
  assign n1982 = n1675 ^ n1676;
  assign n1983 = n1704 ^ n1705;
  assign n1984 = n1608 ^ n1980;
  assign n1985 = n1686 ^ n1687;
  assign n1986 = n1694 ^ n1695;
  assign n1987 = n1673 ^ n1674;
  assign n1988 = n1690 ^ n1691;
  assign n1989 = n1677 ^ n1678;
  assign n1990 = n1698 ^ n1699;
  assign n1991 = n1858 ^ n1859;
  assign n1992 = n1975 & n1555_1 & n1552 & n1546 & ~N_N3999 & n1519 & n1543 & n1549;
  assign n1993 = ~Preset_0_0_ & n1833;
  always @ (posedge clk) begin
    N_N4054 <= n63_1;
    N_N3745 <= n68_1;
    N_N4119 <= n73_1;
    N_N3826 <= n78_1;
    N_N3818 <= n83_1;
    N_N3345 <= n88;
    N_N3924 <= n93_1;
    N_N3815 <= n98_1;
    N_N3691 <= n103;
    N_N3157 <= n108_1;
    N_N3872 <= n113_1;
    N_N3788 <= n118_1;
    N_N3375 <= n123_1;
    N_N3143 <= n128;
    N_N4197 <= n133;
    N_N3843 <= n138_1;
    N_N3426 <= n143_1;
    N_N4118 <= n148_1;
    N_N3580 <= n153_1;
    N_N3175 <= n158_1;
    N_N3071 <= n163_1;
    N_N3808 <= n168_1;
    N_N3923 <= n173_1;
    N_N3250 <= n178_1;
    N_N4221 <= n183_1;
    N_N3069 <= n188_1;
    N_N3464 <= n193_1;
    N_N3535 <= n198_1;
    N_N3871 <= n203_1;
    N_N3248 <= n208_1;
    N_N4180 <= n213_1;
    N_N3311 <= n218_1;
    N_N3442 <= n223_1;
    N_N3981 <= n228_1;
    N_N3842 <= n233;
    N_N3105 <= n238;
    N_N4133 <= n243_1;
    N_N4117 <= n248_1;
    N_N3420 <= n253_1;
    N_N3761 <= n258_1;
    N_N3062 <= n263_1;
    N_N4071 <= n268;
    N_N4227 <= n273;
    N_N3807 <= n278_1;
    N_N4145 <= n283;
    N_N3922 <= n288_1;
    N_N3516 <= n293;
    N_N3489 <= n298;
    N_N4030 <= n303_1;
    N_N3540 <= n308_1;
    N_N3513 <= n313_1;
    N_N4083 <= n318_1;
    N_N3841 <= n323_1;
    N_N4018 <= n328_1;
    N_N3971 <= n333_1;
    N_N4232 <= n338_1;
    N_N4246 <= n343_1;
    N_N3806 <= n348_1;
    N_N3992 <= n353_1;
    N_N4086 <= n358_1;
    N_N4230 <= n363_1;
    N_N4212 <= n368;
    Pnext_0_0_ <= n373;
    N_N3626 <= n377;
    N_N3965 <= n382_1;
    N_N3890 <= n387_1;
    NDN3_11 <= n392_1;
    NDN5_10 <= n397_1;
    N_N3786 <= n402_1;
    N_N4171 <= n407;
    NDN5_16 <= n412_1;
    N_N3799 <= n417_1;
    N_N3844 <= n422_1;
    N_N3196 <= n427;
    N_N4126 <= n432_1;
    N_N3681 <= n437_1;
    N_N3679 <= n442;
    N_N3340 <= n447;
    N_N4116 <= n452_1;
    N_N3810 <= n457;
    N_N3235 <= n462;
    N_N3283 <= n467;
    N_N3716 <= n472;
    N_N3701 <= n477;
    N_N3921 <= n482;
    N_N3625 <= n487_1;
    N_N3751 <= n492;
    N_N3736 <= n497;
    N_N3870 <= n502_1;
    N_N4024 <= n507;
    N_N3876 <= n512;
    N_N3840 <= n517_1;
    N_N4021 <= n522_1;
    N_N3932 <= n527;
    NLC1_2 <= n532;
    N_N3805 <= n537_1;
    N_N3700 <= n542_1;
    N_N3735 <= n547;
    NLak3_2 <= n552;
    NLak3_9 <= n557_1;
    N_N3906 <= n562;
    N_N3388 <= n567_1;
    N_N4057 <= n572;
    N_N3011 <= n577_1;
    N_N3346 <= n582;
    N_N3677 <= n587;
    N_N4165 <= n592;
    N_N4080 <= n597_1;
    N_N3373 <= n602_1;
    N_N3709 <= n607_1;
    N_N4206 <= n612;
    N_N3324 <= n617;
    N_N3575 <= n622;
    N_N4159 <= n627;
    NAK5_2 <= n632;
    N_N3916 <= n637_1;
    N_N3743 <= n642_1;
    N_N4242 <= n647;
    N_N3312 <= n652;
    N_N3733 <= n657;
    N_N3774 <= n662_1;
    N_N4214 <= n667;
    N_N3294 <= n672;
    N_N3796 <= n677;
    N_N3574 <= n682_1;
    N_N3791 <= n687_1;
    N_N3480 <= n692;
    N_N4243 <= n697;
    N_N3940 <= n702_1;
    N_N3509 <= n707;
    N_N4015 <= n712_1;
    N_N2989 <= n717;
    N_N3919 <= n722_1;
    N_N3578 <= n727_1;
    N_N3529 <= n732;
    N_N4222 <= n737;
    N_N3910 <= n742_1;
    N_N3868 <= n747;
    N_N3947 <= n752_1;
    N_N4181 <= n757;
    N_N3793 <= n762;
    N_N3822 <= n767_1;
    N_N3813 <= n772;
    N_N4114 <= n777;
    N_N4134 <= n782;
    N_N3866 <= n787;
    N_N4218 <= n792;
    N_N3939 <= n797;
    N_N3776 <= n802_1;
    N_N3387 <= n807_1;
    N_N4194 <= n812_1;
    N_N3821 <= n817;
    N_N3882 <= n822_1;
    N_N4167 <= n827_1;
    N_N3800 <= n832_1;
    N_N4237 <= n837;
    N_N3417 <= n842_1;
    N_N3918 <= n847_1;
    N_N4158 <= n852_1;
    N_N3630 <= n857_1;
    N_N3344 <= n862;
    N_N4072 <= n867_1;
    N_N3274 <= n872_1;
    N_N3473 <= n877;
    N_N4205 <= n882_1;
    N_N4111 <= n887_1;
    N_N3680 <= n892_1;
    N_N3838 <= n897_1;
    N_N3262 <= n902;
    N_N4099 <= n907;
    N_N3607 <= n912;
    N_N3323 <= n917;
    N_N3612 <= n922;
    N_N4079 <= n927_1;
    PDN <= n932_1;
    N_N3457 <= n936;
    N_N3445 <= n941;
    N_N3794 <= n946_1;
    N_N3663 <= n951_1;
    N_N3715 <= n956_1;
    N_N4039 <= n961_1;
    N_N3280 <= n966_1;
    N_N4239 <= n971_1;
    N_N3988 <= n976;
    N_N3433 <= n981_1;
    N_N4075 <= n986;
    N_N3468 <= n991_1;
    N_N4045 <= n996;
    N_N3482 <= n1001_1;
    N_N3832 <= n1006_1;
    N_N3304 <= n1011;
    N_N3750 <= n1016_1;
    N_N3634 <= n1021;
    N_N3293 <= n1026;
    N_N3659 <= n1031_1;
    N_N4252 <= n1036;
    N_N3912 <= n1041_1;
    N_N3862 <= n1046;
    N_N3221 <= n1051_1;
    N_N3875 <= n1056;
    N_N3949 <= n1061_1;
    N_N3908 <= n1066_1;
    N_N3711 <= n1071;
    N_N3931 <= n1076;
    N_N3469 <= n1081_1;
    N_N3436 <= n1086_1;
    N_N3974 <= n1091_1;
    N_N3905 <= n1096;
    N_N3741 <= n1101;
    N_N3369 <= n1106;
    N_N3164 <= n1111;
    N_N3500 <= n1116_1;
    N_N3996 <= n1121;
    N_N3356 <= n1126;
    N_N4093 <= n1131;
    Pover_0_0_ <= n1136;
    N_N4224 <= n1140;
    N_N4027 <= n1145;
    NDN1_4 <= n1150;
    N_N3384 <= n1155;
    N_N4036 <= n1160;
    N_N3968 <= n1165;
    N_N4183 <= n1170;
    NGFDN_3 <= n1175;
    N_N4090 <= n1180_1;
    N_N4004 <= n1185_1;
    N_N3205 <= n1190;
    N_N4136 <= n1195_1;
    N_N3303 <= n1200_1;
    N_N3533 <= n1205_1;
    N_N3336 <= n1210_1;
    N_N3961 <= n1215;
    N_N3331 <= n1220;
    N_N3203 <= n1225;
    N_N4236 <= n1230_1;
    N_N3884 <= n1235_1;
    N_N3367 <= n1240;
    N_N4140 <= n1245_1;
    NDN2_2 <= n1250_1;
    N_N4106 <= n1255;
    N_N3100 <= n1260;
    N_N4193 <= n1265;
    N_N3470 <= n1270;
    N_N3424 <= n1275_1;
    N_N3959 <= n1280;
    N_N3393 <= n1285_1;
    N_N4042 <= n1290_1;
    N_N3188 <= n1295_1;
    N_N4095 <= n1300;
    N_N3957 <= n1305;
    N_N3517 <= n1310;
    N_N4047 <= n1315;
    N_N3081 <= n1320;
    N_N3541 <= n1325;
    N_N4177 <= n1330;
    NDN3_3 <= n1335;
    N_N4176 <= n1340;
    N_N3585 <= n1345;
    NDN3_8 <= n1350;
    N_N4209 <= n1355;
    N_N3824 <= n1360;
    N_N4208 <= n1365;
    N_N4120 <= n1370;
    N_N3708 <= n1375;
    N_N4220 <= n1380;
    N_N3999 <= n1385;
    N_N4223 <= n1390;
    N_N3179 <= n1395;
    N_N4179 <= n1400;
    N_N3475 <= n1405;
    N_N4132 <= n1410;
    N_N4182 <= n1415;
    N_N3797 <= n1420;
    N_N3214 <= n1425;
    N_N4070 <= n1430;
    N_N4135 <= n1435;
    NLD3_9 <= n1440;
    NDN5_2 <= n1445;
    NDN5_3 <= n1450;
    N_N3778 <= n1455;
    NDN5_4 <= n1460;
    N_N3212 <= n1465;
    NDN5_5 <= n1470;
    NDN5_6 <= n1475;
    NDN5_7 <= n1480;
    NDN5_8 <= n1485;
    N_N4073 <= n1490;
    NDN5_9 <= n1495;
    NEN5_9 <= n1500;
    N_N3684 <= n1505;
    N_N4056 <= n1510;
    N_N3713 <= n1515;
    N_N3829 <= n1520;
    N_N4060 <= n1525;
    NSr3_2 <= n1530;
    NSr5_2 <= n1535;
    NSr5_3 <= n1540;
    N_N3462 <= n1545;
    N_N3460 <= n1550;
    NSr5_4 <= n1555;
    NSr3_9 <= n1560;
    NSr5_5 <= n1565;
    NSr5_7 <= n1570;
    NSr5_8 <= n1575;
    N_N3998 <= n1580;
  end
endmodule


