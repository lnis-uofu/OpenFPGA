`include "./ff_checker.sv"
