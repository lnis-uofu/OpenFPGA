*****************************
*     FPGA SPICE Netlist    *
* Description: Switch Block  [1][0] in FPGA *
*    Author: Xifan TANG     *
* Organization: EPFL/IC/LSI *
* Date: Thu Nov 15 14:26:08 2018
 *
*****************************
***** Switch Box[1][0] Sub-Circuit *****
.subckt sb[1][0] 
***** Inputs/outputs of top side *****
+ chany[1][1]_out[0] chany[1][1]_in[1] chany[1][1]_out[2] chany[1][1]_in[3] chany[1][1]_out[4] chany[1][1]_in[5] chany[1][1]_out[6] chany[1][1]_in[7] chany[1][1]_out[8] chany[1][1]_in[9] chany[1][1]_out[10] chany[1][1]_in[11] chany[1][1]_out[12] chany[1][1]_in[13] chany[1][1]_out[14] chany[1][1]_in[15] chany[1][1]_out[16] chany[1][1]_in[17] chany[1][1]_out[18] chany[1][1]_in[19] chany[1][1]_out[20] chany[1][1]_in[21] chany[1][1]_out[22] chany[1][1]_in[23] chany[1][1]_out[24] chany[1][1]_in[25] chany[1][1]_out[26] chany[1][1]_in[27] chany[1][1]_out[28] chany[1][1]_in[29] chany[1][1]_out[30] chany[1][1]_in[31] chany[1][1]_out[32] chany[1][1]_in[33] chany[1][1]_out[34] chany[1][1]_in[35] chany[1][1]_out[36] chany[1][1]_in[37] chany[1][1]_out[38] chany[1][1]_in[39] chany[1][1]_out[40] chany[1][1]_in[41] chany[1][1]_out[42] chany[1][1]_in[43] chany[1][1]_out[44] chany[1][1]_in[45] chany[1][1]_out[46] chany[1][1]_in[47] chany[1][1]_out[48] chany[1][1]_in[49] chany[1][1]_out[50] chany[1][1]_in[51] chany[1][1]_out[52] chany[1][1]_in[53] chany[1][1]_out[54] chany[1][1]_in[55] chany[1][1]_out[56] chany[1][1]_in[57] chany[1][1]_out[58] chany[1][1]_in[59] chany[1][1]_out[60] chany[1][1]_in[61] chany[1][1]_out[62] chany[1][1]_in[63] chany[1][1]_out[64] chany[1][1]_in[65] chany[1][1]_out[66] chany[1][1]_in[67] chany[1][1]_out[68] chany[1][1]_in[69] chany[1][1]_out[70] chany[1][1]_in[71] chany[1][1]_out[72] chany[1][1]_in[73] chany[1][1]_out[74] chany[1][1]_in[75] chany[1][1]_out[76] chany[1][1]_in[77] chany[1][1]_out[78] chany[1][1]_in[79] chany[1][1]_out[80] chany[1][1]_in[81] chany[1][1]_out[82] chany[1][1]_in[83] chany[1][1]_out[84] chany[1][1]_in[85] chany[1][1]_out[86] chany[1][1]_in[87] chany[1][1]_out[88] chany[1][1]_in[89] chany[1][1]_out[90] chany[1][1]_in[91] chany[1][1]_out[92] chany[1][1]_in[93] chany[1][1]_out[94] chany[1][1]_in[95] chany[1][1]_out[96] chany[1][1]_in[97] chany[1][1]_out[98] chany[1][1]_in[99] 
+ grid[1][1]_pin[0][1][41] grid[1][1]_pin[0][1][45] grid[1][1]_pin[0][1][49] grid[2][1]_pin[0][3][1] grid[2][1]_pin[0][3][3] grid[2][1]_pin[0][3][5] grid[2][1]_pin[0][3][7] grid[2][1]_pin[0][3][9] grid[2][1]_pin[0][3][11] grid[2][1]_pin[0][3][13] grid[2][1]_pin[0][3][15] 
+ ***** Inputs/outputs of right side *****
+ 
+ 
+ ***** Inputs/outputs of bottom side *****
+ 
+ 
+ ***** Inputs/outputs of left side *****
+ chanx[1][0]_in[0] chanx[1][0]_out[1] chanx[1][0]_in[2] chanx[1][0]_out[3] chanx[1][0]_in[4] chanx[1][0]_out[5] chanx[1][0]_in[6] chanx[1][0]_out[7] chanx[1][0]_in[8] chanx[1][0]_out[9] chanx[1][0]_in[10] chanx[1][0]_out[11] chanx[1][0]_in[12] chanx[1][0]_out[13] chanx[1][0]_in[14] chanx[1][0]_out[15] chanx[1][0]_in[16] chanx[1][0]_out[17] chanx[1][0]_in[18] chanx[1][0]_out[19] chanx[1][0]_in[20] chanx[1][0]_out[21] chanx[1][0]_in[22] chanx[1][0]_out[23] chanx[1][0]_in[24] chanx[1][0]_out[25] chanx[1][0]_in[26] chanx[1][0]_out[27] chanx[1][0]_in[28] chanx[1][0]_out[29] chanx[1][0]_in[30] chanx[1][0]_out[31] chanx[1][0]_in[32] chanx[1][0]_out[33] chanx[1][0]_in[34] chanx[1][0]_out[35] chanx[1][0]_in[36] chanx[1][0]_out[37] chanx[1][0]_in[38] chanx[1][0]_out[39] chanx[1][0]_in[40] chanx[1][0]_out[41] chanx[1][0]_in[42] chanx[1][0]_out[43] chanx[1][0]_in[44] chanx[1][0]_out[45] chanx[1][0]_in[46] chanx[1][0]_out[47] chanx[1][0]_in[48] chanx[1][0]_out[49] chanx[1][0]_in[50] chanx[1][0]_out[51] chanx[1][0]_in[52] chanx[1][0]_out[53] chanx[1][0]_in[54] chanx[1][0]_out[55] chanx[1][0]_in[56] chanx[1][0]_out[57] chanx[1][0]_in[58] chanx[1][0]_out[59] chanx[1][0]_in[60] chanx[1][0]_out[61] chanx[1][0]_in[62] chanx[1][0]_out[63] chanx[1][0]_in[64] chanx[1][0]_out[65] chanx[1][0]_in[66] chanx[1][0]_out[67] chanx[1][0]_in[68] chanx[1][0]_out[69] chanx[1][0]_in[70] chanx[1][0]_out[71] chanx[1][0]_in[72] chanx[1][0]_out[73] chanx[1][0]_in[74] chanx[1][0]_out[75] chanx[1][0]_in[76] chanx[1][0]_out[77] chanx[1][0]_in[78] chanx[1][0]_out[79] chanx[1][0]_in[80] chanx[1][0]_out[81] chanx[1][0]_in[82] chanx[1][0]_out[83] chanx[1][0]_in[84] chanx[1][0]_out[85] chanx[1][0]_in[86] chanx[1][0]_out[87] chanx[1][0]_in[88] chanx[1][0]_out[89] chanx[1][0]_in[90] chanx[1][0]_out[91] chanx[1][0]_in[92] chanx[1][0]_out[93] chanx[1][0]_in[94] chanx[1][0]_out[95] chanx[1][0]_in[96] chanx[1][0]_out[97] chanx[1][0]_in[98] chanx[1][0]_out[99] 
+ grid[1][1]_pin[0][2][42] grid[1][1]_pin[0][2][46] grid[1][0]_pin[0][0][1] grid[1][0]_pin[0][0][3] grid[1][0]_pin[0][0][5] grid[1][0]_pin[0][0][7] grid[1][0]_pin[0][0][9] grid[1][0]_pin[0][0][11] grid[1][0]_pin[0][0][13] grid[1][0]_pin[0][0][15] 
+ svdd sgnd
***** top side Multiplexers *****
Xmux_1level_tapbuf_size3[210] grid[1][1]_pin[0][1][41] grid[2][1]_pin[0][3][15] chanx[1][0]_in[0] chany[1][1]_out[0] sram[1852]->outb sram[1852]->out sram[1853]->out sram[1853]->outb sram[1854]->out sram[1854]->outb svdd sgnd mux_1level_tapbuf_size3
***** SRAM bits for MUX[210], level=1, select_path_id=0. *****
*****100*****
Xsram[1852] sram->in sram[1852]->out sram[1852]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1852]->out) 0
.nodeset V(sram[1852]->outb) vsp
Xsram[1853] sram->in sram[1853]->out sram[1853]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1853]->out) 0
.nodeset V(sram[1853]->outb) vsp
Xsram[1854] sram->in sram[1854]->out sram[1854]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1854]->out) 0
.nodeset V(sram[1854]->outb) vsp
Xmux_1level_tapbuf_size3[211] grid[1][1]_pin[0][1][41] grid[2][1]_pin[0][3][15] chanx[1][0]_in[98] chany[1][1]_out[2] sram[1855]->outb sram[1855]->out sram[1856]->out sram[1856]->outb sram[1857]->out sram[1857]->outb svdd sgnd mux_1level_tapbuf_size3
***** SRAM bits for MUX[211], level=1, select_path_id=0. *****
*****100*****
Xsram[1855] sram->in sram[1855]->out sram[1855]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1855]->out) 0
.nodeset V(sram[1855]->outb) vsp
Xsram[1856] sram->in sram[1856]->out sram[1856]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1856]->out) 0
.nodeset V(sram[1856]->outb) vsp
Xsram[1857] sram->in sram[1857]->out sram[1857]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1857]->out) 0
.nodeset V(sram[1857]->outb) vsp
Xmux_1level_tapbuf_size3[212] grid[1][1]_pin[0][1][41] grid[2][1]_pin[0][3][15] chanx[1][0]_in[96] chany[1][1]_out[4] sram[1858]->outb sram[1858]->out sram[1859]->out sram[1859]->outb sram[1860]->out sram[1860]->outb svdd sgnd mux_1level_tapbuf_size3
***** SRAM bits for MUX[212], level=1, select_path_id=0. *****
*****100*****
Xsram[1858] sram->in sram[1858]->out sram[1858]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1858]->out) 0
.nodeset V(sram[1858]->outb) vsp
Xsram[1859] sram->in sram[1859]->out sram[1859]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1859]->out) 0
.nodeset V(sram[1859]->outb) vsp
Xsram[1860] sram->in sram[1860]->out sram[1860]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1860]->out) 0
.nodeset V(sram[1860]->outb) vsp
Xmux_1level_tapbuf_size3[213] grid[1][1]_pin[0][1][41] grid[2][1]_pin[0][3][15] chanx[1][0]_in[94] chany[1][1]_out[6] sram[1861]->outb sram[1861]->out sram[1862]->out sram[1862]->outb sram[1863]->out sram[1863]->outb svdd sgnd mux_1level_tapbuf_size3
***** SRAM bits for MUX[213], level=1, select_path_id=0. *****
*****100*****
Xsram[1861] sram->in sram[1861]->out sram[1861]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1861]->out) 0
.nodeset V(sram[1861]->outb) vsp
Xsram[1862] sram->in sram[1862]->out sram[1862]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1862]->out) 0
.nodeset V(sram[1862]->outb) vsp
Xsram[1863] sram->in sram[1863]->out sram[1863]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1863]->out) 0
.nodeset V(sram[1863]->outb) vsp
Xmux_1level_tapbuf_size3[214] grid[1][1]_pin[0][1][41] grid[2][1]_pin[0][3][15] chanx[1][0]_in[92] chany[1][1]_out[8] sram[1864]->outb sram[1864]->out sram[1865]->out sram[1865]->outb sram[1866]->out sram[1866]->outb svdd sgnd mux_1level_tapbuf_size3
***** SRAM bits for MUX[214], level=1, select_path_id=0. *****
*****100*****
Xsram[1864] sram->in sram[1864]->out sram[1864]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1864]->out) 0
.nodeset V(sram[1864]->outb) vsp
Xsram[1865] sram->in sram[1865]->out sram[1865]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1865]->out) 0
.nodeset V(sram[1865]->outb) vsp
Xsram[1866] sram->in sram[1866]->out sram[1866]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1866]->out) 0
.nodeset V(sram[1866]->outb) vsp
Xmux_1level_tapbuf_size2[215] grid[1][1]_pin[0][1][45] chanx[1][0]_in[90] chany[1][1]_out[10] sram[1867]->outb sram[1867]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[215], level=1, select_path_id=0. *****
*****1*****
Xsram[1867] sram->in sram[1867]->out sram[1867]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1867]->out) 0
.nodeset V(sram[1867]->outb) vsp
Xmux_1level_tapbuf_size2[216] grid[1][1]_pin[0][1][45] chanx[1][0]_in[88] chany[1][1]_out[12] sram[1868]->outb sram[1868]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[216], level=1, select_path_id=0. *****
*****1*****
Xsram[1868] sram->in sram[1868]->out sram[1868]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1868]->out) 0
.nodeset V(sram[1868]->outb) vsp
Xmux_1level_tapbuf_size2[217] grid[1][1]_pin[0][1][45] chanx[1][0]_in[86] chany[1][1]_out[14] sram[1869]->outb sram[1869]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[217], level=1, select_path_id=0. *****
*****1*****
Xsram[1869] sram->in sram[1869]->out sram[1869]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1869]->out) 0
.nodeset V(sram[1869]->outb) vsp
Xmux_1level_tapbuf_size2[218] grid[1][1]_pin[0][1][45] chanx[1][0]_in[84] chany[1][1]_out[16] sram[1870]->outb sram[1870]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[218], level=1, select_path_id=0. *****
*****1*****
Xsram[1870] sram->in sram[1870]->out sram[1870]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1870]->out) 0
.nodeset V(sram[1870]->outb) vsp
Xmux_1level_tapbuf_size2[219] grid[1][1]_pin[0][1][45] chanx[1][0]_in[82] chany[1][1]_out[18] sram[1871]->outb sram[1871]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[219], level=1, select_path_id=0. *****
*****1*****
Xsram[1871] sram->in sram[1871]->out sram[1871]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1871]->out) 0
.nodeset V(sram[1871]->outb) vsp
Xmux_1level_tapbuf_size2[220] grid[1][1]_pin[0][1][49] chanx[1][0]_in[80] chany[1][1]_out[20] sram[1872]->outb sram[1872]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[220], level=1, select_path_id=0. *****
*****1*****
Xsram[1872] sram->in sram[1872]->out sram[1872]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1872]->out) 0
.nodeset V(sram[1872]->outb) vsp
Xmux_1level_tapbuf_size2[221] grid[1][1]_pin[0][1][49] chanx[1][0]_in[78] chany[1][1]_out[22] sram[1873]->outb sram[1873]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[221], level=1, select_path_id=0. *****
*****1*****
Xsram[1873] sram->in sram[1873]->out sram[1873]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1873]->out) 0
.nodeset V(sram[1873]->outb) vsp
Xmux_1level_tapbuf_size2[222] grid[1][1]_pin[0][1][49] chanx[1][0]_in[76] chany[1][1]_out[24] sram[1874]->outb sram[1874]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[222], level=1, select_path_id=0. *****
*****1*****
Xsram[1874] sram->in sram[1874]->out sram[1874]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1874]->out) 0
.nodeset V(sram[1874]->outb) vsp
Xmux_1level_tapbuf_size2[223] grid[1][1]_pin[0][1][49] chanx[1][0]_in[74] chany[1][1]_out[26] sram[1875]->outb sram[1875]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[223], level=1, select_path_id=0. *****
*****1*****
Xsram[1875] sram->in sram[1875]->out sram[1875]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1875]->out) 0
.nodeset V(sram[1875]->outb) vsp
Xmux_1level_tapbuf_size2[224] grid[1][1]_pin[0][1][49] chanx[1][0]_in[72] chany[1][1]_out[28] sram[1876]->outb sram[1876]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[224], level=1, select_path_id=0. *****
*****1*****
Xsram[1876] sram->in sram[1876]->out sram[1876]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1876]->out) 0
.nodeset V(sram[1876]->outb) vsp
Xmux_1level_tapbuf_size2[225] grid[2][1]_pin[0][3][1] chanx[1][0]_in[70] chany[1][1]_out[30] sram[1877]->outb sram[1877]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[225], level=1, select_path_id=0. *****
*****1*****
Xsram[1877] sram->in sram[1877]->out sram[1877]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1877]->out) 0
.nodeset V(sram[1877]->outb) vsp
Xmux_1level_tapbuf_size2[226] grid[2][1]_pin[0][3][1] chanx[1][0]_in[68] chany[1][1]_out[32] sram[1878]->outb sram[1878]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[226], level=1, select_path_id=0. *****
*****1*****
Xsram[1878] sram->in sram[1878]->out sram[1878]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1878]->out) 0
.nodeset V(sram[1878]->outb) vsp
Xmux_1level_tapbuf_size2[227] grid[2][1]_pin[0][3][1] chanx[1][0]_in[66] chany[1][1]_out[34] sram[1879]->outb sram[1879]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[227], level=1, select_path_id=0. *****
*****1*****
Xsram[1879] sram->in sram[1879]->out sram[1879]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1879]->out) 0
.nodeset V(sram[1879]->outb) vsp
Xmux_1level_tapbuf_size2[228] grid[2][1]_pin[0][3][1] chanx[1][0]_in[64] chany[1][1]_out[36] sram[1880]->outb sram[1880]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[228], level=1, select_path_id=0. *****
*****1*****
Xsram[1880] sram->in sram[1880]->out sram[1880]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1880]->out) 0
.nodeset V(sram[1880]->outb) vsp
Xmux_1level_tapbuf_size2[229] grid[2][1]_pin[0][3][1] chanx[1][0]_in[62] chany[1][1]_out[38] sram[1881]->outb sram[1881]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[229], level=1, select_path_id=0. *****
*****1*****
Xsram[1881] sram->in sram[1881]->out sram[1881]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1881]->out) 0
.nodeset V(sram[1881]->outb) vsp
Xmux_1level_tapbuf_size2[230] grid[2][1]_pin[0][3][3] chanx[1][0]_in[60] chany[1][1]_out[40] sram[1882]->outb sram[1882]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[230], level=1, select_path_id=0. *****
*****1*****
Xsram[1882] sram->in sram[1882]->out sram[1882]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1882]->out) 0
.nodeset V(sram[1882]->outb) vsp
Xmux_1level_tapbuf_size2[231] grid[2][1]_pin[0][3][3] chanx[1][0]_in[58] chany[1][1]_out[42] sram[1883]->outb sram[1883]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[231], level=1, select_path_id=0. *****
*****1*****
Xsram[1883] sram->in sram[1883]->out sram[1883]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1883]->out) 0
.nodeset V(sram[1883]->outb) vsp
Xmux_1level_tapbuf_size2[232] grid[2][1]_pin[0][3][3] chanx[1][0]_in[56] chany[1][1]_out[44] sram[1884]->outb sram[1884]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[232], level=1, select_path_id=0. *****
*****1*****
Xsram[1884] sram->in sram[1884]->out sram[1884]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1884]->out) 0
.nodeset V(sram[1884]->outb) vsp
Xmux_1level_tapbuf_size2[233] grid[2][1]_pin[0][3][3] chanx[1][0]_in[54] chany[1][1]_out[46] sram[1885]->outb sram[1885]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[233], level=1, select_path_id=0. *****
*****1*****
Xsram[1885] sram->in sram[1885]->out sram[1885]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1885]->out) 0
.nodeset V(sram[1885]->outb) vsp
Xmux_1level_tapbuf_size2[234] grid[2][1]_pin[0][3][3] chanx[1][0]_in[52] chany[1][1]_out[48] sram[1886]->outb sram[1886]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[234], level=1, select_path_id=0. *****
*****1*****
Xsram[1886] sram->in sram[1886]->out sram[1886]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1886]->out) 0
.nodeset V(sram[1886]->outb) vsp
Xmux_1level_tapbuf_size2[235] grid[2][1]_pin[0][3][5] chanx[1][0]_in[50] chany[1][1]_out[50] sram[1887]->outb sram[1887]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[235], level=1, select_path_id=0. *****
*****1*****
Xsram[1887] sram->in sram[1887]->out sram[1887]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1887]->out) 0
.nodeset V(sram[1887]->outb) vsp
Xmux_1level_tapbuf_size2[236] grid[2][1]_pin[0][3][5] chanx[1][0]_in[48] chany[1][1]_out[52] sram[1888]->outb sram[1888]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[236], level=1, select_path_id=0. *****
*****1*****
Xsram[1888] sram->in sram[1888]->out sram[1888]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1888]->out) 0
.nodeset V(sram[1888]->outb) vsp
Xmux_1level_tapbuf_size2[237] grid[2][1]_pin[0][3][5] chanx[1][0]_in[46] chany[1][1]_out[54] sram[1889]->outb sram[1889]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[237], level=1, select_path_id=0. *****
*****1*****
Xsram[1889] sram->in sram[1889]->out sram[1889]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1889]->out) 0
.nodeset V(sram[1889]->outb) vsp
Xmux_1level_tapbuf_size2[238] grid[2][1]_pin[0][3][5] chanx[1][0]_in[44] chany[1][1]_out[56] sram[1890]->outb sram[1890]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[238], level=1, select_path_id=0. *****
*****1*****
Xsram[1890] sram->in sram[1890]->out sram[1890]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1890]->out) 0
.nodeset V(sram[1890]->outb) vsp
Xmux_1level_tapbuf_size2[239] grid[2][1]_pin[0][3][5] chanx[1][0]_in[42] chany[1][1]_out[58] sram[1891]->outb sram[1891]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[239], level=1, select_path_id=0. *****
*****1*****
Xsram[1891] sram->in sram[1891]->out sram[1891]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1891]->out) 0
.nodeset V(sram[1891]->outb) vsp
Xmux_1level_tapbuf_size2[240] grid[2][1]_pin[0][3][7] chanx[1][0]_in[40] chany[1][1]_out[60] sram[1892]->outb sram[1892]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[240], level=1, select_path_id=0. *****
*****1*****
Xsram[1892] sram->in sram[1892]->out sram[1892]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1892]->out) 0
.nodeset V(sram[1892]->outb) vsp
Xmux_1level_tapbuf_size2[241] grid[2][1]_pin[0][3][7] chanx[1][0]_in[38] chany[1][1]_out[62] sram[1893]->outb sram[1893]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[241], level=1, select_path_id=0. *****
*****1*****
Xsram[1893] sram->in sram[1893]->out sram[1893]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1893]->out) 0
.nodeset V(sram[1893]->outb) vsp
Xmux_1level_tapbuf_size2[242] grid[2][1]_pin[0][3][7] chanx[1][0]_in[36] chany[1][1]_out[64] sram[1894]->outb sram[1894]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[242], level=1, select_path_id=0. *****
*****1*****
Xsram[1894] sram->in sram[1894]->out sram[1894]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1894]->out) 0
.nodeset V(sram[1894]->outb) vsp
Xmux_1level_tapbuf_size2[243] grid[2][1]_pin[0][3][7] chanx[1][0]_in[34] chany[1][1]_out[66] sram[1895]->outb sram[1895]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[243], level=1, select_path_id=0. *****
*****1*****
Xsram[1895] sram->in sram[1895]->out sram[1895]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1895]->out) 0
.nodeset V(sram[1895]->outb) vsp
Xmux_1level_tapbuf_size2[244] grid[2][1]_pin[0][3][7] chanx[1][0]_in[32] chany[1][1]_out[68] sram[1896]->outb sram[1896]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[244], level=1, select_path_id=0. *****
*****1*****
Xsram[1896] sram->in sram[1896]->out sram[1896]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1896]->out) 0
.nodeset V(sram[1896]->outb) vsp
Xmux_1level_tapbuf_size2[245] grid[2][1]_pin[0][3][9] chanx[1][0]_in[30] chany[1][1]_out[70] sram[1897]->outb sram[1897]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[245], level=1, select_path_id=0. *****
*****1*****
Xsram[1897] sram->in sram[1897]->out sram[1897]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1897]->out) 0
.nodeset V(sram[1897]->outb) vsp
Xmux_1level_tapbuf_size2[246] grid[2][1]_pin[0][3][9] chanx[1][0]_in[28] chany[1][1]_out[72] sram[1898]->outb sram[1898]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[246], level=1, select_path_id=0. *****
*****1*****
Xsram[1898] sram->in sram[1898]->out sram[1898]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1898]->out) 0
.nodeset V(sram[1898]->outb) vsp
Xmux_1level_tapbuf_size2[247] grid[2][1]_pin[0][3][9] chanx[1][0]_in[26] chany[1][1]_out[74] sram[1899]->outb sram[1899]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[247], level=1, select_path_id=0. *****
*****1*****
Xsram[1899] sram->in sram[1899]->out sram[1899]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1899]->out) 0
.nodeset V(sram[1899]->outb) vsp
Xmux_1level_tapbuf_size2[248] grid[2][1]_pin[0][3][9] chanx[1][0]_in[24] chany[1][1]_out[76] sram[1900]->outb sram[1900]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[248], level=1, select_path_id=0. *****
*****1*****
Xsram[1900] sram->in sram[1900]->out sram[1900]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1900]->out) 0
.nodeset V(sram[1900]->outb) vsp
Xmux_1level_tapbuf_size2[249] grid[2][1]_pin[0][3][9] chanx[1][0]_in[22] chany[1][1]_out[78] sram[1901]->outb sram[1901]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[249], level=1, select_path_id=0. *****
*****1*****
Xsram[1901] sram->in sram[1901]->out sram[1901]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1901]->out) 0
.nodeset V(sram[1901]->outb) vsp
Xmux_1level_tapbuf_size2[250] grid[2][1]_pin[0][3][11] chanx[1][0]_in[20] chany[1][1]_out[80] sram[1902]->outb sram[1902]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[250], level=1, select_path_id=0. *****
*****1*****
Xsram[1902] sram->in sram[1902]->out sram[1902]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1902]->out) 0
.nodeset V(sram[1902]->outb) vsp
Xmux_1level_tapbuf_size2[251] grid[2][1]_pin[0][3][11] chanx[1][0]_in[18] chany[1][1]_out[82] sram[1903]->outb sram[1903]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[251], level=1, select_path_id=0. *****
*****1*****
Xsram[1903] sram->in sram[1903]->out sram[1903]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1903]->out) 0
.nodeset V(sram[1903]->outb) vsp
Xmux_1level_tapbuf_size2[252] grid[2][1]_pin[0][3][11] chanx[1][0]_in[16] chany[1][1]_out[84] sram[1904]->outb sram[1904]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[252], level=1, select_path_id=0. *****
*****1*****
Xsram[1904] sram->in sram[1904]->out sram[1904]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1904]->out) 0
.nodeset V(sram[1904]->outb) vsp
Xmux_1level_tapbuf_size2[253] grid[2][1]_pin[0][3][11] chanx[1][0]_in[14] chany[1][1]_out[86] sram[1905]->outb sram[1905]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[253], level=1, select_path_id=0. *****
*****1*****
Xsram[1905] sram->in sram[1905]->out sram[1905]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1905]->out) 0
.nodeset V(sram[1905]->outb) vsp
Xmux_1level_tapbuf_size2[254] grid[2][1]_pin[0][3][11] chanx[1][0]_in[12] chany[1][1]_out[88] sram[1906]->outb sram[1906]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[254], level=1, select_path_id=0. *****
*****1*****
Xsram[1906] sram->in sram[1906]->out sram[1906]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1906]->out) 0
.nodeset V(sram[1906]->outb) vsp
Xmux_1level_tapbuf_size2[255] grid[2][1]_pin[0][3][13] chanx[1][0]_in[10] chany[1][1]_out[90] sram[1907]->outb sram[1907]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[255], level=1, select_path_id=0. *****
*****1*****
Xsram[1907] sram->in sram[1907]->out sram[1907]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1907]->out) 0
.nodeset V(sram[1907]->outb) vsp
Xmux_1level_tapbuf_size2[256] grid[2][1]_pin[0][3][13] chanx[1][0]_in[8] chany[1][1]_out[92] sram[1908]->outb sram[1908]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[256], level=1, select_path_id=0. *****
*****1*****
Xsram[1908] sram->in sram[1908]->out sram[1908]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1908]->out) 0
.nodeset V(sram[1908]->outb) vsp
Xmux_1level_tapbuf_size2[257] grid[2][1]_pin[0][3][13] chanx[1][0]_in[6] chany[1][1]_out[94] sram[1909]->outb sram[1909]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[257], level=1, select_path_id=0. *****
*****1*****
Xsram[1909] sram->in sram[1909]->out sram[1909]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1909]->out) 0
.nodeset V(sram[1909]->outb) vsp
Xmux_1level_tapbuf_size2[258] grid[2][1]_pin[0][3][13] chanx[1][0]_in[4] chany[1][1]_out[96] sram[1910]->outb sram[1910]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[258], level=1, select_path_id=0. *****
*****1*****
Xsram[1910] sram->in sram[1910]->out sram[1910]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1910]->out) 0
.nodeset V(sram[1910]->outb) vsp
Xmux_1level_tapbuf_size2[259] grid[2][1]_pin[0][3][13] chanx[1][0]_in[2] chany[1][1]_out[98] sram[1911]->outb sram[1911]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[259], level=1, select_path_id=0. *****
*****1*****
Xsram[1911] sram->in sram[1911]->out sram[1911]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1911]->out) 0
.nodeset V(sram[1911]->outb) vsp
***** right side Multiplexers *****
***** bottom side Multiplexers *****
***** left side Multiplexers *****
Xmux_1level_tapbuf_size2[260] grid[1][0]_pin[0][0][1] chany[1][1]_in[1] chanx[1][0]_out[1] sram[1912]->outb sram[1912]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[260], level=1, select_path_id=0. *****
*****1*****
Xsram[1912] sram->in sram[1912]->out sram[1912]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1912]->out) 0
.nodeset V(sram[1912]->outb) vsp
Xmux_1level_tapbuf_size2[261] grid[1][0]_pin[0][0][1] chany[1][1]_in[99] chanx[1][0]_out[3] sram[1913]->outb sram[1913]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[261], level=1, select_path_id=0. *****
*****1*****
Xsram[1913] sram->in sram[1913]->out sram[1913]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1913]->out) 0
.nodeset V(sram[1913]->outb) vsp
Xmux_1level_tapbuf_size2[262] grid[1][0]_pin[0][0][1] chany[1][1]_in[97] chanx[1][0]_out[5] sram[1914]->outb sram[1914]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[262], level=1, select_path_id=0. *****
*****1*****
Xsram[1914] sram->in sram[1914]->out sram[1914]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1914]->out) 0
.nodeset V(sram[1914]->outb) vsp
Xmux_1level_tapbuf_size2[263] grid[1][0]_pin[0][0][1] chany[1][1]_in[95] chanx[1][0]_out[7] sram[1915]->outb sram[1915]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[263], level=1, select_path_id=0. *****
*****1*****
Xsram[1915] sram->in sram[1915]->out sram[1915]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1915]->out) 0
.nodeset V(sram[1915]->outb) vsp
Xmux_1level_tapbuf_size2[264] grid[1][0]_pin[0][0][1] chany[1][1]_in[93] chanx[1][0]_out[9] sram[1916]->outb sram[1916]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[264], level=1, select_path_id=0. *****
*****1*****
Xsram[1916] sram->in sram[1916]->out sram[1916]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1916]->out) 0
.nodeset V(sram[1916]->outb) vsp
Xmux_1level_tapbuf_size2[265] grid[1][0]_pin[0][0][3] chany[1][1]_in[91] chanx[1][0]_out[11] sram[1917]->outb sram[1917]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[265], level=1, select_path_id=0. *****
*****1*****
Xsram[1917] sram->in sram[1917]->out sram[1917]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1917]->out) 0
.nodeset V(sram[1917]->outb) vsp
Xmux_1level_tapbuf_size2[266] grid[1][0]_pin[0][0][3] chany[1][1]_in[89] chanx[1][0]_out[13] sram[1918]->outb sram[1918]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[266], level=1, select_path_id=0. *****
*****1*****
Xsram[1918] sram->in sram[1918]->out sram[1918]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1918]->out) 0
.nodeset V(sram[1918]->outb) vsp
Xmux_1level_tapbuf_size2[267] grid[1][0]_pin[0][0][3] chany[1][1]_in[87] chanx[1][0]_out[15] sram[1919]->outb sram[1919]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[267], level=1, select_path_id=0. *****
*****1*****
Xsram[1919] sram->in sram[1919]->out sram[1919]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1919]->out) 0
.nodeset V(sram[1919]->outb) vsp
Xmux_1level_tapbuf_size2[268] grid[1][0]_pin[0][0][3] chany[1][1]_in[85] chanx[1][0]_out[17] sram[1920]->outb sram[1920]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[268], level=1, select_path_id=0. *****
*****1*****
Xsram[1920] sram->in sram[1920]->out sram[1920]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1920]->out) 0
.nodeset V(sram[1920]->outb) vsp
Xmux_1level_tapbuf_size2[269] grid[1][0]_pin[0][0][3] chany[1][1]_in[83] chanx[1][0]_out[19] sram[1921]->outb sram[1921]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[269], level=1, select_path_id=0. *****
*****1*****
Xsram[1921] sram->in sram[1921]->out sram[1921]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1921]->out) 0
.nodeset V(sram[1921]->outb) vsp
Xmux_1level_tapbuf_size2[270] grid[1][0]_pin[0][0][5] chany[1][1]_in[81] chanx[1][0]_out[21] sram[1922]->outb sram[1922]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[270], level=1, select_path_id=0. *****
*****1*****
Xsram[1922] sram->in sram[1922]->out sram[1922]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1922]->out) 0
.nodeset V(sram[1922]->outb) vsp
Xmux_1level_tapbuf_size2[271] grid[1][0]_pin[0][0][5] chany[1][1]_in[79] chanx[1][0]_out[23] sram[1923]->outb sram[1923]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[271], level=1, select_path_id=0. *****
*****1*****
Xsram[1923] sram->in sram[1923]->out sram[1923]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1923]->out) 0
.nodeset V(sram[1923]->outb) vsp
Xmux_1level_tapbuf_size2[272] grid[1][0]_pin[0][0][5] chany[1][1]_in[77] chanx[1][0]_out[25] sram[1924]->outb sram[1924]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[272], level=1, select_path_id=0. *****
*****1*****
Xsram[1924] sram->in sram[1924]->out sram[1924]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1924]->out) 0
.nodeset V(sram[1924]->outb) vsp
Xmux_1level_tapbuf_size2[273] grid[1][0]_pin[0][0][5] chany[1][1]_in[75] chanx[1][0]_out[27] sram[1925]->outb sram[1925]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[273], level=1, select_path_id=0. *****
*****1*****
Xsram[1925] sram->in sram[1925]->out sram[1925]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1925]->out) 0
.nodeset V(sram[1925]->outb) vsp
Xmux_1level_tapbuf_size2[274] grid[1][0]_pin[0][0][5] chany[1][1]_in[73] chanx[1][0]_out[29] sram[1926]->outb sram[1926]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[274], level=1, select_path_id=0. *****
*****1*****
Xsram[1926] sram->in sram[1926]->out sram[1926]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1926]->out) 0
.nodeset V(sram[1926]->outb) vsp
Xmux_1level_tapbuf_size2[275] grid[1][0]_pin[0][0][7] chany[1][1]_in[71] chanx[1][0]_out[31] sram[1927]->outb sram[1927]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[275], level=1, select_path_id=0. *****
*****1*****
Xsram[1927] sram->in sram[1927]->out sram[1927]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1927]->out) 0
.nodeset V(sram[1927]->outb) vsp
Xmux_1level_tapbuf_size2[276] grid[1][0]_pin[0][0][7] chany[1][1]_in[69] chanx[1][0]_out[33] sram[1928]->outb sram[1928]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[276], level=1, select_path_id=0. *****
*****1*****
Xsram[1928] sram->in sram[1928]->out sram[1928]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1928]->out) 0
.nodeset V(sram[1928]->outb) vsp
Xmux_1level_tapbuf_size2[277] grid[1][0]_pin[0][0][7] chany[1][1]_in[67] chanx[1][0]_out[35] sram[1929]->outb sram[1929]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[277], level=1, select_path_id=0. *****
*****1*****
Xsram[1929] sram->in sram[1929]->out sram[1929]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1929]->out) 0
.nodeset V(sram[1929]->outb) vsp
Xmux_1level_tapbuf_size2[278] grid[1][0]_pin[0][0][7] chany[1][1]_in[65] chanx[1][0]_out[37] sram[1930]->outb sram[1930]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[278], level=1, select_path_id=0. *****
*****1*****
Xsram[1930] sram->in sram[1930]->out sram[1930]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1930]->out) 0
.nodeset V(sram[1930]->outb) vsp
Xmux_1level_tapbuf_size2[279] grid[1][0]_pin[0][0][7] chany[1][1]_in[63] chanx[1][0]_out[39] sram[1931]->outb sram[1931]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[279], level=1, select_path_id=0. *****
*****1*****
Xsram[1931] sram->in sram[1931]->out sram[1931]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1931]->out) 0
.nodeset V(sram[1931]->outb) vsp
Xmux_1level_tapbuf_size2[280] grid[1][0]_pin[0][0][9] chany[1][1]_in[61] chanx[1][0]_out[41] sram[1932]->outb sram[1932]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[280], level=1, select_path_id=0. *****
*****1*****
Xsram[1932] sram->in sram[1932]->out sram[1932]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1932]->out) 0
.nodeset V(sram[1932]->outb) vsp
Xmux_1level_tapbuf_size2[281] grid[1][0]_pin[0][0][9] chany[1][1]_in[59] chanx[1][0]_out[43] sram[1933]->outb sram[1933]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[281], level=1, select_path_id=0. *****
*****1*****
Xsram[1933] sram->in sram[1933]->out sram[1933]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1933]->out) 0
.nodeset V(sram[1933]->outb) vsp
Xmux_1level_tapbuf_size2[282] grid[1][0]_pin[0][0][9] chany[1][1]_in[57] chanx[1][0]_out[45] sram[1934]->outb sram[1934]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[282], level=1, select_path_id=0. *****
*****1*****
Xsram[1934] sram->in sram[1934]->out sram[1934]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1934]->out) 0
.nodeset V(sram[1934]->outb) vsp
Xmux_1level_tapbuf_size2[283] grid[1][0]_pin[0][0][9] chany[1][1]_in[55] chanx[1][0]_out[47] sram[1935]->outb sram[1935]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[283], level=1, select_path_id=0. *****
*****1*****
Xsram[1935] sram->in sram[1935]->out sram[1935]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1935]->out) 0
.nodeset V(sram[1935]->outb) vsp
Xmux_1level_tapbuf_size2[284] grid[1][0]_pin[0][0][9] chany[1][1]_in[53] chanx[1][0]_out[49] sram[1936]->outb sram[1936]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[284], level=1, select_path_id=0. *****
*****1*****
Xsram[1936] sram->in sram[1936]->out sram[1936]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1936]->out) 0
.nodeset V(sram[1936]->outb) vsp
Xmux_1level_tapbuf_size2[285] grid[1][0]_pin[0][0][11] chany[1][1]_in[51] chanx[1][0]_out[51] sram[1937]->outb sram[1937]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[285], level=1, select_path_id=0. *****
*****1*****
Xsram[1937] sram->in sram[1937]->out sram[1937]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1937]->out) 0
.nodeset V(sram[1937]->outb) vsp
Xmux_1level_tapbuf_size2[286] grid[1][0]_pin[0][0][11] chany[1][1]_in[49] chanx[1][0]_out[53] sram[1938]->outb sram[1938]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[286], level=1, select_path_id=0. *****
*****1*****
Xsram[1938] sram->in sram[1938]->out sram[1938]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1938]->out) 0
.nodeset V(sram[1938]->outb) vsp
Xmux_1level_tapbuf_size2[287] grid[1][0]_pin[0][0][11] chany[1][1]_in[47] chanx[1][0]_out[55] sram[1939]->outb sram[1939]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[287], level=1, select_path_id=0. *****
*****1*****
Xsram[1939] sram->in sram[1939]->out sram[1939]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1939]->out) 0
.nodeset V(sram[1939]->outb) vsp
Xmux_1level_tapbuf_size2[288] grid[1][0]_pin[0][0][11] chany[1][1]_in[45] chanx[1][0]_out[57] sram[1940]->outb sram[1940]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[288], level=1, select_path_id=0. *****
*****1*****
Xsram[1940] sram->in sram[1940]->out sram[1940]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1940]->out) 0
.nodeset V(sram[1940]->outb) vsp
Xmux_1level_tapbuf_size2[289] grid[1][0]_pin[0][0][11] chany[1][1]_in[43] chanx[1][0]_out[59] sram[1941]->outb sram[1941]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[289], level=1, select_path_id=0. *****
*****1*****
Xsram[1941] sram->in sram[1941]->out sram[1941]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1941]->out) 0
.nodeset V(sram[1941]->outb) vsp
Xmux_1level_tapbuf_size2[290] grid[1][0]_pin[0][0][13] chany[1][1]_in[41] chanx[1][0]_out[61] sram[1942]->outb sram[1942]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[290], level=1, select_path_id=0. *****
*****1*****
Xsram[1942] sram->in sram[1942]->out sram[1942]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1942]->out) 0
.nodeset V(sram[1942]->outb) vsp
Xmux_1level_tapbuf_size2[291] grid[1][0]_pin[0][0][13] chany[1][1]_in[39] chanx[1][0]_out[63] sram[1943]->outb sram[1943]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[291], level=1, select_path_id=0. *****
*****1*****
Xsram[1943] sram->in sram[1943]->out sram[1943]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1943]->out) 0
.nodeset V(sram[1943]->outb) vsp
Xmux_1level_tapbuf_size2[292] grid[1][0]_pin[0][0][13] chany[1][1]_in[37] chanx[1][0]_out[65] sram[1944]->outb sram[1944]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[292], level=1, select_path_id=0. *****
*****1*****
Xsram[1944] sram->in sram[1944]->out sram[1944]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1944]->out) 0
.nodeset V(sram[1944]->outb) vsp
Xmux_1level_tapbuf_size2[293] grid[1][0]_pin[0][0][13] chany[1][1]_in[35] chanx[1][0]_out[67] sram[1945]->outb sram[1945]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[293], level=1, select_path_id=0. *****
*****1*****
Xsram[1945] sram->in sram[1945]->out sram[1945]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1945]->out) 0
.nodeset V(sram[1945]->outb) vsp
Xmux_1level_tapbuf_size2[294] grid[1][0]_pin[0][0][13] chany[1][1]_in[33] chanx[1][0]_out[69] sram[1946]->outb sram[1946]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[294], level=1, select_path_id=0. *****
*****1*****
Xsram[1946] sram->in sram[1946]->out sram[1946]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1946]->out) 0
.nodeset V(sram[1946]->outb) vsp
Xmux_1level_tapbuf_size2[295] grid[1][0]_pin[0][0][15] chany[1][1]_in[31] chanx[1][0]_out[71] sram[1947]->outb sram[1947]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[295], level=1, select_path_id=0. *****
*****1*****
Xsram[1947] sram->in sram[1947]->out sram[1947]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1947]->out) 0
.nodeset V(sram[1947]->outb) vsp
Xmux_1level_tapbuf_size2[296] grid[1][0]_pin[0][0][15] chany[1][1]_in[29] chanx[1][0]_out[73] sram[1948]->outb sram[1948]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[296], level=1, select_path_id=0. *****
*****1*****
Xsram[1948] sram->in sram[1948]->out sram[1948]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1948]->out) 0
.nodeset V(sram[1948]->outb) vsp
Xmux_1level_tapbuf_size2[297] grid[1][0]_pin[0][0][15] chany[1][1]_in[27] chanx[1][0]_out[75] sram[1949]->outb sram[1949]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[297], level=1, select_path_id=0. *****
*****1*****
Xsram[1949] sram->in sram[1949]->out sram[1949]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1949]->out) 0
.nodeset V(sram[1949]->outb) vsp
Xmux_1level_tapbuf_size2[298] grid[1][0]_pin[0][0][15] chany[1][1]_in[25] chanx[1][0]_out[77] sram[1950]->outb sram[1950]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[298], level=1, select_path_id=0. *****
*****1*****
Xsram[1950] sram->in sram[1950]->out sram[1950]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1950]->out) 0
.nodeset V(sram[1950]->outb) vsp
Xmux_1level_tapbuf_size2[299] grid[1][0]_pin[0][0][15] chany[1][1]_in[23] chanx[1][0]_out[79] sram[1951]->out sram[1951]->outb svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[299], level=1, select_path_id=1. *****
*****0*****
Xsram[1951] sram->in sram[1951]->out sram[1951]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1951]->out) 0
.nodeset V(sram[1951]->outb) vsp
Xmux_1level_tapbuf_size2[300] grid[1][1]_pin[0][2][42] chany[1][1]_in[21] chanx[1][0]_out[81] sram[1952]->outb sram[1952]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[300], level=1, select_path_id=0. *****
*****1*****
Xsram[1952] sram->in sram[1952]->out sram[1952]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1952]->out) 0
.nodeset V(sram[1952]->outb) vsp
Xmux_1level_tapbuf_size2[301] grid[1][1]_pin[0][2][42] chany[1][1]_in[19] chanx[1][0]_out[83] sram[1953]->outb sram[1953]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[301], level=1, select_path_id=0. *****
*****1*****
Xsram[1953] sram->in sram[1953]->out sram[1953]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1953]->out) 0
.nodeset V(sram[1953]->outb) vsp
Xmux_1level_tapbuf_size2[302] grid[1][1]_pin[0][2][42] chany[1][1]_in[17] chanx[1][0]_out[85] sram[1954]->outb sram[1954]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[302], level=1, select_path_id=0. *****
*****1*****
Xsram[1954] sram->in sram[1954]->out sram[1954]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1954]->out) 0
.nodeset V(sram[1954]->outb) vsp
Xmux_1level_tapbuf_size2[303] grid[1][1]_pin[0][2][42] chany[1][1]_in[15] chanx[1][0]_out[87] sram[1955]->outb sram[1955]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[303], level=1, select_path_id=0. *****
*****1*****
Xsram[1955] sram->in sram[1955]->out sram[1955]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1955]->out) 0
.nodeset V(sram[1955]->outb) vsp
Xmux_1level_tapbuf_size2[304] grid[1][1]_pin[0][2][42] chany[1][1]_in[13] chanx[1][0]_out[89] sram[1956]->outb sram[1956]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[304], level=1, select_path_id=0. *****
*****1*****
Xsram[1956] sram->in sram[1956]->out sram[1956]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1956]->out) 0
.nodeset V(sram[1956]->outb) vsp
Xmux_1level_tapbuf_size2[305] grid[1][1]_pin[0][2][46] chany[1][1]_in[11] chanx[1][0]_out[91] sram[1957]->outb sram[1957]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[305], level=1, select_path_id=0. *****
*****1*****
Xsram[1957] sram->in sram[1957]->out sram[1957]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1957]->out) 0
.nodeset V(sram[1957]->outb) vsp
Xmux_1level_tapbuf_size2[306] grid[1][1]_pin[0][2][46] chany[1][1]_in[9] chanx[1][0]_out[93] sram[1958]->outb sram[1958]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[306], level=1, select_path_id=0. *****
*****1*****
Xsram[1958] sram->in sram[1958]->out sram[1958]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1958]->out) 0
.nodeset V(sram[1958]->outb) vsp
Xmux_1level_tapbuf_size2[307] grid[1][1]_pin[0][2][46] chany[1][1]_in[7] chanx[1][0]_out[95] sram[1959]->outb sram[1959]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[307], level=1, select_path_id=0. *****
*****1*****
Xsram[1959] sram->in sram[1959]->out sram[1959]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1959]->out) 0
.nodeset V(sram[1959]->outb) vsp
Xmux_1level_tapbuf_size2[308] grid[1][1]_pin[0][2][46] chany[1][1]_in[5] chanx[1][0]_out[97] sram[1960]->outb sram[1960]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[308], level=1, select_path_id=0. *****
*****1*****
Xsram[1960] sram->in sram[1960]->out sram[1960]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1960]->out) 0
.nodeset V(sram[1960]->outb) vsp
Xmux_1level_tapbuf_size2[309] grid[1][1]_pin[0][2][46] chany[1][1]_in[3] chanx[1][0]_out[99] sram[1961]->outb sram[1961]->out svdd sgnd mux_1level_tapbuf_size2
***** SRAM bits for MUX[309], level=1, select_path_id=0. *****
*****1*****
Xsram[1961] sram->in sram[1961]->out sram[1961]->outb gvdd_sram_sbs sgnd  sram6T
.nodeset V(sram[1961]->out) 0
.nodeset V(sram[1961]->outb) vsp
.eom
