//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog netlist for pre-configured FPGA fabric by design: and2
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

//----- Default net type -----
`default_nettype none

module and2_top_formal_verification (
input [0:0] a,
input [0:0] b,
output [0:0] c);

// ----- Local wires for FPGA fabric -----
wire [0:63] gfpga_pad_GPIO_PAD_fm;
wire [0:0] ccff_head_fm;
wire [0:0] ccff_tail_fm;
wire [0:0] pReset_fm;
wire [0:0] prog_clk_fm;
wire [0:0] set_fm;
wire [0:0] reset_fm;
wire [0:0] clk_fm;

// ----- FPGA top-level module to be capsulated -----
	fpga_top U0_formal_verification (
		.pReset(pReset_fm[0]),
		.prog_clk(prog_clk_fm[0]),
		.set(set_fm[0]),
		.reset(reset_fm[0]),
		.clk(clk_fm[0]),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD_fm[0:63]),
		.ccff_head(ccff_head_fm[0]),
		.ccff_tail(ccff_tail_fm[0]));

// ----- Begin Connect Global ports of FPGA top module -----
	assign set_fm[0] = 1'b0;
	assign reset_fm[0] = 1'b0;
	assign clk_fm[0] = 1'b0;
	assign pReset_fm[0] = 1'b0;
	assign prog_clk_fm[0] = 1'b0;
// ----- End Connect Global ports of FPGA top module -----

// ----- Link BLIF Benchmark I/Os to FPGA I/Os -----
// ----- Blif Benchmark input a is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[22] -----
	assign gfpga_pad_GPIO_PAD_fm[22] = a[0];

// ----- Blif Benchmark input b is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[26] -----
	assign gfpga_pad_GPIO_PAD_fm[26] = b[0];

// ----- Blif Benchmark output c is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[9] -----
	assign c[0] = gfpga_pad_GPIO_PAD_fm[9];

// ----- Wire unused FPGA I/Os to constants -----
	assign gfpga_pad_GPIO_PAD_fm[0] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[1] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[2] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[3] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[4] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[5] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[6] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[7] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[8] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[10] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[11] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[12] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[13] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[14] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[15] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[16] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[17] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[18] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[19] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[20] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[21] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[23] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[24] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[25] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[27] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[28] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[29] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[30] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[31] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[32] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[33] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[34] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[35] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[36] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[37] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[38] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[39] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[40] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[41] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[42] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[43] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[44] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[45] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[46] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[47] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[48] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[49] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[50] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[51] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[52] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[53] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[54] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[55] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[56] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[57] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[58] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[59] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[60] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[61] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[62] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[63] = 1'b0;

// ----- Begin load bitstream to configuration memories -----
// ----- Begin assign bitstream to configuration memories -----
initial begin
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_out[0:16] = 17'b00000000110000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_DFFR_mem.mem_outb[0:16] = 17'b11111111001111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:9] = 10'b0000110000;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:9] = 10'b1111001111;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:9] = 10'b0100010000;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:9] = 10'b1011101111;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:9] = 10'b0000000001;
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:9] = 10'b1111111110;
	force U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.sb_0__0_.mem_top_track_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_0__1_.mem_top_track_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_0__1_.mem_top_track_8.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_0__1_.mem_top_track_8.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_0__1_.mem_top_track_16.mem_out[0:5] = 6'b001001;
	force U0_formal_verification.sb_0__1_.mem_top_track_16.mem_outb[0:5] = 6'b110110;
	force U0_formal_verification.sb_0__1_.mem_right_track_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_2.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__1_.mem_right_track_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__1_.mem_right_track_4.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__1_.mem_right_track_4.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__1_.mem_right_track_6.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_0__1_.mem_right_track_6.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_0__1_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_0__2_.mem_right_track_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__0_.mem_top_track_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__0_.mem_top_track_2.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__0_.mem_top_track_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__0_.mem_top_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_1__0_.mem_right_track_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__0_.mem_right_track_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_1__0_.mem_right_track_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__0_.mem_right_track_16.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_1__0_.mem_right_track_16.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__0_.mem_left_track_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_1__0_.mem_left_track_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__0_.mem_left_track_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_1__0_.mem_left_track_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__0_.mem_left_track_17.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_1__0_.mem_left_track_17.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__1_.mem_top_track_0.mem_out[0:7] = 8'b01000001;
	force U0_formal_verification.sb_1__1_.mem_top_track_0.mem_outb[0:7] = 8'b10111110;
	force U0_formal_verification.sb_1__1_.mem_top_track_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_1__1_.mem_top_track_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__1_.mem_top_track_16.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_1__1_.mem_top_track_16.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__1_.mem_right_track_0.mem_out[0:7] = 8'b01000100;
	force U0_formal_verification.sb_1__1_.mem_right_track_0.mem_outb[0:7] = 8'b10111011;
	force U0_formal_verification.sb_1__1_.mem_right_track_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_1__1_.mem_right_track_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__1_.mem_right_track_16.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_1__1_.mem_right_track_16.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_out[0:7] = 8'b01000001;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_outb[0:7] = 8'b10111110;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_17.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_17.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__1_.mem_left_track_1.mem_out[0:7] = 8'b01000001;
	force U0_formal_verification.sb_1__1_.mem_left_track_1.mem_outb[0:7] = 8'b10111110;
	force U0_formal_verification.sb_1__1_.mem_left_track_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_1__1_.mem_left_track_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__1_.mem_left_track_17.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_1__1_.mem_left_track_17.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__2_.mem_right_track_0.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_1__2_.mem_right_track_0.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__2_.mem_right_track_8.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_1__2_.mem_right_track_8.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__2_.mem_right_track_16.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__2_.mem_right_track_16.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_3.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_3.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_1__2_.mem_left_track_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__2_.mem_left_track_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_1__2_.mem_left_track_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_1__2_.mem_left_track_17.mem_out[0:5] = 6'b010001;
	force U0_formal_verification.sb_1__2_.mem_left_track_17.mem_outb[0:5] = 6'b101110;
	force U0_formal_verification.sb_2__0_.mem_top_track_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_12.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_12.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_0.mem_out[0:7] = 8'b00010100;
	force U0_formal_verification.sb_2__1_.mem_top_track_0.mem_outb[0:7] = 8'b11101011;
	force U0_formal_verification.sb_2__1_.mem_top_track_8.mem_out[0:7] = 8'b00011000;
	force U0_formal_verification.sb_2__1_.mem_top_track_8.mem_outb[0:7] = 8'b11100111;
	force U0_formal_verification.sb_2__1_.mem_top_track_16.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_2__1_.mem_top_track_16.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_9.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_9.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_17.mem_out[0:7] = 8'b00000001;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_17.mem_outb[0:7] = 8'b11111110;
	force U0_formal_verification.sb_2__1_.mem_left_track_1.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_2__1_.mem_left_track_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_2__1_.mem_left_track_3.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_2__1_.mem_left_track_3.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_2__1_.mem_left_track_5.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_2__1_.mem_left_track_5.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_2__1_.mem_left_track_7.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.sb_2__1_.mem_left_track_7.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.sb_2__1_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_3.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_3.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_1.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_2.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_3.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_3.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_4.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_4.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_5.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_5.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_6.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_6.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_7.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_7.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_3.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_3.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_4.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_4.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_5.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_5.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_6.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_6.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_7.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_7.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_1.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_2.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_3.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_3.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_4.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_4.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_5.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_5.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_6.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_6.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_7.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_7.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.mem_out[0:5] = 6'b010100;
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.mem_outb[0:5] = 6'b101011;
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_3.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_3.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_4.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_4.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_5.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_5.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_6.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_6.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_7.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_7.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_0__1_.mem_left_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_1.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_2.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_3.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_3.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_4.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_4.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_5.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_5.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_6.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_6.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_7.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_0__1_.mem_right_ipin_7.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_1.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_2.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_3.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_3.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_4.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_4.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_5.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_5.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_6.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_6.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_7.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_0__2_.mem_right_ipin_7.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_1__1_.mem_left_ipin_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_1__1_.mem_left_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_3.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_3.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_4.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_4.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_5.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_1__1_.mem_right_ipin_5.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_1__2_.mem_left_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_3.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_3.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_4.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_4.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_5.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_5.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_1.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_2.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_3.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_3.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_4.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_4.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_5.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_5.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_6.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_6.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_7.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_2__1_.mem_left_ipin_7.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__1_.mem_right_ipin_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_2__1_.mem_right_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__1_.mem_right_ipin_1.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_2__1_.mem_right_ipin_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__1_.mem_right_ipin_2.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_2__1_.mem_right_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__1_.mem_right_ipin_3.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_2__1_.mem_right_ipin_3.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__1_.mem_right_ipin_4.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_2__1_.mem_right_ipin_4.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__1_.mem_right_ipin_5.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_2__1_.mem_right_ipin_5.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_1.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_1.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_2.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_3.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_3.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_4.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_4.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_5.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_5.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_6.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_6.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_7.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_2__2_.mem_left_ipin_7.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_0.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_0.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_1.mem_out[0:5] = 6'b100100;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_1.mem_outb[0:5] = 6'b011011;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_2.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_2.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_3.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_3.mem_outb[0:5] = 6'b111110;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_4.mem_out[0:5] = 6'b001100;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_4.mem_outb[0:5] = 6'b110011;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_5.mem_out[0:5] = 6'b000001;
	force U0_formal_verification.cby_2__2_.mem_right_ipin_5.mem_outb[0:5] = 6'b111110;
end
// ----- End assign bitstream to configuration memories -----
// ----- End load bitstream to configuration memories -----
endmodule
// ----- END Verilog module for and2_top_formal_verification -----

//----- Default net type -----
`default_nettype none

