// Benchmark "TOP" written by ABC on Mon Feb  4 17:32:57 2019

module misex3 ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n,
    r2, s2, t2, u2, n2, o2, p2, q2, h2, i2, j2, k2, m2, l2  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n;
  output r2, s2, t2, u2, n2, o2, p2, q2, h2, i2, j2, k2, m2, l2;
  wire n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
    n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
    n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
    n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
    n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
    n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
    n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
    n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
    n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
    n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
    n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
    n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
    n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
    n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
    n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
    n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
    n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
    n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
    n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
    n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
    n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
    n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
    n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
    n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
    n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
    n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
    n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
    n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
    n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
    n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
    n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
    n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
    n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
    n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
    n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
    n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
    n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
    n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
    n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
    n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
    n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
    n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
    n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
    n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
    n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
    n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
    n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
    n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
    n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
    n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
    n758, n759, n760, n761, n762;
  assign r2 = ~n293;
  assign s2 = ~n74;
  assign t2 = ~n217;
  assign u2 = ~n148;
  assign n2 = ~n68;
  assign o2 = ~n62;
  assign p2 = ~n388;
  assign q2 = ~n349;
  assign h2 = ~n56;
  assign i2 = ~n569;
  assign j2 = ~n55;
  assign k2 = ~n50;
  assign m2 = ~n456;
  assign l2 = ~n757 | ~n759 | n46 | ~n747 | n44 | n45 | n42 | n43;
  assign n42 = f & (~n680 | ~n739 | ~n740);
  assign n43 = ~f & (n475 | n476 | ~n735);
  assign n44 = ~n & (~n722 | ~n724 | ~n728);
  assign n45 = n & (~n518 | ~n730 | ~n731);
  assign n46 = n548 | ~n744 | n544 | n547 | n542 | ~n543 | ~n540 | n541;
  assign n47 = n675 | n676 | n372 | i | l;
  assign n48 = n438 | n549 | n189;
  assign n49 = n434 & n662 & n661 & n51 & n437 & n439;
  assign n50 = n49 & n47 & n48;
  assign n51 = n657 & n573 & n656 & n431 & n425 & n428;
  assign n52 = n443 & n442 & n440 & n441;
  assign n53 = n675 | n189 | n438;
  assign n54 = n179 | n480 | n550 | n551;
  assign n55 = n54 & n53 & n51 & n52;
  assign n56 = n579 & n578 & n577 & n576 & n575 & n574 & n572 & n573;
  assign n57 = (n95 | n408) & (n409 | n88);
  assign n58 = n96 | n121;
  assign n59 = n648 & ~n404 & n361 & n402;
  assign n60 = n83 | n317;
  assign n61 = (n362 | n300) & (n363 | n426);
  assign n62 = ~n416 & ~n415 & ~n414 & n61 & n60 & n59 & n57 & n58;
  assign n63 = j | n243 | n119 | n591;
  assign n64 = (n177 | n362) & (n684 | n409);
  assign n65 = ~n297 & (n95 | n253 | n298);
  assign n66 = n620 & n619 & n572 & n618 & n617 & n69 & n574 & n211;
  assign n67 = ~n422 & (n591 | (n710 & n711));
  assign n68 = ~n420 & ~n419 & n67 & n66 & n65 & n64 & n59 & n63;
  assign n69 = n92 | n407 | n91;
  assign n70 = n595 | n92;
  assign n71 = n264 | ~d | n248;
  assign n72 = n701 & (n236 | n79);
  assign n73 = n232 & (n152 | n632);
  assign n74 = ~n267 & ~n266 & ~n265 & n73 & n72 & n71 & n69 & n70;
  assign n75 = ~h | ~k;
  assign n76 = n75 | l;
  assign n77 = n623 | ~n658;
  assign n78 = ~n167 & (n77 | ~n586);
  assign n79 = ~c | n459;
  assign n80 = e | n521;
  assign n81 = n612 & n302;
  assign n82 = n81 & n79 & n80;
  assign n83 = ~k | n199;
  assign n84 = m | j | ~l;
  assign n85 = n83 & (~n | n84);
  assign n86 = n684 | n83;
  assign n87 = (n192 | n605) & (n206 | n604);
  assign n88 = ~g | n603;
  assign n89 = n86 & n87 & (n85 | n88);
  assign n90 = (n110 | n156) & (n113 | n275);
  assign n91 = ~i | n538;
  assign n92 = ~a | n521;
  assign n93 = n90 & (n91 | n92);
  assign n94 = ~g | n600;
  assign n95 = n285 & n397;
  assign n96 = ~k | n167;
  assign n97 = n96 | n94 | n95;
  assign n98 = n601 | n199;
  assign n99 = ~i | n368;
  assign n100 = n98 & (~n | n99);
  assign n101 = ~h | n538;
  assign n102 = ~n | n129;
  assign n103 = h | n538;
  assign n104 = (n100 | n103) & (n101 | n102);
  assign n105 = ~g | n249;
  assign n106 = h | n197;
  assign n107 = (n100 | n106) & (n102 | n105);
  assign n108 = ~k | n179;
  assign n109 = n108 & (n | n84);
  assign n110 = n608 & n287 & n607;
  assign n111 = (n101 | n92) & (n110 | n105);
  assign n112 = n135 | n119;
  assign n113 = n218 & n295;
  assign n114 = ~g | n393;
  assign n115 = n112 & n111 & (n113 | n114);
  assign n116 = (n110 | n164) & (n113 | n189);
  assign n117 = e | n609;
  assign n118 = n116 & (n92 | n117);
  assign n119 = ~a | n271;
  assign n120 = ~e | n609;
  assign n121 = n118 & (n119 | n120);
  assign n122 = (n110 | n106) & (n113 | n202);
  assign n123 = n122 & (n92 | n103);
  assign n124 = n153 | n399;
  assign n125 = ~n610 | ~g | n237;
  assign n126 = j | n154;
  assign n127 = ~i | n609;
  assign n128 = n124 & n125 & (n126 | n127);
  assign n129 = n401 & n512 & n527 & n760;
  assign n130 = (n106 | n99) & (n129 | n105);
  assign n131 = n519 | ~i | n121;
  assign n132 = (n123 | n588) & (n95 | n128);
  assign n133 = ~e | n271;
  assign n134 = n131 & n132 & (n130 | n133);
  assign n135 = ~h | n243;
  assign n136 = h | n243;
  assign n137 = (n100 | n136) & (n135 | n102);
  assign n138 = ~n137 & (~n625 | (b & ~n479));
  assign n139 = ~n89 & (~n325 | ~n606);
  assign n140 = ~n167 & (~n683 | (~n121 & ~n601));
  assign n141 = ~n95 & (~n687 | (~n96 & ~n127));
  assign n142 = n133 | n601 | n179 | n106;
  assign n143 = n590 | n591;
  assign n144 = n136 | n587 | n588;
  assign n145 = ~n139 & ~n140 & (n | n134);
  assign n146 = (n93 | n591) & (n104 | n616);
  assign n147 = n688 & (n107 | n269);
  assign n148 = n147 & n146 & n145 & n144 & n143 & n142 & n66 & ~n138;
  assign n149 = n689 | n108;
  assign n150 = (n372 | n193) & (n613 | n624);
  assign n151 = ~f | n603;
  assign n152 = n149 & n150 & (n109 | n151);
  assign n153 = ~m | n611;
  assign n154 = ~l | ~m;
  assign n155 = n153 & (i | n154);
  assign n156 = ~i | n197;
  assign n157 = j | n197;
  assign n158 = n156 & n157;
  assign n159 = (n155 | n105) & (n158 | n589);
  assign n160 = n690 & (n164 | n126);
  assign n161 = n644 & n647;
  assign n162 = i | n197;
  assign n163 = n159 & n160 & (n161 | n162);
  assign n164 = g | n249;
  assign n165 = (n164 | n96) & (n | n163);
  assign n166 = n75 | ~m | n;
  assign n167 = ~m | n;
  assign n168 = ~l | ~h | j;
  assign n169 = n166 & (n167 | n168);
  assign n170 = ~f | n243;
  assign n171 = ~e | n196;
  assign n172 = (n169 | n171) & (~n78 | n170);
  assign n173 = n196 | d | n169;
  assign n174 = d | n197;
  assign n175 = n173 & (~n78 | n174);
  assign n176 = j | n75;
  assign n177 = n176 & (i | n75);
  assign n178 = n299 & n300 & n76 & n177;
  assign n179 = m | n;
  assign n180 = j | n603;
  assign n181 = ~l | n179;
  assign n182 = (n180 | n181) & (n178 | n179);
  assign n183 = ~e | n615;
  assign n184 = ~n | n183;
  assign n185 = (n99 | n184) & (n98 | n183);
  assign n186 = ~n184 & ~n761 & (~n114 | ~n189);
  assign n187 = ~n186 & (n185 | (n202 & n676));
  assign n188 = n183 | n391;
  assign n189 = g | n393;
  assign n190 = n187 & (n188 | (n114 & n189));
  assign n191 = (n206 | n624) & (n689 | n83);
  assign n192 = k | n199;
  assign n193 = ~j | n249;
  assign n194 = n191 & (n192 | n193);
  assign n195 = n194 & (n85 | n151);
  assign n196 = ~f | g;
  assign n197 = ~f | ~g;
  assign n198 = (n169 | n196) & (~n78 | n197);
  assign n199 = m | ~n;
  assign n200 = ~l | n199;
  assign n201 = (n180 | n200) & (n178 | n199);
  assign n202 = h | n570;
  assign n203 = (n100 | n202) & (n102 | n114);
  assign n204 = n203 & (n201 | (n170 & n171));
  assign n205 = n691 & n692 & (n85 | n314);
  assign n206 = l | n199;
  assign n207 = ~k | n393;
  assign n208 = n89 & n205 & (n206 | n207);
  assign n209 = ~n152 & (~n133 | ~n430);
  assign n210 = n595 | n599;
  assign n211 = n595 | n353;
  assign n212 = n693 & (~e | n195 | n324);
  assign n213 = ~n209 & (n285 | (n165 & n595));
  assign n214 = n208 | n315;
  assign n215 = (n172 | n119) & (n175 | n287);
  assign n216 = n694 & (n182 | n302);
  assign n217 = n216 & n190 & n215 & n214 & n213 & n212 & n210 & n211;
  assign n218 = ~a | n560;
  assign n219 = n167 | n218;
  assign n220 = (n168 | n219) & (n218 | n166);
  assign n221 = ~n658 | ~n586 | n623;
  assign n222 = ~f & ~n538;
  assign n223 = ~n219 & n221 & (n222 | ~n261);
  assign n224 = e | n488;
  assign n225 = e | n196;
  assign n226 = ~n223 & (n220 | (n224 & n225));
  assign n227 = n393 | ~j | n372;
  assign n228 = (n613 | n207) & (n109 | n314);
  assign n229 = n640 & n643;
  assign n230 = n227 & n228 & (n229 | n108);
  assign n231 = ~e | n626;
  assign n232 = n190 & n226 & (n230 | n231);
  assign n233 = ~n83 & (~n252 | ~n639);
  assign n234 = (n192 | n322) & (n256 | n206);
  assign n235 = g | n603;
  assign n236 = ~n233 & n234 & (n85 | n235);
  assign n237 = k | n154;
  assign n238 = (i | n161) & (~j | n237);
  assign n239 = ~n591 & (~n91 | (~j & ~n538));
  assign n240 = ~n239 & (n | (n699 & n700));
  assign n241 = n165 & n240 & (n96 | n117);
  assign n242 = ~i | n243;
  assign n243 = ~e | ~g;
  assign n244 = n242 & (j | n243);
  assign n245 = n96 | n120;
  assign n246 = n697 & (n120 | n126);
  assign n247 = n696 & n695 & (n244 | n589);
  assign n248 = n245 & (n | (n246 & n247));
  assign n249 = ~f | ~h;
  assign n250 = n249 | n102 | e;
  assign n251 = n629 & n88;
  assign n252 = j | n609;
  assign n253 = i | n602;
  assign n254 = ~g | n360;
  assign n255 = n254 & n253 & n251 & n252;
  assign n256 = g | n75;
  assign n257 = n698 & (n376 | (n628 & n649));
  assign n258 = (n94 | n96) & (n629 | n630);
  assign n259 = ~l | n167;
  assign n260 = n257 & n258 & (n255 | n259);
  assign n261 = ~f | n538;
  assign n262 = (n169 | n225) & (~n78 | n261);
  assign n263 = ~n260 & (~n655 | (d & ~n524));
  assign n264 = a | ~b;
  assign n265 = ~n201 & (~n325 | (~n261 & ~n616));
  assign n266 = ~n352 & (~n262 | n263);
  assign n267 = ~n526 & (~n250 | (~n100 & ~n631));
  assign n268 = n344 & (n83 | n633);
  assign n269 = ~b | n598;
  assign n270 = n268 & (n194 | n269);
  assign n271 = ~c | d;
  assign n272 = n79 & (~f | n271);
  assign n273 = (n100 | n634) & (n164 | n102);
  assign n274 = n273 & n107;
  assign n275 = ~i | n570;
  assign n276 = j | n570;
  assign n277 = n275 & n276;
  assign n278 = (n155 | n114) & (n277 | n589);
  assign n279 = n749 & (n189 | n126);
  assign n280 = i | n570;
  assign n281 = n278 & n279 & (n161 | n280);
  assign n282 = (n96 | n189) & (n | n281);
  assign n283 = n286 | g | n169;
  assign n284 = n283 & (d | ~n78 | n243);
  assign n285 = ~e | n264;
  assign n286 = d | ~e;
  assign n287 = c | ~a | ~b;
  assign n288 = n285 & (n286 | n287);
  assign n289 = (n236 | n635) & (n104 | n616);
  assign n290 = (n260 | n288) & (n284 | ~n545);
  assign n291 = n107 | n315;
  assign n292 = (n182 | n272) & (n274 | n625);
  assign n293 = n292 & n291 & n290 & n289 & n270 & n232;
  assign n294 = n123 & (n119 | n136);
  assign n295 = n596 & n594;
  assign n296 = n112 & n111 & (n295 | n114);
  assign n297 = ~n636 & (~n355 | (~n167 & ~n296));
  assign n298 = n | n126;
  assign n299 = ~h | n360;
  assign n300 = ~k | n603;
  assign n301 = n180 & n300 & n299 & n176;
  assign n302 = ~c | n524;
  assign n303 = n302 & (~c | n196);
  assign n304 = (n113 | n646) & (~j | n645);
  assign n305 = ~j | n197;
  assign n306 = n304 & (n110 | n305);
  assign n307 = n121 & (n95 | n94);
  assign n308 = ~n95 & ~n644 & (~n88 | ~n660);
  assign n309 = ~n308 & (n329 | n339 | n435);
  assign n310 = (n118 | n126) & (n306 | n237);
  assign n311 = ~l | n519;
  assign n312 = n309 & n310 & (n307 | n311);
  assign n313 = n183 & n390;
  assign n314 = f | n603;
  assign n315 = ~b | n286;
  assign n316 = (n314 | n315) & (n313 | n235);
  assign n317 = n633 & n316;
  assign n318 = (n80 & (~n | n371)) | (n & n371);
  assign n319 = (n88 | n318) & (~n | n317);
  assign n320 = n393 | ~j | n315;
  assign n321 = n269 | n193;
  assign n322 = ~j | n609;
  assign n323 = n320 & n321 & (n313 | n322);
  assign n324 = b | ~c;
  assign n325 = ~f | n324;
  assign n326 = (n315 | n643) & (n313 | n252);
  assign n327 = j | n249;
  assign n328 = n326 & (n269 | n327);
  assign n329 = ~h | n621;
  assign n330 = n328 & (n325 | n329);
  assign n331 = (n316 | n84) & (n330 | n435);
  assign n332 = m | k | ~l;
  assign n333 = n331 & (n323 | n332);
  assign n334 = (n315 | n640) & (n313 | n639);
  assign n335 = i | n249;
  assign n336 = n334 & (n269 | n335);
  assign n337 = ~n199 & (~n336 | (~n253 & ~n371));
  assign n338 = ~n337 & (n80 | n179 | n253);
  assign n339 = n303 & n637;
  assign n340 = (n339 | n181) & (n325 | n200);
  assign n341 = ~n318 & (~n704 | (~n332 & ~n605));
  assign n342 = n243 | n490 | ~j | n119;
  assign n343 = n298 | n119 | n120;
  assign n344 = n633 | ~n | n84;
  assign n345 = n705 & (n301 | n340);
  assign n346 = n65 & (n319 | n435);
  assign n347 = (n312 & (~n | n333)) | (n & n333);
  assign n348 = (n682 | n641) & (n338 | n433);
  assign n349 = n348 & n347 & n346 & n345 & n344 & n343 & ~n341 & n342;
  assign n350 = (n113 | n280) & (i | n645);
  assign n351 = n350 & (n110 | n162);
  assign n352 = ~a | n324;
  assign n353 = ~b | n597;
  assign n354 = n353 & n287 & n352;
  assign n355 = n114 | n219;
  assign n356 = (n599 | n105) & (n295 | n114);
  assign n357 = n112 & (n92 | (n105 & n101));
  assign n358 = n355 & (n167 | (n356 & n357));
  assign n359 = n707 & (n285 | n630 | n605);
  assign n360 = ~j | k;
  assign n361 = n359 & (n358 | n360);
  assign n362 = (n339 | n179) & (n325 | n199);
  assign n363 = (n339 | n108) & (n325 | n83);
  assign n364 = ~n88 & (~n706 | (~n167 & ~n433));
  assign n365 = ~n364 & (n629 | (n259 & n630));
  assign n366 = n365 & (n96 | n322);
  assign n367 = n519 | n | n121;
  assign n368 = ~k | m;
  assign n369 = (n253 | n318) & (~n | n336);
  assign n370 = n367 & (n368 | (n369 & n319));
  assign n371 = n395 & n315 & n606;
  assign n372 = k | n179;
  assign n373 = (n372 | n80) & (n371 | n192);
  assign n374 = ~i | k | ~l | n167;
  assign n375 = ~k | ~n610;
  assign n376 = l | n167;
  assign n377 = n374 & (n375 | (n376 & n259));
  assign n378 = ~j | n603;
  assign n379 = n378 & n329;
  assign n380 = n644 | n587 | n627;
  assign n381 = n647 | n587 | n627;
  assign n382 = n351 | n | n161;
  assign n383 = (n294 | n377) & (n363 | n379);
  assign n384 = n373 | n605;
  assign n385 = (n95 | n366) & (~j | n370);
  assign n386 = n362 | n299;
  assign n387 = n361 & (n323 | n192);
  assign n388 = n387 & n386 & n385 & n384 & n383 & n382 & n380 & n381;
  assign n389 = ~n372 & (~n303 | ~n637);
  assign n390 = n635 & n638;
  assign n391 = ~n | n401;
  assign n392 = n188 & (n390 | n391);
  assign n393 = f | ~h;
  assign n394 = (n393 | n315) & (n249 | n269);
  assign n395 = n616 & n625;
  assign n396 = e | n324;
  assign n397 = ~b | n524;
  assign n398 = n397 & n396 & n395 & n315;
  assign n399 = ~i | n602;
  assign n400 = (n398 | n399) & (~i | n394);
  assign n401 = m | n360;
  assign n402 = n399 | n | n80 | n401;
  assign n403 = h & n610;
  assign n404 = n403 & (n389 | (~n192 & ~n325));
  assign n405 = n253 | n641;
  assign n406 = (n256 | n167) & (n376 | n176);
  assign n407 = n | n592;
  assign n408 = n405 & n406 & (n407 | n399);
  assign n409 = (n108 | n80) & (n371 | n83);
  assign n410 = i & ~n394;
  assign n411 = n & (n410 | (~n127 & ~n313));
  assign n412 = j | i;
  assign n413 = n412 | ~k | n259;
  assign n414 = ~n115 & (~n413 | (n77 & ~n167));
  assign n415 = ~n527 & (n411 | (~n318 & ~n399));
  assign n416 = ~n591 & (~n709 | (~n110 & ~n327));
  assign n417 = ~n433 & (~n351 | (~n119 & ~n627));
  assign n418 = ~n311 & ~n & ~n251;
  assign n419 = ~n95 & (n418 | (~n376 & ~n649));
  assign n420 = ~n83 & (~n328 | ~n336);
  assign n421 = i & k;
  assign n422 = ~n167 & (n417 | (~n294 & n421));
  assign n423 = n654 | ~f | n598;
  assign n424 = j | k;
  assign n425 = n259 | n399 | n423 | n424;
  assign n426 = ~h | n600;
  assign n427 = n651 | ~n | n557;
  assign n428 = n427 | n426 | n332;
  assign n429 = n650 | n114 | n181;
  assign n430 = ~e | n521;
  assign n431 = n429 | n430;
  assign n432 = ~n545 | n655;
  assign n433 = ~l | ~j | ~k;
  assign n434 = n399 | n167 | n432 | n433;
  assign n435 = ~l | n368;
  assign n436 = n170 | n526;
  assign n437 = n436 | ~n403 | n435;
  assign n438 = n181 | n375;
  assign n439 = n438 | n231 | n105;
  assign n440 = n652 | n202 | n632;
  assign n441 = ~n653 | n435 | n445;
  assign n442 = n181 | n202 | n430 | ~n473;
  assign n443 = n712 & (n332 | n427 | n378);
  assign n444 = n106 | n613 | n231 | n658;
  assign n445 = h | n621;
  assign n446 = m | k | l;
  assign n447 = n444 & (n436 | n445 | n446);
  assign n448 = n551 | n | n446;
  assign n449 = n448 & (n179 | n127 | n433);
  assign n450 = k | n189 | n181 | n632;
  assign n451 = n332 | n651 | ~h | n224;
  assign n452 = n450 & n451;
  assign n453 = n641 | n654 | n660 | n477;
  assign n454 = n105 | n181 | n549 | n650;
  assign n455 = (n449 | n480) & (n452 | n412);
  assign n456 = n455 & n454 & n453 & n49 & n52 & n447;
  assign n457 = i | n179;
  assign n458 = (~k | n457) & (n179 | ~n412);
  assign n459 = e | ~f;
  assign n460 = a | n526;
  assign n461 = j & ~n630 & (n459 | n460);
  assign n462 = ~n758 & (~h | n438 | ~n479);
  assign n463 = f | ~c | e;
  assign n464 = ~n461 & n462 & (n458 | n463);
  assign n465 = b | n199;
  assign n466 = n200 & n83 & n465 & n298;
  assign n467 = (b | n200) & (c | n181);
  assign n468 = ~n167 & (~n737 | (~b & ~n479));
  assign n469 = h | j | n199;
  assign n470 = (j | n83) & (~i | n663);
  assign n471 = ~j | n199;
  assign n472 = n469 & n470 & (~h | n471);
  assign n473 = ~k & n610;
  assign n474 = n473 & b & ~n199;
  assign n475 = ~h & (n474 | (~i & ~n206));
  assign n476 = ~n673 & (~n521 | (~e & n324));
  assign n477 = f | n659;
  assign n478 = n477 & (f | a | e);
  assign n479 = c | d;
  assign n480 = f | n479;
  assign n481 = n669 | c | e;
  assign n482 = b | e | ~n | n669;
  assign n483 = n375 | ~n615 | ~h | n259;
  assign n484 = (d | n734) & (n457 | n480);
  assign n485 = n199 | n675;
  assign n486 = ~n762 & n485 & n484 & n483 & n481 & n482;
  assign n487 = c & ~n655;
  assign n488 = f | g;
  assign n489 = b | n488;
  assign n490 = n | n237;
  assign n491 = (j | n490) & (n199 | ~n626);
  assign n492 = ~n199 & (~n741 | (~j & ~n525));
  assign n493 = n742 & (n670 | n671);
  assign n494 = ~n492 & ~n756 & (i | n491);
  assign n495 = n493 & n494 & (n457 | n271);
  assign n496 = c | n488;
  assign n497 = n664 & n463;
  assign n498 = (n106 | n231) & (~j | n497);
  assign n499 = (n716 | n167) & (n498 | n179);
  assign n500 = n496 | n372;
  assign n501 = (n527 | n671) & (n719 | n613);
  assign n502 = n718 & (n436 | (n206 & n192));
  assign n503 = n502 & n501 & n499 & n500;
  assign n504 = ~j & ~n372 & (~n271 | ~n302);
  assign n505 = (b | n199) & (c | n179);
  assign n506 = ~b | ~e | ~n | n666;
  assign n507 = e | n505 | n650;
  assign n508 = (n525 | n471) & (n457 | n479);
  assign n509 = n478 | n167;
  assign n510 = ~n626 | j | n192;
  assign n511 = n510 & n509 & n508 & n507 & ~n504 & n506;
  assign n512 = i | n368;
  assign n513 = m | n603;
  assign n514 = i | m;
  assign n515 = n512 & n513 & (~l | n514);
  assign n516 = n253 & n127;
  assign n517 = (n426 | n446) & (n516 | n666);
  assign n518 = n517 & (n401 | n151);
  assign n519 = ~k | ~m;
  assign n520 = n519 & (j | ~m);
  assign n521 = c | ~d;
  assign n522 = n81 & (g | n521);
  assign n523 = ~n311 & n403 & (~n174 | ~n261);
  assign n524 = ~e | f;
  assign n525 = b | n524;
  assign n526 = ~d | n615;
  assign n527 = j | n368;
  assign n528 = n99 & n527;
  assign n529 = n717 & (h | n524 | n636);
  assign n530 = (n521 | n525) & (~j | n716);
  assign n531 = (i | n432) & (n254 | n665);
  assign n532 = n634 & n550 & (n135 | n650);
  assign n533 = n532 & n531 & n529 & n530;
  assign n534 = ~c & ~n524;
  assign n535 = (~n180 | ~n628) & (~n463 | n534);
  assign n536 = ~j & (~n660 | (~n156 & ~n231));
  assign n537 = n396 & (a | c | e);
  assign n538 = e | ~g;
  assign n539 = ~n162 & (~n108 | ~n181);
  assign n540 = n375 | n259 | n114;
  assign n541 = ~n489 & (~n206 | ~n663);
  assign n542 = ~n613 & (~n497 | (~c & ~n660));
  assign n543 = n438 | n101;
  assign n544 = ~n231 & (n539 | (~n156 & ~n613));
  assign n545 = a & ~n615;
  assign n546 = n545 & ~n655 & (~n630 | ~n672);
  assign n547 = ~n457 & (~n631 | (~n105 & ~n231));
  assign n548 = ~n179 & (n535 | n536 | ~n715);
  assign n549 = ~e | n479;
  assign n550 = l | n424;
  assign n551 = i | g | h;
  assign n552 = n112 | n155 | n;
  assign n553 = n119 | n245;
  assign n554 = f | n167;
  assign n555 = (n168 | n554) & (f | n166);
  assign n556 = n555 | ~e | g;
  assign n557 = f | n243;
  assign n558 = n556 & (~n78 | n557);
  assign n559 = ~n99 & ~g & n;
  assign n560 = ~b | ~d;
  assign n561 = (n203 | n560) & (n526 | ~n748);
  assign n562 = (n175 | n287) & (n282 | n594);
  assign n563 = n236 | n638;
  assign n564 = (n352 | n558) & (~e | n561);
  assign n565 = n608 | n172;
  assign n566 = n677 & n553 & n552 & n342 & n143 & n63;
  assign n567 = n226 & n270 & (n89 | n625);
  assign n568 = n750 & n752 & n656 & n661 & n441 & n657 & n440 & n662;
  assign n569 = n568 & n567 & n447 & n566 & n565 & n564 & n562 & n563;
  assign n570 = f | ~g;
  assign n571 = (g | n555) & (~n78 | n570);
  assign n572 = n595 | n352;
  assign n573 = n652 | n106 | n549;
  assign n574 = n593 | n596;
  assign n575 = n626 | ~a | n262;
  assign n576 = n571 | ~d | ~n545;
  assign n577 = n753 & (n654 | (n175 & n248));
  assign n578 = n282 | n596;
  assign n579 = n566 & (n165 | n352);
  assign n580 = l | ~n421;
  assign n581 = ~l | ~h | i;
  assign n582 = (~l & n622) | (n603 & (l | n622));
  assign n583 = ~h | n611;
  assign n584 = ~l | n360;
  assign n585 = ~l | n621;
  assign n586 = n585 & n584 & n583 & n582 & n580 & n581;
  assign n587 = n | n119;
  assign n588 = ~i | n154;
  assign n589 = l | n519;
  assign n590 = n119 | n242;
  assign n591 = n | n589;
  assign n592 = j | n519;
  assign n593 = n407 | n275;
  assign n594 = ~a | n286;
  assign n595 = n156 | n407;
  assign n596 = ~e | ~a | ~c;
  assign n597 = d | a;
  assign n598 = ~d | e;
  assign n599 = ~a | n598;
  assign n600 = ~i | j;
  assign n601 = ~l | n600;
  assign n602 = ~g | ~h;
  assign n603 = h | ~i;
  assign n604 = ~g | n75;
  assign n605 = ~j | n602;
  assign n606 = n396 & n397;
  assign n607 = n599 & n353;
  assign n608 = n92 & n352;
  assign n609 = g | ~h;
  assign n610 = i & j;
  assign n611 = ~j | l;
  assign n612 = ~f | n521;
  assign n613 = l | n179;
  assign n614 = ~g | ~n421;
  assign n615 = ~b | ~c;
  assign n616 = d | n615;
  assign n617 = n590 | n407;
  assign n618 = n593 | n594;
  assign n619 = n97 & n70 & n210;
  assign n620 = (n595 | n287) & (n593 | n218);
  assign n621 = i | ~j;
  assign n622 = j | ~k;
  assign n623 = k & ~n600;
  assign n624 = ~k | n249;
  assign n625 = ~b | n521;
  assign n626 = ~c | ~d;
  assign n627 = i | n243;
  assign n628 = n614 & n605;
  assign n629 = ~g | n621;
  assign n630 = k | n167;
  assign n631 = h | n459;
  assign n632 = e | n626;
  assign n633 = n269 | n151;
  assign n634 = h | n196;
  assign n635 = ~b | n459;
  assign n636 = ~l | n412;
  assign n637 = n612 & n272;
  assign n638 = ~f | n560;
  assign n639 = i | n609;
  assign n640 = i | n393;
  assign n641 = n622 | ~l | n167;
  assign n642 = j | n602;
  assign n643 = j | n393;
  assign n644 = ~j | n154;
  assign n645 = n538 | n92;
  assign n646 = ~j | n570;
  assign n647 = ~m | n360;
  assign n648 = (n392 | n127) & (n400 | n391);
  assign n649 = ~g | n622;
  assign n650 = k | n600;
  assign n651 = b | n626;
  assign n652 = n621 | ~k | n181;
  assign n653 = n222 & ~n526;
  assign n654 = a | n615;
  assign n655 = ~f | ~d | ~e;
  assign n656 = ~n653 | n332 | n426;
  assign n657 = n632 | n429;
  assign n658 = k | n621;
  assign n659 = d | e;
  assign n660 = i | ~g | h;
  assign n661 = n445 | n435 | n427;
  assign n662 = n430 | n202 | n652;
  assign n663 = n83 & n471;
  assign n664 = ~g | n479;
  assign n665 = a | n598;
  assign n666 = m | n424;
  assign n667 = ~h | n514;
  assign n668 = k | n514;
  assign n669 = h | n514;
  assign n670 = m | n600;
  assign n671 = n | n479;
  assign n672 = h | n167;
  assign n673 = g | n199;
  assign n674 = h & ~n650;
  assign n675 = e | n479;
  assign n676 = h | n488;
  assign n677 = n343 & n144 & n454 & n617 & n381 & n380;
  assign n678 = (e & ~n119) | (~n92 & (~e | ~n119));
  assign n679 = (n479 & n674) | (~g & (~n479 | n674));
  assign n680 = n755 & (i | n466 | h);
  assign n681 = ~n610 | l | n115;
  assign n682 = n590 & n93;
  assign n683 = n681 & (n682 | n584);
  assign n684 = n642 & n253;
  assign n685 = (n684 | n108) & (n109 | n88);
  assign n686 = (n605 | n372) & (n604 | n613);
  assign n687 = (n614 | n376) & (n88 | n259);
  assign n688 = ~n141 & (n82 | (n685 & n686));
  assign n689 = n335 & n327;
  assign n690 = (n588 | n106) & (n237 | n305);
  assign n691 = n229 | n83;
  assign n692 = n393 | ~j | n192;
  assign n693 = ~a | b | ~d | n198;
  assign n694 = (n607 | n165) & (n204 | n625);
  assign n695 = (n161 | n627) & (n155 | n135);
  assign n696 = n243 | ~j | n237;
  assign n697 = (n588 | n136) & (n242 | n592);
  assign n698 = n256 | n167;
  assign n699 = (n155 | n101) & (n238 | n538);
  assign n700 = (n588 | n103) & (n117 | n126);
  assign n701 = (n182 | n612) & (n241 | n92);
  assign n702 = ~n294 & (~n585 | (l & n610));
  assign n703 = ~n95 & (~n252 | ~n254 | ~n256);
  assign n704 = (n84 | n88) & (n642 | n435);
  assign n705 = (n167 | ~n702) & (n259 | ~n703);
  assign n706 = n490 & (n96 | n611);
  assign n707 = n354 | n360 | n167 | n105;
  assign n708 = ~h | j;
  assign n709 = (n113 | n643) & (~n678 | n708);
  assign n710 = (n95 | n88) & (j | n645);
  assign n711 = (n110 | n157) & (n113 | n276);
  assign n712 = n167 | n127 | n584 | n423;
  assign n713 = (d | n525) & (j | n436);
  assign n714 = (b | c) & (n127 | n433);
  assign n715 = (n253 | n463) & (n103 | ~n473);
  assign n716 = n676 & n478;
  assign n717 = a | b;
  assign n718 = n433 | n487 | ~h | n199;
  assign n719 = n496 & ~n534;
  assign n720 = n478 & n665 & n432;
  assign n721 = ~n523 & (g | n520 | n720);
  assign n722 = n721 & (n670 | (n496 & n480));
  assign n723 = (n522 | n669) & (n164 | n666);
  assign n724 = n723 & (n668 | (n202 & n664));
  assign n725 = n231 | n156 | n401;
  assign n726 = n592 | n432;
  assign n727 = n725 & n726 & (n719 | n667);
  assign n728 = n518 & n727 & (n496 | n515);
  assign n729 = (n436 | n667) & (n525 | n528);
  assign n730 = n729 & (n515 | n436);
  assign n731 = (n669 | n397) & (n525 | n668);
  assign n732 = n526 | e | n472;
  assign n733 = n672 | ~n597 | n636;
  assign n734 = n754 & (~h | n438);
  assign n735 = n732 & n733 & (~c | n734);
  assign n736 = n | a | ~g;
  assign n737 = (i | n665) & (~n545 | n659);
  assign n738 = ~n468 & (n311 | ~n403 | n736);
  assign n739 = n738 & (n665 | (n672 & n96));
  assign n740 = (n549 | n673) & (n179 | ~n679);
  assign n741 = n489 & (e | n254);
  assign n742 = ~n629 | k | n206;
  assign n743 = ~n546 & (n537 | n554);
  assign n744 = n743 & (n199 | (n714 & n713));
  assign n745 = (n720 | n376) & (n533 | n167);
  assign n746 = (n192 | n327) & (~i | n503);
  assign n747 = n745 & n746 & (n591 | n445);
  assign n748 = ~h & (n559 | (~n601 & ~n673));
  assign n749 = (n588 | n202) & (n237 | n646);
  assign n750 = n53 & n47 & n618;
  assign n751 = n526 | n102 | n120;
  assign n752 = n751 & (n651 | (n104 & n195));
  assign n753 = n449 | n480;
  assign n754 = ~n473 | h | n179;
  assign n755 = n467 | ~h | n375;
  assign n756 = i & ~k & (~n376 | ~n613);
  assign n757 = (n495 & (~h | n511)) | (h & n511);
  assign n758 = ~h & (~n96 | (c & ~n457));
  assign n759 = (n464 & (~g | n486)) | (g & n486);
  assign n760 = l | n368;
  assign n761 = n760 & n512 & n527;
  assign n762 = n674 & ~n167 & n460;
endmodule


