// Benchmark "TOP" written by ABC on Mon Feb  4 10:08:03 2019

module alu4 ( 
    i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_,
    i_11_, i_12_, i_13_,
    o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_  );
  input  i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_,
    i_10_, i_11_, i_12_, i_13_;
  output o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_;
  wire n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
    n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
    n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
    n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
    n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
    n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
    n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
    n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
    n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
    n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
    n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
    n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
    n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
    n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
    n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
    n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
    n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
    n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
    n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
    n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
    n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
    n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
    n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
    n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
    n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
    n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
    n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
    n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
    n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
    n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
    n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
    n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
    n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
    n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
    n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
    n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
    n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
    n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
    n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
    n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751;
  assign o_0_ = ~n42;
  assign o_1_ = ~n509;
  assign o_2_ = ~n502;
  assign o_3_ = ~n488;
  assign o_4_ = ~n41;
  assign o_5_ = ~n659 | ~n662 | n40 | ~n658 | n38 | n39 | n36 | n37;
  assign o_6_ = ~n35;
  assign o_7_ = ~n636 | ~n637 | n34 | ~n576 | n32 | n33 | n30 | n31;
  assign n30 = ~i_9_ & (~n163 | n165 | n168);
  assign n31 = i_9_ & n65 & n419;
  assign n32 = ~i_5_ & (~n625 | (~n238 & n250));
  assign n33 = i_9_ & (n66 | ~n621 | ~n622);
  assign n34 = n244 | n246 | n240 | n242 | ~n630 | ~n632 | n248 | n249;
  assign n35 = n278 & n279 & (~i_2_ | n277);
  assign n36 = i_11_ & (~n650 | (~n266 & n360));
  assign n37 = i_2_ & n361 & n272;
  assign n38 = ~n71 & ~n532;
  assign n39 = ~n562 & (~n648 | (~i_13_ & ~n532));
  assign n40 = ~i_4_ & (~n647 | (~n59 & ~n281));
  assign n41 = n473 & n472 & n471 & n470 & n469 & ~n465 & ~n459 & ~n461;
  assign n42 = ~n46 & n510 & (~i_0_ | n511);
  assign n43 = ~i_1_ | ~i_3_;
  assign n44 = ~i_5_ | n43;
  assign n45 = ~i_8_ & i_10_;
  assign n46 = i_3_ & (n45 | ~n435);
  assign n47 = ~n67 & (~i_6_ | ~i_10_);
  assign n48 = (n521 | n52) & (n56 | n120);
  assign n49 = i_1_ | n445;
  assign n50 = i_11_ | n116;
  assign n51 = n48 & (n49 | n50);
  assign n52 = i_12_ | n116;
  assign n53 = i_0_ | n225;
  assign n54 = (i_11_ | n53) & (n49 | n52);
  assign n55 = ~i_6_ | i_7_;
  assign n56 = i_0_ | n212;
  assign n57 = ~i_2_ | i_0_ | i_1_;
  assign n58 = (i_6_ | n57) & (n55 | n56);
  assign n59 = ~i_3_ | n225;
  assign n60 = ~i_3_ | n445;
  assign n61 = (~i_6_ | n60) & (~i_5_ | n59);
  assign n62 = i_0_ | n63;
  assign n63 = i_3_ | i_2_;
  assign n64 = n62 & (~i_5_ | n63);
  assign n65 = ~i_12_ & i_13_;
  assign n66 = n65 & (~n613 | (i_8_ & ~n379));
  assign n67 = i_6_ & n519;
  assign n68 = ~n158 & (~n615 | (n67 & ~n400));
  assign n69 = (i_7_ | n200) & (i_6_ | n62);
  assign n70 = n69 & (i_8_ | n56);
  assign n71 = ~i_12_ | n116;
  assign n72 = (~i_1_ | n71) & (~i_6_ | ~n348);
  assign n73 = ~i_1_ & i_6_;
  assign n74 = (~i_0_ | n73) & (~i_1_ | i_5_);
  assign n75 = ~n304 & ~i_9_ & ~n77;
  assign n76 = i_3_ & (n75 | (~n71 & ~n98));
  assign n77 = ~i_11_ | n116;
  assign n78 = i_8_ | i_6_;
  assign n79 = n77 | n78 | ~i_2_ | i_9_;
  assign n80 = ~i_0_ | n63;
  assign n81 = ~i_0_ | n195;
  assign n82 = (i_7_ | n81) & (i_6_ | n80);
  assign n83 = i_0_ & (n76 | ~n79 | ~n627);
  assign n84 = i_3_ | ~i_11_ | n56 | ~n348;
  assign n85 = n116 | n400 | ~i_3_ | i_9_;
  assign n86 = n178 | ~i_5_ | n72;
  assign n87 = n516 | n177 | ~n338;
  assign n88 = i_9_ | n74 | n522 | n77;
  assign n89 = n88 & n87 & n86 & n85 & ~n83 & n84;
  assign n90 = (n99 | n157) & (n134 | n521);
  assign n91 = ~i_6_ | n522;
  assign n92 = n90 & (n91 | n49);
  assign n93 = (~n102 | n521) & (~n67 | n157);
  assign n94 = (n518 | n49) & (n520 | n400);
  assign n95 = n93 & n94;
  assign n96 = (~n103 | n134) & (n53 | n107);
  assign n97 = n96 & (n57 | n91);
  assign n98 = ~i_6_ | n272;
  assign n99 = i_8_ | ~i_6_ | ~i_7_;
  assign n100 = n98 & n97 & (n99 | n56);
  assign n101 = i_5_ & n365;
  assign n102 = ~i_6_ & n519;
  assign n103 = ~i_2_ & ~i_0_ & i_1_;
  assign n104 = n101 & (~n607 | (n102 & n103));
  assign n105 = i_11_ | ~n166;
  assign n106 = i_10_ | n304;
  assign n107 = i_6_ | n522;
  assign n108 = (n107 | n50) & (n105 | n106);
  assign n109 = i_12_ | n113;
  assign n110 = i_11_ | n113;
  assign n111 = (~n67 | n109) & (n99 | n110);
  assign n112 = i_11_ | i_12_;
  assign n113 = i_9_ | i_13_;
  assign n114 = i_3_ | i_10_ | n112 | n113;
  assign n115 = i_5_ | n312;
  assign n116 = i_10_ | i_13_;
  assign n117 = (~i_10_ | n115) & (n116 | ~n164);
  assign n118 = i_13_ & (~n600 | (~n547 & ~n548));
  assign n119 = i_5_ | n515;
  assign n120 = i_12_ | ~n338;
  assign n121 = (n119 | n120) & (~n164 | ~n239);
  assign n122 = n65 & (~n599 | (~i_3_ & ~i_11_));
  assign n123 = n555 | n518 | n554;
  assign n124 = n553 | n134 | n552;
  assign n125 = n522 | n198 | ~n247;
  assign n126 = ~n348 | ~n67 | ~n101;
  assign n127 = n449 | n107 | ~n338;
  assign n128 = n524 | n99 | ~n319;
  assign n129 = (n544 | n546) & (n121 | n520);
  assign n130 = n129 & n128 & n127 & n126 & n125 & n124 & ~n122 & n123;
  assign n131 = (n107 | ~n419) & (n91 | ~n402);
  assign n132 = (n171 | n151) & (n150 | n551);
  assign n133 = n597 & n598 & (n545 | n550);
  assign n134 = ~i_7_ | n78;
  assign n135 = ~n101 | ~n239;
  assign n136 = n132 & n133 & (n134 | n135);
  assign n137 = i_4_ | ~i_0_ | ~i_1_;
  assign n138 = i_4_ | n445;
  assign n139 = (~i_6_ | n138) & (~i_7_ | n137);
  assign n140 = ~n524 & ~n220 & i_2_ & ~i_8_;
  assign n141 = n546 | n549;
  assign n142 = n162 | n107 | n158;
  assign n143 = n555 | ~n102 | n554;
  assign n144 = n553 | n91 | n552;
  assign n145 = (n194 | n151) & (n198 | n551);
  assign n146 = (n134 | n543) & (n547 | n550);
  assign n147 = n146 & n145 & n144 & n143 & n141 & n142;
  assign n148 = (n171 | n551) & (n99 | n543);
  assign n149 = n595 & n596 & (n545 | n549);
  assign n150 = ~i_5_ | n201;
  assign n151 = ~n65 | ~n264;
  assign n152 = n148 & n149 & (n150 | n151);
  assign n153 = (n99 | ~n402) & (n91 | ~n419);
  assign n154 = (n544 | n547) & (n172 | n198);
  assign n155 = n593 & n594 & (n542 | n546);
  assign n156 = n154 & n155 & (n91 | n135);
  assign n157 = ~i_0_ | n212;
  assign n158 = ~i_5_ | n312;
  assign n159 = n158 | n157 | n134;
  assign n160 = n115 | n99 | ~n103;
  assign n161 = i_2_ | n312;
  assign n162 = ~i_10_ | ~n319;
  assign n163 = n161 | n162 | ~i_5_ | n91;
  assign n164 = ~i_5_ & i_3_ & i_4_;
  assign n165 = n164 & ~n77 & i_1_ & ~i_7_;
  assign n166 = ~i_12_ & ~i_13_;
  assign n167 = i_10_ & i_11_;
  assign n168 = n166 & n167 & (~n159 | ~n160);
  assign n169 = (n542 | n545) & (n541 | n150);
  assign n170 = (n107 | n135) & (~n446 | n544);
  assign n171 = i_3_ | n539;
  assign n172 = ~n65 | ~n437;
  assign n173 = n169 & n170 & (n171 | n172);
  assign n174 = (~n446 | n542) & (n171 | n541);
  assign n175 = (n544 | n545) & (n91 | n543);
  assign n176 = n174 & n175 & (n172 | n150);
  assign n177 = i_10_ | n522;
  assign n178 = ~i_8_ | n272;
  assign n179 = n177 & n178;
  assign n180 = (~n460 | n591) & (n179 | ~n463);
  assign n181 = n592 & (n533 | n56);
  assign n182 = n106 & n98;
  assign n183 = n180 & n181 & (n182 | ~n385);
  assign n184 = (~n340 | n535) & (n106 | n449);
  assign n185 = i_8_ | n534;
  assign n186 = ~i_4_ | n212;
  assign n187 = n184 & (n185 | n186);
  assign n188 = (~n536 | n537) & (n335 | n538);
  assign n189 = (n186 | n474) & (n98 | ~n101);
  assign n190 = ~i_5_ | n272;
  assign n191 = n188 & n189 & (n190 | ~n340);
  assign n192 = (n518 | n521) & (n520 | n157);
  assign n193 = n192 & (n49 | ~n102);
  assign n194 = i_3_ | n214;
  assign n195 = i_1_ | i_3_;
  assign n196 = n194 & (~i_5_ | n195);
  assign n197 = ~i_6_ | i_0_ | i_3_;
  assign n198 = i_3_ | n516;
  assign n199 = n198 & (i_5_ | n195);
  assign n200 = i_0_ | n195;
  assign n201 = i_3_ | i_6_;
  assign n202 = n200 & n199 & (i_0_ | n201);
  assign n203 = ~i_6_ | ~i_0_ | ~i_3_;
  assign n204 = i_1_ & ~i_6_;
  assign n205 = (i_2_ | ~i_6_) & (~i_7_ | n204);
  assign n206 = n517 | i_6_ | n749;
  assign n207 = n517 | i_1_ | i_7_;
  assign n208 = i_11_ | n435;
  assign n209 = n206 & n207 & (n205 | n208);
  assign n210 = i_5_ | n63;
  assign n211 = i_2_ | n516;
  assign n212 = i_1_ | i_2_;
  assign n213 = n211 & (i_5_ | n212);
  assign n214 = ~i_5_ | ~i_6_;
  assign n215 = (~i_5_ | n212) & (i_2_ | n214);
  assign n216 = (~i_5_ | n225) & (~i_2_ | n214);
  assign n217 = ~i_6_ | n445;
  assign n218 = n216 & n217;
  assign n219 = ~i_7_ | ~i_1_ | ~i_5_;
  assign n220 = ~i_1_ & ~i_6_;
  assign n221 = n219 & (~i_0_ | ~i_7_ | n220);
  assign n222 = i_10_ & ~n435 & (~n218 | ~n221);
  assign n223 = ~i_2_ | n516;
  assign n224 = i_6_ | n445;
  assign n225 = ~i_1_ | ~i_2_;
  assign n226 = n223 & n224 & (i_5_ | n225);
  assign n227 = n226 & (i_7_ | n74);
  assign n228 = (~i_0_ | i_6_) & (~i_1_ | i_5_);
  assign n229 = (i_6_ | n138) & (i_7_ | n137);
  assign n230 = n73 | n119 | ~i_2_ | ~i_8_;
  assign n231 = n230 & (n229 | ~n475);
  assign n232 = (n53 | ~n67) & (~n103 | n518);
  assign n233 = n232 & (n57 | ~n102);
  assign n234 = ~i_4_ | n225;
  assign n235 = ~i_4_ | n557;
  assign n236 = (i_6_ | n235) & (i_8_ | n234);
  assign n237 = i_4_ & (~n623 | (~i_1_ & ~n177));
  assign n238 = ~n237 & (i_6_ | i_10_ | ~n536);
  assign n239 = ~i_9_ & n338;
  assign n240 = n239 & n164 & ~n233;
  assign n241 = n406 & ~i_10_ & ~i_13_;
  assign n242 = ~n119 & (~n580 | (~n92 & n241));
  assign n243 = ~i_3_ & ~i_8_;
  assign n244 = ~n525 & (n140 | (~n139 & n243));
  assign n245 = n383 & ~i_9_ & ~i_13_;
  assign n246 = ~n524 & (~n582 | (~n193 & n245));
  assign n247 = ~i_11_ & i_13_;
  assign n248 = n247 & (~n584 | (~n223 & ~n528));
  assign n249 = n65 & (~n586 | ~n588 | ~n590);
  assign n250 = n338 & i_12_;
  assign n251 = n250 & (~n183 | ~n187 | ~n191);
  assign n252 = ~n71 & (~n609 | ~n610 | ~n611);
  assign n253 = ~n247 & (i_4_ | ~i_8_ | ~n406);
  assign n254 = (~i_3_ | n208) & (~n338 | n533);
  assign n255 = n253 & n254 & (n120 | ~n475);
  assign n256 = ~i_7_ | i_10_;
  assign n257 = i_4_ | ~n383;
  assign n258 = (~i_7_ | n257) & (n256 | ~n318);
  assign n259 = i_7_ & n45;
  assign n260 = (i_8_ | n258) & (~n259 | n559);
  assign n261 = n260 & ~n731 & (i_7_ | n255);
  assign n262 = ~i_7_ | ~i_9_;
  assign n263 = n262 & (i_7_ | ~i_10_);
  assign n264 = i_10_ & ~i_7_ & i_8_;
  assign n265 = i_12_ & (n264 | ~n548);
  assign n266 = ~i_10_ | n522;
  assign n267 = i_8_ | n262;
  assign n268 = ~n265 & (~i_11_ | (n266 & n267));
  assign n269 = (n110 | ~n243) & (n109 | ~n475);
  assign n270 = ~i_4_ | n116;
  assign n271 = n270 & (~i_8_ | n52);
  assign n272 = ~i_7_ | i_9_;
  assign n273 = ~i_4_ | n272;
  assign n274 = (i_7_ | n271) & (i_13_ | n273);
  assign n275 = n282 & (i_4_ | n268);
  assign n276 = n556 & n638 & (i_3_ | n274);
  assign n277 = n275 & n276 & (~i_13_ | n263);
  assign n278 = ~n750 & (n548 | n559);
  assign n279 = n644 & n645 & (i_2_ | n261);
  assign n280 = ~i_6_ | ~i_9_;
  assign n281 = n280 & (i_6_ | ~i_10_);
  assign n282 = n332 | n116;
  assign n283 = (n523 & (~i_7_ | n733)) | (i_7_ & n733);
  assign n284 = i_2_ | i_13_;
  assign n285 = n282 & (n283 | n284);
  assign n286 = i_10_ | i_7_;
  assign n287 = i_11_ | n286;
  assign n288 = i_11_ | i_13_;
  assign n289 = (~n166 | n287) & (n177 | n288);
  assign n290 = i_8_ | n272;
  assign n291 = (n288 | n290) & (~n166 | n178);
  assign n292 = (n289 & (~i_6_ | n291)) | (i_6_ & n291);
  assign n293 = (n523 & (~i_8_ | n733)) | (i_8_ & n733);
  assign n294 = n292 & (i_13_ | n293);
  assign n295 = (~i_7_ & n566) | (n565 & (i_7_ | n566));
  assign n296 = i_7_ | n435;
  assign n297 = n295 & (~i_6_ | ~i_11_ | n296);
  assign n298 = n287 & (i_12_ | n256);
  assign n299 = ~i_2_ & ~n751 & (i_6_ | ~n298);
  assign n300 = ~n299 & (~i_4_ | ~n578);
  assign n301 = n591 | i_2_ | ~i_4_;
  assign n302 = n300 & n301 & (n182 | ~n365);
  assign n303 = ~i_7_ | n280;
  assign n304 = i_6_ | i_7_;
  assign n305 = n303 & (~i_10_ | (~i_9_ & n304));
  assign n306 = (i_6_ & ~n540) | (~n266 & (~i_6_ | ~n540));
  assign n307 = ~i_4_ & (~n577 | (i_11_ & n306));
  assign n308 = (n294 & (~i_3_ | n297)) | (i_3_ & n297);
  assign n309 = (~i_13_ & n302) | (n281 & (i_13_ | n302));
  assign n310 = ~n307 & n656 & (~i_2_ | n305);
  assign n311 = n310 & n309 & n308 & n285;
  assign n312 = ~i_3_ | i_4_;
  assign n313 = (n312 | ~n406) & (n284 | ~n383);
  assign n314 = (~i_4_ | ~n338) & (i_3_ | n120);
  assign n315 = ~n247 & (~i_3_ | ~n406 | n548);
  assign n316 = (~i_2_ | n530) & (~i_7_ | n313);
  assign n317 = n315 & n316 & (n314 | n178);
  assign n318 = i_4_ & n348;
  assign n319 = ~i_11_ & n348;
  assign n320 = ~n177 & (n318 | (~i_3_ & n319));
  assign n321 = ~n402 | ~i_2_ | i_7_;
  assign n322 = ~n319 | n563;
  assign n323 = ~n383 | ~i_3_ | n266;
  assign n324 = n257 | ~i_2_ | i_8_;
  assign n325 = ~n65 & (i_7_ | n312 | ~n383);
  assign n326 = n325 & n324 & n323 & n322 & ~n320 & n321;
  assign n327 = i_11_ | ~n496 | n558 | ~n563;
  assign n328 = (n317 & (~i_6_ | n326)) | (i_6_ & n326);
  assign n329 = n327 & n328 & (n91 | n257);
  assign n330 = ~i_11_ | n514;
  assign n331 = ~n166 | ~n475;
  assign n332 = ~i_4_ | i_9_;
  assign n333 = (n332 | n77) & (n330 | n331);
  assign n334 = ~n517 & i_3_ & i_12_;
  assign n335 = i_1_ | n63;
  assign n336 = ~i_11_ | ~n166;
  assign n337 = (n335 | n336) & (n186 | ~n239);
  assign n338 = i_11_ & ~i_13_;
  assign n339 = i_4_ & (~n652 | (~n335 & n338));
  assign n340 = ~i_1_ & n365;
  assign n341 = i_7_ & (n334 | (n340 & n239));
  assign n342 = n734 & (~i_8_ | n337);
  assign n343 = (n208 | n561) & (n404 | n356);
  assign n344 = (n517 | n557) & (~n45 | n59);
  assign n345 = n344 & n343 & n342 & ~n341 & n333 & ~n339;
  assign n346 = ~i_2_ | i_12_;
  assign n347 = (~i_8_ | n59) & (n346 | ~n391);
  assign n348 = i_12_ & ~i_13_;
  assign n349 = n348 & (~n654 | (i_4_ & ~n335));
  assign n350 = n655 & (i_8_ | ~n402 | n561);
  assign n351 = ~n349 & n350 & (~i_9_ | n347);
  assign n352 = ~i_8_ | i_9_;
  assign n353 = (~n263 | ~n340) & (n186 | n352);
  assign n354 = i_10_ | n78;
  assign n355 = ~i_6_ | n352;
  assign n356 = ~i_1_ | n312;
  assign n357 = (n303 | n356) & (~n259 | ~n360);
  assign n358 = ~n573 & (~i_4_ | i_13_ | ~n496);
  assign n359 = ~n512 & (i_6_ | i_11_);
  assign n360 = i_3_ & n204;
  assign n361 = ~i_6_ & n419;
  assign n362 = ~i_9_ | ~i_11_;
  assign n363 = ~i_12_ | n362;
  assign n364 = ~i_4_ | n113;
  assign n365 = ~i_3_ & i_4_;
  assign n366 = ~i_9_ | ~i_12_;
  assign n367 = n364 & (n365 | n366);
  assign n368 = (~i_9_ & n572) | (~i_13_ & (i_9_ | n572));
  assign n369 = i_3_ | n111;
  assign n370 = ~n166 | i_2_ | n98;
  assign n371 = (~i_1_ | n280) & (n363 | ~n391);
  assign n372 = (~n67 | n367) & (i_4_ | n363);
  assign n373 = ~n737 & n372 & n371 & n370 & n368 & n369;
  assign n374 = ~i_4_ & (~n564 | (~n107 & n167));
  assign n375 = ~n736 & (~i_10_ | (~i_13_ & ~n204));
  assign n376 = ~n374 & n687 & (n107 | n270);
  assign n377 = n375 & n376 & (i_3_ | n108);
  assign n378 = i_7_ | n516;
  assign n379 = ~i_7_ | n214;
  assign n380 = (n113 | n379) & (n378 | n116);
  assign n381 = ~i_2_ & (~n686 | (~n270 & ~n440));
  assign n382 = ~n53 & i_3_ & ~i_8_;
  assign n383 = i_11_ & ~i_12_;
  assign n384 = n383 & i_10_ & ~i_0_ & i_2_;
  assign n385 = ~i_0_ & n365;
  assign n386 = ~i_6_ & (n384 | (~n71 & n385));
  assign n387 = (n56 | ~n319) & (n53 | ~n402);
  assign n388 = i_0_ | n43;
  assign n389 = ~n386 & n387 & (n257 | n388);
  assign n390 = (~i_7_ | n81) & (~i_6_ | n80);
  assign n391 = i_8_ & i_3_;
  assign n392 = ~n400 & (i_7_ | n391);
  assign n393 = (i_3_ & n553) | (~n241 & (~i_3_ | n553));
  assign n394 = n257 & n393 & (~i_4_ | n71);
  assign n395 = ~i_12_ | n572;
  assign n396 = ~n65 & (i_2_ | n106 | ~n319);
  assign n397 = n395 & n396 & (n394 | n107);
  assign n398 = ~i_7_ | n362;
  assign n399 = (i_2_ | n355) & (n204 | n178);
  assign n400 = ~i_1_ | n445;
  assign n401 = (~i_8_ | n400) & (~i_6_ | n60);
  assign n402 = i_10_ & ~i_12_;
  assign n403 = n402 & (n382 | (~i_0_ & n204));
  assign n404 = i_7_ | ~n167;
  assign n405 = n167 & (~n718 | (~i_8_ & ~n400));
  assign n406 = ~i_11_ & i_12_;
  assign n407 = n406 & (~n674 | (i_8_ & ~n53));
  assign n408 = ~i_0_ | n43;
  assign n409 = ~n405 & ~n407 & (n404 | n408);
  assign n410 = ~n247 & (~i_1_ | i_11_ | n280);
  assign n411 = n672 & (~n67 | (~n423 & n673));
  assign n412 = n410 & n411 & (~n73 | n336);
  assign n413 = ~n385 | ~i_6_ | ~n239;
  assign n414 = ~n166 | ~i_11_ | n56;
  assign n415 = n413 & n414 & (n200 | ~n423);
  assign n416 = n238 & (~i_4_ | i_6_ | n177);
  assign n417 = ~i_7_ & n419;
  assign n418 = n417 & i_2_ & i_12_;
  assign n419 = i_10_ & ~i_11_;
  assign n420 = n116 | ~i_4_ | i_8_;
  assign n421 = n420 & (n50 | ~n243);
  assign n422 = ~n53 & (~n530 | (i_3_ & ~n208));
  assign n423 = i_4_ & n239;
  assign n424 = i_6_ & (n418 | (~n62 & n423));
  assign n425 = (n517 | n59) & (i_4_ | n409);
  assign n426 = (~i_7_ | n415) & (i_0_ | n412);
  assign n427 = (n82 | n271) & (~n338 | n416);
  assign n428 = (~i_1_ | ~n361) & (~n423 | n671);
  assign n429 = (n157 | n421) & (n400 | ~n670);
  assign n430 = ~n422 & (n56 | n120 | ~n475);
  assign n431 = n430 & n429 & n428 & n427 & n426 & n425 & n333 & ~n424;
  assign n432 = n183 & (~i_4_ | i_10_ | n70);
  assign n433 = i_7_ | i_9_ | i_11_;
  assign n434 = n191 & (n215 | n433);
  assign n435 = ~i_8_ | ~i_9_;
  assign n436 = i_5_ & ~n558 & (~n540 | ~n568);
  assign n437 = i_10_ & n519;
  assign n438 = ~i_4_ & ~n539 & (n437 | ~n568);
  assign n439 = ~i_8_ | n214;
  assign n440 = i_8_ | n516;
  assign n441 = (n366 | n439) & (~n167 | n440);
  assign n442 = ~i_12_ & (~n158 | n417 | ~n530);
  assign n443 = n435 | ~i_3_ | n112;
  assign n444 = ~n442 & n443 & (i_11_ | n115);
  assign n445 = ~i_0_ | ~i_2_;
  assign n446 = ~i_6_ & i_3_ & i_5_;
  assign n447 = n383 & (~n684 | (~i_7_ & n446));
  assign n448 = n406 & (~n685 | (i_7_ & ~n545));
  assign n449 = i_5_ | ~n365;
  assign n450 = (~n338 | n449) & (~n101 | ~n348);
  assign n451 = i_5_ | n522;
  assign n452 = (n80 | n440) & (n81 | n451);
  assign n453 = ~i_5_ | ~n519;
  assign n454 = (n453 | n81) & (n439 | n80);
  assign n455 = n137 & n408;
  assign n456 = ~i_0_ | n312;
  assign n457 = (n379 | n456) & (n455 | n453);
  assign n458 = ~i_5_ & i_0_ & i_3_;
  assign n459 = n167 & (~n663 | (~n107 & n458));
  assign n460 = i_4_ & ~i_0_ & ~i_2_;
  assign n461 = ~n569 & (~n664 | (n239 & n460));
  assign n462 = ~i_5_ & n519;
  assign n463 = i_4_ & ~i_0_ & ~i_1_;
  assign n464 = n462 & (~n665 | (n239 & n463));
  assign n465 = ~n570 & (~n666 | (~n71 & n463));
  assign n466 = ~n571 & (~n667 | (~n71 & n460));
  assign n467 = n406 & (n438 | (n259 & ~n545));
  assign n468 = n383 & (n436 | (~n296 & n446));
  assign n469 = (n450 | n56) & (n441 | n60);
  assign n470 = ~n464 & (~i_9_ | n158 | n400);
  assign n471 = n702 & n701 & (n452 | n50);
  assign n472 = n699 & n698 & (n457 | n366);
  assign n473 = ~n740 & ~n739 & n709 & n707 & n706 & n705 & n703 & n704;
  assign n474 = ~i_5_ | n352;
  assign n475 = ~i_3_ & i_8_;
  assign n476 = ~n56 & (i_7_ | n475);
  assign n477 = (i_1_ | n537) & (n589 | n178);
  assign n478 = ~n476 & n715 & (n335 | n474);
  assign n479 = n477 & n478 & (i_0_ | ~i_5_);
  assign n480 = ~n56 & (~i_7_ | n243);
  assign n481 = n300 & (i_1_ | n359);
  assign n482 = n746 & (i_5_ | n416);
  assign n483 = n187 & (i_3_ | n293);
  assign n484 = (n56 | ~n365) & (i_12_ | n479);
  assign n485 = (n213 | n298) & (n215 | n574);
  assign n486 = n716 & (i_1_ | n359 | n534);
  assign n487 = n717 & (i_11_ | (n714 & n711));
  assign n488 = n487 & n486 & n485 & n484 & n483 & n482 & n432 & n434;
  assign n489 = ~i_7_ | n366;
  assign n490 = ~i_10_ | ~i_12_;
  assign n491 = n489 & ~n496 & (i_7_ | n490);
  assign n492 = (n747 & (~i_5_ | n748)) | (i_5_ & n748);
  assign n493 = n492 & (~i_0_ | n281);
  assign n494 = i_8_ | ~i_11_;
  assign n495 = ~n496 & n494 & ~i_3_ & n263;
  assign n496 = i_8_ & i_12_;
  assign n497 = n496 & (~n221 | ~n379);
  assign n498 = (n218 | n491) & (~i_1_ | n493);
  assign n499 = n726 & (~i_12_ | (n61 & n723));
  assign n500 = n725 & (~i_11_ | (n719 & n722));
  assign n501 = n724 & (n494 | (n227 & n378));
  assign n502 = n501 & n500 & n498 & n499;
  assign n503 = i_12_ | ~n475;
  assign n504 = ~n46 & n503 & (i_11_ | ~n243);
  assign n505 = (~n243 | ~n338) & (n113 | ~n391);
  assign n506 = (~n243 | ~n247) & (~n65 | ~n475);
  assign n507 = (n504 & (~i_4_ | n505)) | (i_4_ & n505);
  assign n508 = n727 & n728 & (~i_13_ | ~n46);
  assign n509 = n508 & n506 & n507;
  assign n510 = (~i_1_ | n281) & (~i_2_ | n263);
  assign n511 = (~i_5_ & ~i_10_) | (~i_9_ & (i_5_ | ~i_10_));
  assign n512 = i_6_ & ~i_12_;
  assign n513 = i_9_ & (n392 | (n512 & i_1_));
  assign n514 = i_9_ | i_10_;
  assign n515 = i_3_ | i_4_;
  assign n516 = i_5_ | i_6_;
  assign n517 = i_8_ | ~n419;
  assign n518 = ~i_8_ | n55;
  assign n519 = i_8_ & i_7_;
  assign n520 = ~i_8_ | n304;
  assign n521 = i_2_ | ~i_0_ | ~i_1_;
  assign n522 = i_8_ | i_7_;
  assign n523 = i_11_ | n514;
  assign n524 = ~i_5_ | n515;
  assign n525 = ~n348 | n523;
  assign n526 = ~i_9_ | ~i_10_;
  assign n527 = i_7_ | n526;
  assign n528 = ~i_3_ | n526;
  assign n529 = ~i_7_ | n526;
  assign n530 = i_11_ | n262;
  assign n531 = ~i_5_ | ~i_3_ | ~i_4_;
  assign n532 = ~i_6_ | n332;
  assign n533 = ~i_8_ | n332;
  assign n534 = i_5_ | i_10_;
  assign n535 = i_7_ | n534;
  assign n536 = ~i_2_ & n365;
  assign n537 = i_9_ | n214;
  assign n538 = ~i_5_ | n332;
  assign n539 = i_5_ | ~i_6_;
  assign n540 = ~i_9_ | n522;
  assign n541 = ~n247 | n540;
  assign n542 = ~n65 | ~n259;
  assign n543 = ~n239 | n449;
  assign n544 = ~n247 | n296;
  assign n545 = ~i_3_ | n539;
  assign n546 = ~i_3_ | n516;
  assign n547 = ~i_3_ | n214;
  assign n548 = ~i_7_ | n435;
  assign n549 = ~n247 | n548;
  assign n550 = ~n65 | n266;
  assign n551 = ~n247 | n267;
  assign n552 = i_13_ | n115;
  assign n553 = ~i_11_ | ~n402;
  assign n554 = i_13_ | n158;
  assign n555 = ~i_9_ | ~n406;
  assign n556 = n114 & n528;
  assign n557 = ~i_2_ | ~i_3_;
  assign n558 = i_4_ | i_6_;
  assign n559 = ~i_3_ | i_12_;
  assign n560 = i_4_ | n225;
  assign n561 = i_1_ | n557;
  assign n562 = ~i_1_ | n63;
  assign n563 = i_7_ | i_2_;
  assign n564 = ~i_11_ | n490;
  assign n565 = ~i_9_ | n490;
  assign n566 = ~i_9_ | ~n167;
  assign n567 = ~i_8_ | n286;
  assign n568 = i_0_ | n557;
  assign n569 = ~i_8_ | n539;
  assign n570 = ~i_5_ | n522;
  assign n571 = ~i_5_ | n78;
  assign n572 = ~n220 | n288;
  assign n573 = n243 & n319;
  assign n574 = i_12_ | n272;
  assign n575 = (~i_5_ & n419) | (n402 & (i_5_ | n419));
  assign n576 = (~i_4_ & n729) | (n89 & (i_4_ | n729));
  assign n577 = (~i_6_ & n564) | (n363 & (i_6_ | n564));
  assign n578 = (i_6_ & ~n178) | (~n177 & (~i_6_ | ~n178));
  assign n579 = i_10_ | i_13_ | ~n383 | n520;
  assign n580 = n579 & (n233 | ~n245);
  assign n581 = i_9_ | i_13_ | n99 | ~n406;
  assign n582 = n581 & (n97 | ~n241);
  assign n583 = n527 | ~i_3_ | n228;
  assign n584 = n583 & (i_8_ | n227 | n526);
  assign n585 = (n213 | n517) & (n210 | ~n361);
  assign n586 = ~n222 & n585 & (n208 | n215);
  assign n587 = n547 & n408 & n44 & n203;
  assign n588 = (n587 | n529) & (i_0_ | n209);
  assign n589 = n196 & n200 & n197;
  assign n590 = (n530 | n589) & (n202 | ~n417);
  assign n591 = n355 & n354;
  assign n592 = (n273 | n200) & (n62 | n532);
  assign n593 = n541 | n194;
  assign n594 = n113 | n153 | n158;
  assign n595 = ~n402 | n107 | n158;
  assign n596 = ~n446 | n550;
  assign n597 = ~n446 | n549;
  assign n598 = n113 | n131 | n158;
  assign n599 = (~n259 | n547) & (n194 | ~n519);
  assign n600 = n528 & (n546 | n266);
  assign n601 = n531 | ~n67 | n113;
  assign n602 = n601 & (n117 | n107);
  assign n603 = (n99 | n135) & (n198 | n151);
  assign n604 = n602 & n603 & (n194 | n551);
  assign n605 = (n108 | n119) & (n111 | n524);
  assign n606 = ~n118 & n605 & (i_4_ | n556);
  assign n607 = (n518 | n57) & (n53 | n520);
  assign n608 = (n95 | n449) & (n92 | ~n164);
  assign n609 = ~n104 & n608 & (n100 | n531);
  assign n610 = (n537 | n235) & (n474 | n234);
  assign n611 = (n273 | n408) & (n538 | n59);
  assign n612 = n64 | ~i_6_ | i_11_;
  assign n613 = n612 & (~i_10_ | n61);
  assign n614 = i_10_ | ~n103 | ~n319 | n520;
  assign n615 = n614 & (n58 | n162);
  assign n616 = i_10_ | n157 | ~n319 | n518;
  assign n617 = n616 & (n47 | n57 | n120);
  assign n618 = n617 & (n520 | n521 | n50);
  assign n619 = (n54 | ~n67) & (n51 | ~n102);
  assign n620 = n161 | n534 | ~n102 | n120;
  assign n621 = n620 & (i_4_ | n59 | ~n575);
  assign n622 = ~n68 & (n115 | (n618 & n619));
  assign n623 = (i_2_ | n354) & (i_10_ | n335);
  assign n624 = i_11_ | n266 | n59 | n558;
  assign n625 = n624 & (i_9_ | n236 | n77);
  assign n626 = n355 | ~i_2_ | n71;
  assign n627 = n626 & (n220 | n71 | n178);
  assign n628 = n332 | i_10_ | ~n250;
  assign n629 = n628 & (~n166 | n231 | n330);
  assign n630 = n629 & (~i_13_ | n378 | n517);
  assign n631 = n531 | n193 | ~n239;
  assign n632 = ~n251 & n631 & (~n103 | n176);
  assign n633 = (n156 | n521) & (n173 | n157);
  assign n634 = n633 & (n152 | n53);
  assign n635 = (n136 | n49) & (n147 | n57);
  assign n636 = n635 & n634 & (n130 | n56);
  assign n637 = ~n252 & (n400 | (n604 & n606));
  assign n638 = n730 & (~i_7_ | n269);
  assign n639 = ~n435 | ~i_4_ | n77;
  assign n640 = n639 & (i_8_ | i_13_ | n235);
  assign n641 = (i_11_ | n161) & (~n338 | ~n536);
  assign n642 = n235 | ~i_8_ | i_13_;
  assign n643 = n642 & (~n348 | (n533 & ~n536));
  assign n644 = n312 | ~i_2_ | n263;
  assign n645 = ~n732 & (i_7_ | (n640 & n641));
  assign n646 = ~n563 | ~n361 | ~n496;
  assign n647 = n646 & (n359 | n561);
  assign n648 = (n288 | n354) & (~n166 | n355);
  assign n649 = ~i_8_ | i_3_ | i_6_ | n749 | i_10_ | ~n166;
  assign n650 = n649 & (~n348 | n353);
  assign n651 = i_10_ | i_13_ | n749 | n494;
  assign n652 = n651 & (n116 | n562);
  assign n653 = i_10_ | i_8_;
  assign n654 = (n286 | ~n340) & (n186 | n653);
  assign n655 = n335 | i_8_ | ~n319;
  assign n656 = n365 | n548 | ~i_6_ | ~i_12_;
  assign n657 = ~i_3_ | ~i_9_ | ~n383 | n518;
  assign n658 = n657 & (n281 | ~n496 | n560);
  assign n659 = (n358 | n98) & (n346 | n303);
  assign n660 = (n345 & (~i_6_ | n351)) | (i_6_ & n351);
  assign n661 = (~i_1_ & n329) | (n311 & (i_1_ | n329));
  assign n662 = n660 & n661 & (~i_12_ | n357);
  assign n663 = (n378 | n456) & (n455 | n451);
  assign n664 = (n555 | n568) & (n62 | ~n245);
  assign n665 = (n388 | n555) & (n200 | ~n245);
  assign n666 = (n388 | n553) & (n200 | ~n241);
  assign n667 = (n553 | n568) & (n62 | ~n241);
  assign n668 = (n288 | n535) & (~n166 | n190);
  assign n669 = (n116 | n449) & (~n101 | n113);
  assign n670 = i_10_ & (~i_7_ | (i_3_ & ~i_8_));
  assign n671 = ~i_8_ | n56;
  assign n672 = n741 & (~i_2_ | n303 | ~n406);
  assign n673 = (i_3_ & n555) | (~n245 & (~i_3_ | n555));
  assign n674 = (~i_7_ | n388) & (i_0_ | ~n67);
  assign n675 = ~n383 | i_8_ | n53;
  assign n676 = n675 & (n401 | n366);
  assign n677 = n157 | ~i_8_ | n113;
  assign n678 = n677 & (~n348 | n399);
  assign n679 = n346 | i_6_ | n398;
  assign n680 = n679 & (n390 | n364);
  assign n681 = (~n243 | n525) & (n157 | n269);
  assign n682 = n680 & n681 & (n56 | ~n573);
  assign n683 = (i_7_ | n389) & (i_0_ | n397);
  assign n684 = (~i_2_ | n571) & (~i_1_ | n570);
  assign n685 = (~i_2_ | n569) & (~i_1_ | ~n462);
  assign n686 = (n364 | n439) & (n105 | n537);
  assign n687 = n288 | i_2_ | n106;
  assign n688 = (n451 | n270) & (n364 | n453);
  assign n689 = n211 | i_10_ | n105;
  assign n690 = n689 & (~i_9_ | n536 | n564);
  assign n691 = ~n381 & n690 & (~n365 | n380);
  assign n692 = i_3_ | i_13_ | n293;
  assign n693 = n735 & (~i_6_ | ~i_12_ | n529);
  assign n694 = n285 & n692 & (~i_3_ | n693);
  assign n695 = (~i_5_ & n377) | (n373 & (i_5_ | n377));
  assign n696 = n695 & ~n738 & (~i_1_ | n526);
  assign n697 = n564 | i_8_ | ~n458;
  assign n698 = n697 & (n213 | n256 | n336);
  assign n699 = n400 | ~i_10_ | n115;
  assign n700 = n567 | n199 | n120;
  assign n701 = n700 & (n454 | n109);
  assign n702 = ~n319 | n196 | n290;
  assign n703 = ~n466 & (n157 | (n668 & n669));
  assign n704 = (n444 | n53) & (n217 | n565);
  assign n705 = ~n467 & ~n468 & (n138 | n441);
  assign n706 = (~n348 | n434) & (~n250 | n432);
  assign n707 = (n538 | n71) & (n566 | n224);
  assign n708 = n445 | i_5_ | n512 | n404;
  assign n709 = n708 & ~n745 & (i_5_ | n431);
  assign n710 = (n589 | n290) & (n202 | n177);
  assign n711 = ~n480 & n710 & (n62 | n354);
  assign n712 = (n185 | n335) & (n210 | n354);
  assign n713 = ~n220 | ~i_5_ | i_9_;
  assign n714 = n713 & n712 & (i_0_ | i_5_);
  assign n715 = (n202 | n567) & (n64 | n355);
  assign n716 = i_10_ | n332;
  assign n717 = (i_2_ | n283) & (i_0_ | n481);
  assign n718 = i_6_ | n60;
  assign n719 = ~i_12_ & n718 & (i_5_ | n59);
  assign n720 = n228 | ~i_3_ | i_7_;
  assign n721 = n720 & (i_7_ | n408);
  assign n722 = n721 & (n546 | (~i_2_ & i_7_));
  assign n723 = (~i_7_ | n587) & (~i_2_ | n547);
  assign n724 = ~n497 & (n226 | (n398 & n404));
  assign n725 = ~i_0_ | n511;
  assign n726 = n495 | n400;
  assign n727 = ~n435 | ~i_3_ | n270;
  assign n728 = ~n365 | ~i_8_ | ~n348;
  assign n729 = ~i_5_ | n59 | ~n512 | n548;
  assign n730 = ~n243 | i_7_ | n50;
  assign n731 = i_7_ & (n573 | n65);
  assign n732 = i_7_ & (~n643 | (~i_12_ & ~n161));
  assign n733 = i_12_ | n514;
  assign n734 = n560 | i_8_ | ~n167;
  assign n735 = n527 | i_6_ | ~i_11_;
  assign n736 = ~i_10_ & (~n572 | (n73 & n166));
  assign n737 = i_2_ & i_12_ & (~n303 | ~n398);
  assign n738 = ~i_1_ & (~n688 | (n166 & ~n537));
  assign n739 = ~i_0_ & ~i_4_ & (n447 | n448);
  assign n740 = i_0_ & (~n691 | ~n694 | ~n696);
  assign n741 = i_2_ | n98 | n120;
  assign n742 = i_4_ & (~n678 | (~n70 & ~n71));
  assign n743 = ~i_4_ & (~n676 | (~n408 & ~n489));
  assign n744 = ~n682 | n403 | n513 | n743 | ~n683 | n742;
  assign n745 = i_5_ & n744;
  assign n746 = n399 | ~i_4_ | ~i_5_;
  assign n747 = (i_6_ & n362) | (~n167 & (~i_6_ | n362));
  assign n748 = (~i_6_ & n490) | (n366 & (i_6_ | n490));
  assign n749 = i_2_ & i_7_;
  assign n750 = n417 & n533 & i_3_;
  assign n751 = i_6_ & n574 & n433;
endmodule


