// Benchmark "TOP" written by ABC on Mon Feb  4 17:31:22 2019

module ex1010 ( 
    i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_,
    o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_  );
  input  i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_;
  output o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_;
  wire n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
    n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
    n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
    n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
    n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
    n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
    n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
    n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
    n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
    n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
    n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
    n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
    n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
    n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
    n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
    n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
    n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
    n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
    n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
    n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
    n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
    n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
    n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
    n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
    n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
    n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
    n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
    n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
    n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
    n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
    n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
    n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
    n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
    n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
    n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
    n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
    n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
    n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
    n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
    n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
    n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
    n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
    n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
    n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
    n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
    n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
    n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
    n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
    n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
    n868, n869;
  assign o_0_ = ~n418;
  assign o_1_ = ~n31;
  assign o_2_ = ~n403;
  assign o_3_ = ~n378;
  assign o_4_ = ~n349;
  assign o_5_ = ~n30;
  assign o_6_ = ~n270;
  assign o_7_ = ~n216;
  assign o_8_ = ~n170;
  assign o_9_ = ~n109;
  assign n30 = n155 & n50 & n301 & n302 & n303 & n304 & n305 & n306;
  assign n31 = n97 & n404 & n151 & n405 & n406 & n407 & n408 & n409;
  assign n32 = (n436 | n458) & (n219 | n479);
  assign n33 = ~i_9_ | n429;
  assign n34 = n423 | n446;
  assign n35 = n32 & (n33 | n34);
  assign n36 = (n222 | n481) & (n43 | n480);
  assign n37 = ~i_9_ | n419;
  assign n38 = n423 | n457;
  assign n39 = n36 & (n37 | n38);
  assign n40 = i_9_ | n440;
  assign n41 = n420 | n441;
  assign n42 = n419 | n450;
  assign n43 = i_9_ | n421;
  assign n44 = (n42 | n43) & (n40 | n41);
  assign n45 = n219 | n103;
  assign n46 = n439 | n290;
  assign n47 = n565 & n320 & n566;
  assign n48 = n563 & n564 & (n272 | n476);
  assign n49 = n561 & n562 & n125 & n556 & n560 & n557;
  assign n50 = n45 & n46 & n44 & n35 & n39 & n47 & n48 & n49;
  assign n51 = n40 | n456;
  assign n52 = n436 | n203;
  assign n53 = ~i_9_ | n427;
  assign n54 = n426 | n446;
  assign n55 = n51 & n52 & (n53 | n54);
  assign n56 = n37 | n262;
  assign n57 = n272 | n487;
  assign n58 = n319 & (n219 | n488);
  assign n59 = n555 & n55 & (n91 | n489);
  assign n60 = n53 | n92;
  assign n61 = n219 | n485;
  assign n62 = n33 | n486;
  assign n63 = n388 & n554 & (n53 | n483);
  assign n64 = n56 & n57 & n58 & n59 & n60 & n61 & n62 & n63;
  assign n65 = n552 & (n37 | n490);
  assign n66 = n436 | n491;
  assign n67 = (n33 | n469) & (n96 | n43);
  assign n68 = n219 | n339;
  assign n69 = (n37 | n478) & (n439 | n494);
  assign n70 = n553 & n328 & (n309 | n481);
  assign n71 = n65 & n66 & n67 & n68 & n69 & n70;
  assign n72 = n91 | n496;
  assign n73 = n100 | n41;
  assign n74 = (n309 | n463) & (n222 | n495);
  assign n75 = (n222 | n463) & (n43 | n255);
  assign n76 = (n422 | n462) & (n43 | n223);
  assign n77 = n72 & n73 & n74 & n75 & n76;
  assign n78 = n219 | n498;
  assign n79 = n436 | n480;
  assign n80 = (n436 | n447) & (n222 | n497);
  assign n81 = (n86 | n475) & (n258 | n499);
  assign n82 = (n309 | n480) & (n40 | n493);
  assign n83 = n78 & n79 & n80 & n81 & n82;
  assign n84 = (n443 | n86) & (n462 | n502);
  assign n85 = n225 & n551 & (n258 | n500);
  assign n86 = i_9_ | n460;
  assign n87 = n433 | n466;
  assign n88 = n84 & n85 & (n86 | n87);
  assign n89 = (n222 | n203) & (n33 | n150);
  assign n90 = n549 & n550 & (n219 | n199);
  assign n91 = ~i_9_ | n466;
  assign n92 = n435 | n442;
  assign n93 = n89 & n90 & (n91 | n92);
  assign n94 = n462 | n507;
  assign n95 = n548 & n124 & (n100 | n506);
  assign n96 = n441 | n442;
  assign n97 = n94 & n95 & (n96 | n86);
  assign n98 = (n219 | n92) & (n53 | n469);
  assign n99 = n431 | n432;
  assign n100 = i_9_ | n457;
  assign n101 = n98 & (n99 | n100);
  assign n102 = (n100 | n508) & (n33 | n489);
  assign n103 = n423 | n460;
  assign n104 = n102 & (n37 | n103);
  assign n105 = (n86 | n465) & (n464 | n219);
  assign n106 = n64 & n71 & n50 & n83 & n88 & n77;
  assign n107 = n589 & n593 & n592 & n586 & n585 & n588;
  assign n108 = n580 & n584 & n583 & n579 & n577 & n575;
  assign n109 = n97 & n101 & n93 & n105 & n104 & n106 & n107 & n108;
  assign n110 = n623 & (n100 | n514);
  assign n111 = n37 | n507;
  assign n112 = n86 | (n468 & n492);
  assign n113 = n622 & (n462 | n498);
  assign n114 = n620 & n621 & (n43 | n310);
  assign n115 = n619 & n285 & n561 & n209 & n56 & n618 & n299 & n616;
  assign n116 = n110 & n111 & n112 & n113 & n114 & n115;
  assign n117 = (n37 | n471) & (n33 | n520);
  assign n118 = n53 | n34;
  assign n119 = (n91 | n523) & (n462 | n488);
  assign n120 = n609 & n608 & (n100 | n475);
  assign n121 = n312 & n613 & (n309 | n458);
  assign n122 = n611 & n610 & (n447 | n43);
  assign n123 = n117 & n118 & n119 & n120 & n121 & n122;
  assign n124 = n462 | n505;
  assign n125 = n43 | n468;
  assign n126 = n73 & (n222 | n518);
  assign n127 = (n86 | n525) & (n272 | n465);
  assign n128 = n606 & (n309 | n524);
  assign n129 = n603 & (n462 | n526);
  assign n130 = n601 & n602 & (n439 | n498);
  assign n131 = n605 & n604 & (n37 | n461);
  assign n132 = n124 & n125 & n126 & n127 & n128 & n129 & n130 & n131;
  assign n133 = (n272 | n495) & (n91 | n103);
  assign n134 = n454 | n100;
  assign n135 = n600 & (n309 | n484);
  assign n136 = n462 | n477;
  assign n137 = n598 & n599 & (n219 | n500);
  assign n138 = n596 & n597 & (n222 | n42);
  assign n139 = n133 & n134 & n135 & n136 & n137 & n138;
  assign n140 = (n91 | n511) & (n272 | n528);
  assign n141 = n594 & n595 & (n91 | n34);
  assign n142 = n420 | n432;
  assign n143 = n140 & n141 & (n86 | n142);
  assign n144 = (n272 | n529) & (n258 | n503);
  assign n145 = n86 | n530;
  assign n146 = (n53 | n103) & (n424 | n462);
  assign n147 = n144 & n145 & n146 & n61;
  assign n148 = (n309 | n531) & (n436 | n456);
  assign n149 = (n86 | n532) & (n100 | n472);
  assign n150 = n421 | n442;
  assign n151 = n148 & n149 & (n91 | n150);
  assign n152 = (n40 & n436) | n533;
  assign n153 = n380 & (n53 | n496);
  assign n154 = n423 | n435;
  assign n155 = n152 & n153 & (n91 | n154);
  assign n156 = (n100 | n531) & (n91 | n534);
  assign n157 = n426 | n466;
  assign n158 = n156 & (n86 | n157);
  assign n159 = (n33 | n505) & (n91 | n38);
  assign n160 = n433 | n460;
  assign n161 = n159 & (n33 | n160);
  assign n162 = (n436 | n513) & (n33 | n92);
  assign n163 = (n53 | n509) & (n222 | n512);
  assign n164 = (n222 | n513) & (n37 | n467);
  assign n165 = (n258 | n467) & (n43 | n501);
  assign n166 = n626 & n625 & (n309 | n42);
  assign n167 = n633 & n634 & n631 & n630 & n629 & n387 & n628 & n627;
  assign n168 = n139 & n143 & n147 & n151 & n123 & n132 & n116 & n644;
  assign n169 = n640 & n641 & n639 & n638 & n637 & n642 & n636 & n635;
  assign n170 = n162 & n163 & n164 & n165 & n166 & n167 & n168 & n169;
  assign n171 = (n37 | n92) & (n43 | n484);
  assign n172 = n648 & n649 & (n458 | n86);
  assign n173 = n647 & (n100 | n294);
  assign n174 = n645 & n646 & (n219 | n540);
  assign n175 = n171 & n172 & n173 & n174;
  assign n176 = n33 | n477;
  assign n177 = n272 | n255;
  assign n178 = (n91 | n538) & (n452 | n43);
  assign n179 = n91 | n504;
  assign n180 = (n100 | n492) & (n258 | n504);
  assign n181 = n559 & (n53 | n290);
  assign n182 = n176 & n177 & n178 & n179 & n180 & n181;
  assign n183 = n428 | n100;
  assign n184 = n219 | n34;
  assign n185 = (n436 | n472) & (n43 | n474);
  assign n186 = n40 | n542;
  assign n187 = (n91 | n339) & (n445 | n219);
  assign n188 = (n40 | n525) & (n219 | n505);
  assign n189 = n183 & n184 & n185 & n186 & n187 & n188;
  assign n190 = n436 | n525;
  assign n191 = n86 | n512;
  assign n192 = (n86 | n480) & (n436 | n544);
  assign n193 = n53 | n486;
  assign n194 = n309 | n543;
  assign n195 = (n258 | n251) & (n222 | n294);
  assign n196 = n190 & n191 & n192 & n193 & n194 & n195;
  assign n197 = (n96 | n100) & (n272 | n532);
  assign n198 = n350 & n351 & (n40 | n513);
  assign n199 = n450 | n457;
  assign n200 = n197 & n198 & (n53 | n199);
  assign n201 = (n462 | n496) & (n37 | n522);
  assign n202 = (n309 | n517) & (n439 | n539);
  assign n203 = n423 | n432;
  assign n204 = n201 & n202 & (n86 | n203);
  assign n205 = (n222 | n142) & (n272 | n521);
  assign n206 = (n439 | n496) & (n33 | n470);
  assign n207 = n205 & n206;
  assign n208 = (n86 | n519) & (n100 | n537);
  assign n209 = n53 | n150;
  assign n210 = n674 & n673 & (n272 | n514);
  assign n211 = n566 & n563 & n234 & n605 & n672 & n671;
  assign n212 = n64 & n139 & (n461 | n91);
  assign n213 = n676 & n675 & (n53 | n539);
  assign n214 = n196 & n200 & n204 & n207 & n182 & n189 & n175;
  assign n215 = n670 & n227 & n668 & n667 & n663 & n662 & n666 & n661;
  assign n216 = n208 & n209 & n210 & n211 & n212 & n213 & n214 & n215;
  assign n217 = n258 | n92;
  assign n218 = (n309 | n542) & (n40 | n518);
  assign n219 = ~i_9_ | n451;
  assign n220 = n217 & n218 & (n219 | n38);
  assign n221 = (n86 | n513) & (n462 | n545);
  assign n222 = i_9_ | n425;
  assign n223 = n442 | n466;
  assign n224 = n221 & (n222 | n223);
  assign n225 = n272 | n501;
  assign n226 = n438 | n439;
  assign n227 = n456 | n100;
  assign n228 = n45 & n72 & (n43 | n525);
  assign n229 = n686 & n685 & (n309 | n294);
  assign n230 = n276 & n652 & n684 & n277;
  assign n231 = n224 & n158 & n220 & n44 & n404 & n693 & n692 & n690;
  assign n232 = n225 & n226 & n227 & n176 & n228 & n229 & n230 & n231;
  assign n233 = n434 | n33;
  assign n234 = n462 | n478;
  assign n235 = n674 & (n40 | n536);
  assign n236 = (n258 | n527) & (n222 | n510);
  assign n237 = n33 | n523;
  assign n238 = (n40 | n519) & (n37 | n259);
  assign n239 = n439 | (n339 & n516);
  assign n240 = n682 & n683 & (n100 | n541);
  assign n241 = n233 & n234 & n235 & n236 & n237 & n238 & n239 & n240;
  assign n242 = (n53 | n534) & (n462 | n54);
  assign n243 = n96 | n272;
  assign n244 = n681 & (n86 | n501);
  assign n245 = n43 | n491;
  assign n246 = n46 & n615 & (n91 | n479);
  assign n247 = n679 & n680 & (n436 | n508);
  assign n248 = n242 & n243 & n244 & n245 & n246 & n247;
  assign n249 = n392 & (n40 | n492);
  assign n250 = n678 & n677 & (n33 | n546);
  assign n251 = n442 | n446;
  assign n252 = n249 & n250 & (n53 | n251);
  assign n253 = n272 | n536;
  assign n254 = (n258 | n540) & (n86 | n515);
  assign n255 = n431 | n441;
  assign n256 = n253 & n254 & (n40 | n255);
  assign n257 = (n91 | n520) & (n456 | n43);
  assign n258 = ~i_9_ | n441;
  assign n259 = n420 | n440;
  assign n260 = n257 & (n258 | n259);
  assign n261 = (n222 | n468) & (n258 | n339);
  assign n262 = n420 | n449;
  assign n263 = n261 & (n53 | n262);
  assign n264 = (n37 | n290) & (n454 | n86);
  assign n265 = (n219 | n511) & (n33 | n494);
  assign n266 = n710 & n709 & (n309 | n506);
  assign n267 = n713 & n712 & (n33 | n479);
  assign n268 = n252 & n256 & n260 & n263 & n241 & n248 & n232 & n717;
  assign n269 = n700 & n177 & n699 & n698 & n695 & n694 & n697 & n708;
  assign n270 = n264 & n265 & n266 & n267 & n268 & n269;
  assign n271 = (n100 | n535) & (n439 | n251);
  assign n272 = i_9_ | n449;
  assign n273 = n271 & (n272 | n42);
  assign n274 = n91 | n546;
  assign n275 = n439 | n546;
  assign n276 = n436 | n476;
  assign n277 = n219 | n150;
  assign n278 = n253 & n719 & (n309 | n528);
  assign n279 = n714 & (n91 | n526);
  assign n280 = n321 & (n37 | n438);
  assign n281 = n721 & n720 & (n86 | n41);
  assign n282 = n274 & n275 & n276 & n277 & n278 & n279 & n280 & n281;
  assign n283 = n219 | n478;
  assign n284 = n428 | n436;
  assign n285 = n100 | n521;
  assign n286 = n665 & (n455 | n219);
  assign n287 = n161 & n283 & n263 & n284 & n285 & n286;
  assign n288 = (n40 | n497) & (n37 | n539);
  assign n289 = n718 & (n219 | n486);
  assign n290 = n453 | n460;
  assign n291 = n288 & n289 & (n290 | n91);
  assign n292 = n43 | (n476 & n506);
  assign n293 = n686 & (n53 | n473);
  assign n294 = n423 | n466;
  assign n295 = n292 & n293 & (n272 | n294);
  assign n296 = n219 | n469;
  assign n297 = n100 | n533;
  assign n298 = (n272 | n543) & (n462 | n486);
  assign n299 = n455 | n53;
  assign n300 = n296 & n297 & n298 & n299;
  assign n301 = (n436 | n529) & (n219 | n547);
  assign n302 = n749 & n748 & (n91 | n516);
  assign n303 = n282 & n287 & n291 & n295 & n300 & n252 & n224 & n196;
  assign n304 = n747 & n746 & n745 & n744 & n743 & n742 & n741 & n740;
  assign n305 = n738 & n739 & n730 & n732 & n731 & n737 & n736 & n735;
  assign n306 = n729 & n728 & n727 & n726 & n725 & n724 & n723 & n722;
  assign n307 = n678 & (n219 | n490);
  assign n308 = (n219 | n507) & (n459 | n462);
  assign n309 = i_9_ | n446;
  assign n310 = n419 | n433;
  assign n311 = n307 & n308 & (n309 | n310);
  assign n312 = n53 | n503;
  assign n313 = n710 & n632 & (n309 | n501);
  assign n314 = n753 & n590 & n190 & n78 & n79 & n51;
  assign n315 = n469 | n91;
  assign n316 = n669 & n649 & (n37 | n477);
  assign n317 = n751 & n752 & (n439 | n92);
  assign n318 = n311 & n312 & n313 & n314 & n315 & n234 & n316 & n317;
  assign n319 = n447 | n100;
  assign n320 = n219 | n477;
  assign n321 = n219 | n154;
  assign n322 = (n439 | n461) & (n100 | n530);
  assign n323 = n222 | n472;
  assign n324 = n654 & (n91 | n259);
  assign n325 = (n222 | n537) & (n37 | n482);
  assign n326 = n750 & n738 & (n272 | n484);
  assign n327 = n319 & n320 & n321 & n322 & n323 & n324 & n325 & n326;
  assign n328 = n436 | n492;
  assign n329 = n53 | n489;
  assign n330 = n452 | n100;
  assign n331 = (n465 | n43) & (n272 | n512);
  assign n332 = (n439 | n538) & (n37 | n527);
  assign n333 = n462 | n538;
  assign n334 = (n462 | n520) & (n424 | n219);
  assign n335 = n258 | n490;
  assign n336 = n328 & n329 & n330 & n331 & n332 & n333 & n334 & n335;
  assign n337 = n53 | n520;
  assign n338 = n43 | n203;
  assign n339 = n420 | n425;
  assign n340 = n337 & n338 & (n53 | n339);
  assign n341 = n759 & n758 & (n462 | n527);
  assign n342 = n602 & n757 & (n258 | n479);
  assign n343 = n614 & n756 & (n43 | n497);
  assign n344 = n755 & n754 & (n43 | n294);
  assign n345 = n599 & n274 & n761 & n763 & n762 & n765 & n764 & n766;
  assign n346 = n773 & n621 & n772 & n771;
  assign n347 = n769 & n770 & n552 & n562 & n768 & n767;
  assign n348 = n340 & n300 & n248 & n220 & n327 & n336 & n318 & n777;
  assign n349 = n341 & n342 & n343 & n344 & n345 & n346 & n347 & n348;
  assign n350 = n99 | n272;
  assign n351 = n462 | n103;
  assign n352 = n340 & (n459 | n219);
  assign n353 = (n436 | n468) & (n33 | n467);
  assign n354 = n94 & n582 & (n43 | n541);
  assign n355 = n315 & n782 & (n258 | n511);
  assign n356 = n739 & n780 & (n222 | n491);
  assign n357 = n297 & n350 & n351 & n352 & n353 & n354 & n355 & n356;
  assign n358 = (n436 | n532) & (n91 | n470);
  assign n359 = n40 | n528;
  assign n360 = (n43 | n515) & (n424 | n53);
  assign n361 = n222 | n536;
  assign n362 = n779 & n676 & (n100 | n142);
  assign n363 = n778 & n760 & (n91 | n477);
  assign n364 = n358 & n359 & n360 & n361 & n362 & n363;
  assign n365 = (n222 | n524) & (n436 | n537);
  assign n366 = n100 | n532;
  assign n367 = (n91 | n498) & (n40 | n541);
  assign n368 = (n33 | n154) & (n222 | n541);
  assign n369 = n53 | n502;
  assign n370 = n569 & (n436 | n157);
  assign n371 = n365 & n366 & n367 & n368 & n369 & n370;
  assign n372 = n801 & n800 & (n455 | n462);
  assign n373 = n798 & n797 & (n272 | n530);
  assign n374 = n364 & n371 & n357 & n804 & n88 & n55 & n116 & n803;
  assign n375 = n795 & n794 & (n290 | n219);
  assign n376 = n792 & n791 & (n100 | n493);
  assign n377 = n788 & n789 & n787 & n786 & n785 & n217 & n784 & n783;
  assign n378 = n372 & n373 & n374 & n375 & n376 & n377;
  assign n379 = n462 | (n444 & n534);
  assign n380 = n258 | n507;
  assign n381 = n808 & (n53 | n471);
  assign n382 = n809 & n810 & (n100 | n501);
  assign n383 = n806 & n807 & (n53 | n461);
  assign n384 = n759 & n805 & (n40 | n484);
  assign n385 = n379 & n380 & n381 & n382 & n383 & n384;
  assign n386 = n86 | n514;
  assign n387 = n219 | n496;
  assign n388 = n91 | n482;
  assign n389 = n101 & (n272 | n519);
  assign n390 = n40 | n514;
  assign n391 = n37 | n154;
  assign n392 = n430 | n100;
  assign n393 = n596 & n597 & (n439 | n520);
  assign n394 = n386 & n387 & n388 & n389 & n390 & n391 & n392 & n393;
  assign n395 = (n222 | n447) & (n37 | n339);
  assign n396 = n43 | (n454 & n510);
  assign n397 = n811 & (n37 | n434);
  assign n398 = n813 & (n462 | n546);
  assign n399 = n812 & (n53 | n498);
  assign n400 = n817 & n818 & (n439 | n103);
  assign n401 = n816 & n815 & (n272 | n508);
  assign n402 = n182 & n143 & n260 & n827 & n93 & n828 & n826 & n822;
  assign n403 = n395 & n396 & n397 & n398 & n399 & n400 & n401 & n402;
  assign n404 = n33 | n534;
  assign n405 = (n37 | n502) & (n86 | n524);
  assign n406 = (n100 | n518) & (n222 | n454);
  assign n407 = n318 & n287 & n256 & n200 & n394 & n364 & n273;
  assign n408 = n111 & n606 & n808 & n849 & n848 & n847 & n846 & n845;
  assign n409 = n843 & n564 & n842 & n840 & n832 & n831 & n830 & n836;
  assign n410 = (n86 | n533) & (n439 | n199);
  assign n411 = n438 | n91;
  assign n412 = n858 & n555 & (n43 | n533);
  assign n413 = n721 & n857 & (n100 | n517);
  assign n414 = n781 & n856 & (n462 | n499);
  assign n415 = n855 & n854 & (n309 | n468);
  assign n416 = n852 & n851 & (n33 | n444);
  assign n417 = n132 & n83 & n175 & n868 & n867 & n869 & n866 & n862;
  assign n418 = n410 & n411 & n412 & n413 & n414 & n415 & n416 & n417;
  assign n419 = i_8_ | i_6_ | ~i_7_;
  assign n420 = ~i_5_ | ~i_3_ | i_4_;
  assign n421 = ~i_0_ | ~i_1_ | ~i_2_;
  assign n422 = n420 | n421;
  assign n423 = i_5_ | i_3_ | ~i_4_;
  assign n424 = n421 | n423;
  assign n425 = ~i_0_ | ~i_1_ | i_2_;
  assign n426 = ~i_3_ | ~i_4_ | i_5_;
  assign n427 = ~i_6_ | ~i_7_ | i_8_;
  assign n428 = n426 | n427;
  assign n429 = ~i_6_ | ~i_7_ | ~i_8_;
  assign n430 = n420 | n429;
  assign n431 = ~i_5_ | i_3_ | i_4_;
  assign n432 = i_8_ | i_6_ | i_7_;
  assign n433 = i_5_ | i_3_ | i_4_;
  assign n434 = n425 | n433;
  assign n435 = ~i_2_ | ~i_0_ | i_1_;
  assign n436 = i_9_ | n435;
  assign n437 = i_8_ | ~i_6_ | i_7_;
  assign n438 = n433 | n435;
  assign n439 = ~i_9_ | n437;
  assign n440 = i_2_ | ~i_0_ | i_1_;
  assign n441 = ~i_8_ | ~i_6_ | i_7_;
  assign n442 = ~i_3_ | ~i_4_ | ~i_5_;
  assign n443 = n419 | n442;
  assign n444 = n431 | n440;
  assign n445 = n433 | n440;
  assign n446 = ~i_2_ | i_0_ | ~i_1_;
  assign n447 = n419 | n420;
  assign n448 = n431 | n437;
  assign n449 = i_2_ | i_0_ | ~i_1_;
  assign n450 = i_5_ | ~i_3_ | i_4_;
  assign n451 = ~i_8_ | i_6_ | ~i_7_;
  assign n452 = n450 | n451;
  assign n453 = ~i_5_ | i_3_ | ~i_4_;
  assign n454 = n429 | n453;
  assign n455 = n423 | n449;
  assign n456 = n423 | n441;
  assign n457 = ~i_2_ | i_0_ | i_1_;
  assign n458 = n429 | n431;
  assign n459 = n433 | n457;
  assign n460 = i_2_ | i_0_ | i_1_;
  assign n461 = n450 | n460;
  assign n462 = ~i_9_ | n432;
  assign n463 = n423 | n429;
  assign n464 = n431 | n460;
  assign n465 = n427 | n433;
  assign n466 = ~i_8_ | i_6_ | i_7_;
  assign n467 = n421 | n450;
  assign n468 = n423 | n437;
  assign n469 = n421 | n431;
  assign n470 = n425 | n426;
  assign n471 = n425 | n453;
  assign n472 = n433 | n441;
  assign n473 = n426 | n440;
  assign n474 = n453 | n466;
  assign n475 = n423 | n451;
  assign n476 = n432 | n450;
  assign n477 = n426 | n457;
  assign n478 = n420 | n460;
  assign n479 = n420 | n435;
  assign n480 = n432 | n453;
  assign n481 = n426 | n429;
  assign n482 = n421 | n426;
  assign n483 = n421 | n453;
  assign n484 = n427 | n453;
  assign n485 = n425 | n431;
  assign n486 = n431 | n446;
  assign n487 = n420 | n427;
  assign n488 = n431 | n449;
  assign n489 = n453 | n457;
  assign n490 = n425 | n450;
  assign n491 = n420 | n466;
  assign n492 = n429 | n450;
  assign n493 = n441 | n453;
  assign n494 = n442 | n449;
  assign n495 = n429 | n433;
  assign n496 = n426 | n460;
  assign n497 = n431 | n466;
  assign n498 = n431 | n435;
  assign n499 = n449 | n453;
  assign n500 = n440 | n450;
  assign n501 = n442 | n451;
  assign n502 = n431 | n457;
  assign n503 = n423 | n440;
  assign n504 = n426 | n449;
  assign n505 = n435 | n453;
  assign n506 = n420 | n437;
  assign n507 = n442 | n460;
  assign n508 = n419 | n423;
  assign n509 = n423 | n425;
  assign n510 = n437 | n453;
  assign n511 = n420 | n457;
  assign n512 = n441 | n450;
  assign n513 = n419 | n426;
  assign n514 = n432 | n433;
  assign n515 = n433 | n451;
  assign n516 = n435 | n450;
  assign n517 = n426 | n451;
  assign n518 = n433 | n437;
  assign n519 = n451 | n453;
  assign n520 = n421 | n433;
  assign n521 = n437 | n442;
  assign n522 = n426 | n435;
  assign n523 = n442 | n457;
  assign n524 = n429 | n442;
  assign n525 = n427 | n442;
  assign n526 = n420 | n446;
  assign n527 = n440 | n442;
  assign n528 = n431 | n451;
  assign n529 = n426 | n441;
  assign n530 = n420 | n451;
  assign n531 = n437 | n450;
  assign n532 = n427 | n431;
  assign n533 = n427 | n450;
  assign n534 = n433 | n446;
  assign n535 = n419 | n453;
  assign n536 = n432 | n442;
  assign n537 = n423 | n427;
  assign n538 = n446 | n453;
  assign n539 = n449 | n450;
  assign n540 = n433 | n449;
  assign n541 = n426 | n432;
  assign n542 = n419 | n431;
  assign n543 = n426 | n437;
  assign n544 = n450 | n466;
  assign n545 = n446 | n450;
  assign n546 = n440 | n453;
  assign n547 = n425 | n442;
  assign n548 = n462 | n259;
  assign n549 = n439 | n504;
  assign n550 = n91 | n503;
  assign n551 = (n222 | n493) & (n424 | n33);
  assign n552 = n53 | n479;
  assign n553 = n436 | n493;
  assign n554 = (n222 | n484) & (n33 | n339);
  assign n555 = n456 | n86;
  assign n556 = n315 & n338 & (n462 | n470);
  assign n557 = n323 & n411 & (n33 | n471);
  assign n558 = n40 | n157;
  assign n559 = n91 | n473;
  assign n560 = n558 & n559 & (n309 | n474);
  assign n561 = n53 | n467;
  assign n562 = n157 | n43;
  assign n563 = n309 | n475;
  assign n564 = n272 | n203;
  assign n565 = n428 | n86;
  assign n566 = n33 | n478;
  assign n567 = (n219 | n467) & (n422 | n37);
  assign n568 = (n37 | n424) & (n91 | n483);
  assign n569 = n222 | n430;
  assign n570 = n569 & (n428 | n222);
  assign n571 = (n222 | n99) & (n258 | n485);
  assign n572 = (n436 | n510) & (n434 | n439);
  assign n573 = n99 | n436;
  assign n574 = n33 | n509;
  assign n575 = n572 & n573 & n571 & n233 & n570 & n574 & n568 & n567;
  assign n576 = n96 | n40;
  assign n577 = n576 & n226 & (n40 | n443);
  assign n578 = (n33 | n445) & (n37 | n444);
  assign n579 = n578 & (n439 | n54);
  assign n580 = n309 | (n447 & n448);
  assign n581 = n272 | n454;
  assign n582 = n272 | n452;
  assign n583 = n581 & n582 & (n272 | n493);
  assign n584 = n443 | n272;
  assign n585 = (n33 & n258) | n455;
  assign n586 = (n33 | n511) & (n272 | n456);
  assign n587 = n100 | n42;
  assign n588 = n587 & n330 & (n100 | n203);
  assign n589 = (n459 | n53) & (n100 | n458);
  assign n590 = n463 | n86;
  assign n591 = n290 | n462;
  assign n592 = n590 & n591 & (n448 | n86);
  assign n593 = n258 | n461;
  assign n594 = n40 | n476;
  assign n595 = n91 | n527;
  assign n596 = n458 | n43;
  assign n597 = n439 | n505;
  assign n598 = n40 | n524;
  assign n599 = n40 | n465;
  assign n600 = n91 | n262;
  assign n601 = n258 | n498;
  assign n602 = n436 | n223;
  assign n603 = n40 | n521;
  assign n604 = (n258 | n477) & (n309 | n510);
  assign n605 = n439 | n38;
  assign n606 = n430 | n436;
  assign n607 = n100 | n481;
  assign n608 = n607 & (n100 | n484);
  assign n609 = n100 | n463;
  assign n610 = n549 & n584 & (n43 | n521);
  assign n611 = n422 | n258;
  assign n612 = n222 | n456;
  assign n613 = n612 & (n439 | n485);
  assign n614 = n219 | n520;
  assign n615 = n436 | n518;
  assign n616 = n614 & n615 & (n219 | n470);
  assign n617 = n40 | n508;
  assign n618 = n617 & (n219 | n503);
  assign n619 = n86 | n472;
  assign n620 = n222 | n443;
  assign n621 = n462 | n339;
  assign n622 = (n436 | n42) & (n439 | n522);
  assign n623 = n219 | n259;
  assign n624 = n40 | (n491 & n529);
  assign n625 = n391 & n624 & (n436 | n514);
  assign n626 = (n40 | n458) & (n33 | n500);
  assign n627 = (n272 | n497) & (n258 | n262);
  assign n628 = (n33 | n38) & (n272 | n87);
  assign n629 = (n33 | n502) & (n100 | n468);
  assign n630 = (n33 | n461) & (n91 | n478);
  assign n631 = (n219 | n482) & (n86 | n294);
  assign n632 = n462 | n467;
  assign n633 = n632 & (n43 | n495);
  assign n634 = n222 | n501;
  assign n635 = (n436 | n443) & (n222 | n515);
  assign n636 = (n37 | n479) & (n462 | n92);
  assign n637 = (n40 | n517) & (n37 | n516);
  assign n638 = n309 | (n491 & n497);
  assign n639 = (n272 | n518) & (n37 | n499);
  assign n640 = (n100 | n519) & (n219 | n489);
  assign n641 = n100 | n87;
  assign n642 = n91 | n251;
  assign n643 = (n258 | n464) & (n86 | n535);
  assign n644 = n158 & n161 & n155 & n71 & n35 & n643;
  assign n645 = n436 | n454;
  assign n646 = n43 | n87;
  assign n647 = n272 | n310;
  assign n648 = n86 | n541;
  assign n649 = n439 | n502;
  assign n650 = n43 | (n493 & n513);
  assign n651 = (n258 | n520) & (n43 | n475);
  assign n652 = n53 | n470;
  assign n653 = n652 & (n439 | n470);
  assign n654 = n222 | n532;
  assign n655 = n654 & (n91 | n509);
  assign n656 = (n434 | n91) & (n222 | n528);
  assign n657 = (n436 | n536) & (n222 | n87);
  assign n658 = n436 | n484;
  assign n659 = n658 & (n462 | n516);
  assign n660 = n462 | n154;
  assign n661 = n659 & n660 & n657 & n656 & n655 & n653 & n651 & n650;
  assign n662 = (n40 | n42) & (n436 | n465);
  assign n663 = n40 | (n510 & n537);
  assign n664 = (n37 | n445) & (n40 | n448);
  assign n665 = n258 | n54;
  assign n666 = n665 & n664 & (n309 | n536);
  assign n667 = (n272 | n517) & (n37 | n34);
  assign n668 = (n100 | n529) & (n53 | n523);
  assign n669 = n462 | n199;
  assign n670 = n669 & (n100 | n513);
  assign n671 = (n37 | n503) & (n33 | n527);
  assign n672 = (n219 | n538) & (n444 | n91);
  assign n673 = (n272 | n524) & (n258 | n34);
  assign n674 = n272 | n463;
  assign n675 = (n219 | n526) & (n309 | n157);
  assign n676 = n439 | n507;
  assign n677 = (n439 | n479) & (n258 | n150);
  assign n678 = n309 | n537;
  assign n679 = n436 | n531;
  assign n680 = n430 | n43;
  assign n681 = n309 | n530;
  assign n682 = n272 | n492;
  assign n683 = n309 | n508;
  assign n684 = n219 | n483;
  assign n685 = (n33 | n545) & (n439 | n473);
  assign n686 = n33 | n488;
  assign n687 = n43 | n528;
  assign n688 = n687 & (n33 | n490);
  assign n689 = n53 | n494;
  assign n690 = n689 & n688 & (n53 | n527);
  assign n691 = n462 | n540;
  assign n692 = n691 & n623 & (n272 | n535);
  assign n693 = (n219 | n509) & (n37 | n523);
  assign n694 = (n462 | n509) & (n43 | n518);
  assign n695 = (n40 | n487) & (n53 | n505);
  assign n696 = (n444 | n53) & (n40 | n544);
  assign n697 = n390 & n696 & (n428 | n309);
  assign n698 = (n37 | n538) & (n258 | n545);
  assign n699 = n179 & (n91 | n494);
  assign n700 = (n439 | n262) & (n272 | n41);
  assign n701 = (n91 | n199) & (n258 | n523);
  assign n702 = (n258 | n38) & (n100 | n476);
  assign n703 = n619 & (n86 | n518);
  assign n704 = (n222 | n448) & (n43 | n142);
  assign n705 = (n436 | n530) & (n462 | n522);
  assign n706 = (n436 | n515) & (n219 | n516);
  assign n707 = n706 & (n436 | n310);
  assign n708 = n550 & n60 & n703 & n702 & n701 & n705 & n704 & n707;
  assign n709 = (n309 | n512) & (n53 | n545);
  assign n710 = n40 | n515;
  assign n711 = n351 & (n99 | n86);
  assign n712 = n620 & n711 & (n43 | n543);
  assign n713 = (n272 | n472) & (n91 | n54);
  assign n714 = n309 | n535;
  assign n715 = n714 & (n430 | n40);
  assign n716 = (n219 | n494) & (n33 | n540);
  assign n717 = n207 & n123 & n104 & n39 & n716 & n715;
  assign n718 = (n40 | n506) & (n258 | n470);
  assign n719 = (n272 | n542) & (n53 | n499);
  assign n720 = (n436 | n517) & (n43 | n544);
  assign n721 = n53 | n477;
  assign n722 = (n53 | n482) & (n439 | n150);
  assign n723 = (n439 | n483) & (n422 | n219);
  assign n724 = (n43 | n508) & (n424 | n258);
  assign n725 = (n33 & n258) | n547;
  assign n726 = n222 | (n487 & n543);
  assign n727 = (n33 | n516) & (n439 | n490);
  assign n728 = n598 & (n436 | n528);
  assign n729 = n595 & (n462 | n500);
  assign n730 = (n40 | n535) & (n37 | n546);
  assign n731 = n186 & (n309 | n142);
  assign n732 = n309 | (n255 & n519);
  assign n733 = (n430 | n272) & (n309 | n514);
  assign n734 = n100 | n524;
  assign n735 = n734 & n733 & (n272 | n475);
  assign n736 = (n258 | n489) & (n100 | n536);
  assign n737 = (n258 | n103) & (n462 | n38);
  assign n738 = n444 | n219;
  assign n739 = n462 | n503;
  assign n740 = n386 & (n258 | n160);
  assign n741 = (n422 | n33) & (n43 | n524);
  assign n742 = (n222 | n521) & (n448 | n43);
  assign n743 = n436 | (n495 & n512);
  assign n744 = n681 & (n37 | n494);
  assign n745 = (n219 | n523) & (n272 | n541);
  assign n746 = (n37 | n496) & (n258 | n199);
  assign n747 = n612 & (n434 | n258);
  assign n748 = (n219 | n502) & (n272 | n537);
  assign n749 = n219 | n522;
  assign n750 = n219 | n262;
  assign n751 = (n222 | n506) & (n43 | n472);
  assign n752 = n595 & n194 & (n436 | n448);
  assign n753 = n462 | n471;
  assign n754 = (n258 | n483) & (n43 | n531);
  assign n755 = n424 | n91;
  assign n756 = n222 | (n529 & n530);
  assign n757 = (n434 | n219) & (n222 | n542);
  assign n758 = (n37 | n498) & (n436 | n294);
  assign n759 = n258 | n546;
  assign n760 = n40 | n472;
  assign n761 = n760 & (n445 | n258);
  assign n762 = (n309 | n525) & (n439 | n445);
  assign n763 = (n309 | n493) & (n462 | n251);
  assign n764 = n118 & (n219 | n534);
  assign n765 = n272 | (n157 & n506);
  assign n766 = n600 & n607 & (n33 | n539);
  assign n767 = (n86 | n536) & (n37 | n511);
  assign n768 = (n219 | n160) & (n86 | n517);
  assign n769 = n222 | n519;
  assign n770 = n222 | n525;
  assign n771 = n40 | (n468 & n543);
  assign n772 = (n91 | n486) & (n33 | n526);
  assign n773 = n100 | (n495 & n544);
  assign n774 = (n436 | n542) & (n222 | n517);
  assign n775 = (n439 | n34) & (n40 | n463);
  assign n776 = n258 | n534;
  assign n777 = n189 & n147 & n77 & n776 & n775 & n774;
  assign n778 = n309 | n476;
  assign n779 = n436 | n519;
  assign n780 = n680 & n652 & (n33 | n483);
  assign n781 = n439 | n499;
  assign n782 = n781 & n734 & (n37 | n486);
  assign n783 = (n422 | n53) & (n43 | n517);
  assign n784 = (n222 | n452) & (n258 | n469);
  assign n785 = (n222 | n535) & (n462 | n490);
  assign n786 = (n436 | n475) & (n91 | n522);
  assign n787 = (n438 | n219) & (n33 | n498);
  assign n788 = (n219 | n546) & (n37 | n500);
  assign n789 = n445 | n91;
  assign n790 = (n447 | n272) & (n37 | n504);
  assign n791 = n184 & n790 & (n40 | n87);
  assign n792 = (n53 & n258) | n488;
  assign n793 = (n100 | n310) & (n91 | n502);
  assign n794 = n793 & (n86 | n223);
  assign n795 = n86 | (n491 & n529);
  assign n796 = n558 & (n86 | n537);
  assign n797 = n769 & n796 & (n43 | n542);
  assign n798 = n753 & (n258 | n516);
  assign n799 = (n258 | n526) & (n100 | n512);
  assign n800 = n691 & n799 & (n272 | n531);
  assign n801 = (n272 | n491) & (n33 | n504);
  assign n802 = (n86 | n310) & (n37 | n199);
  assign n803 = n44 & n802 & (n439 | n477);
  assign n804 = n241 & n204 & n282;
  assign n805 = n658 & n755 & (n91 | n500);
  assign n806 = (n459 | n91) & (n53 | n504);
  assign n807 = n57 & (n219 | n471);
  assign n808 = n422 | n439;
  assign n809 = n749 & (n222 | n465);
  assign n810 = (n428 | n43) & (n462 | n150);
  assign n811 = (n37 | n485) & (n222 | n533);
  assign n812 = n436 | (n463 & n524);
  assign n813 = n40 | (n142 & n530);
  assign n814 = (n445 | n462) & (n444 | n258);
  assign n815 = n814 & (n443 | n309);
  assign n816 = (n272 | n481) & (n309 | n529);
  assign n817 = (n258 | n478) & (n53 | n511);
  assign n818 = n68 & n62 & (n439 | n160);
  assign n819 = (n467 | n91) & (n462 | n482);
  assign n820 = n687 & n819 & (n439 | n509);
  assign n821 = (n33 | n473) & (n53 | n516);
  assign n822 = n821 & n820 & (n40 | n531);
  assign n823 = n91 | n499;
  assign n824 = n823 & n689 & (n53 | n540);
  assign n825 = (n436 | n543) & (n86 | n495);
  assign n826 = n825 & n824 & (n258 | n505);
  assign n827 = (n42 | n86) & (n428 | n272);
  assign n828 = n394 & n357 & n385 & n311 & n295 & n336;
  assign n829 = (n43 | n514) & (n462 | n483);
  assign n830 = n684 & n829 & (n443 | n43);
  assign n831 = (n91 | n490) & (n222 | n41);
  assign n832 = (n436 | n501) & (n462 | n485);
  assign n833 = (n436 | n41) & (n33 | n522);
  assign n834 = n645 & n833 & (n438 | n258);
  assign n835 = n603 & (n40 | n474);
  assign n836 = n835 & n834 & (n309 | n521);
  assign n837 = (n219 | n499) & (n272 | n142);
  assign n838 = n683 & n837 & (n462 | n262);
  assign n839 = (n272 | n458) & (n455 | n91);
  assign n840 = n839 & n838 & (n439 | n488);
  assign n841 = n647 & (n100 | n223);
  assign n842 = n609 & n841 & (n439 | n511);
  assign n843 = n33 | (n459 & n464);
  assign n844 = (n436 | n506) & (n53 | n490);
  assign n845 = n565 & n844 & (n43 | n41);
  assign n846 = (n219 | n251) & (n91 | n505);
  assign n847 = n37 | (n54 & n251);
  assign n848 = (n439 | n540) & (n430 | n309);
  assign n849 = n611 & (n462 | n464);
  assign n850 = (n436 | n535) & (n43 | n487);
  assign n851 = n275 & n850 & (n40 | n452);
  assign n852 = n617 & (n40 | n475);
  assign n853 = (n96 | n309) & (n40 | n310);
  assign n854 = n853 & (n309 | n492);
  assign n855 = (n258 | n538) & (n309 | n544);
  assign n856 = (n219 | n504) & (n462 | n494);
  assign n857 = n37 | n455;
  assign n858 = n43 | n536;
  assign n859 = (n37 & n53) | n547;
  assign n860 = n779 & n859 & (n222 | n508);
  assign n861 = n53 | (n154 & n259);
  assign n862 = n861 & n860 & (n40 | n512);
  assign n863 = (n53 | n538) & (n439 | n500);
  assign n864 = n863 & (n100 | n543);
  assign n865 = (n462 | n489) & (n100 | n510);
  assign n866 = n865 & n864 & (n448 | n100);
  assign n867 = (n436 | n481) & (n462 | n34);
  assign n868 = (n436 | n474) & (n258 | n494);
  assign n869 = n385 & n371 & n273 & n291 & n232 & n327;
endmodule


