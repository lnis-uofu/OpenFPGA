*****************************
*     FPGA SPICE Netlist    *
* Description: Connection Block Y-channel  [1][1] in FPGA *
*    Author: Xifan TANG     *
* Organization: EPFL/IC/LSI *
* Date: Thu Nov 15 14:26:08 2018
 *
*****************************
.subckt cby[1][1] 
+ chany[1][1]_midout[0] 
+ chany[1][1]_midout[1] 
+ chany[1][1]_midout[2] 
+ chany[1][1]_midout[3] 
+ chany[1][1]_midout[4] 
+ chany[1][1]_midout[5] 
+ chany[1][1]_midout[6] 
+ chany[1][1]_midout[7] 
+ chany[1][1]_midout[8] 
+ chany[1][1]_midout[9] 
+ chany[1][1]_midout[10] 
+ chany[1][1]_midout[11] 
+ chany[1][1]_midout[12] 
+ chany[1][1]_midout[13] 
+ chany[1][1]_midout[14] 
+ chany[1][1]_midout[15] 
+ chany[1][1]_midout[16] 
+ chany[1][1]_midout[17] 
+ chany[1][1]_midout[18] 
+ chany[1][1]_midout[19] 
+ chany[1][1]_midout[20] 
+ chany[1][1]_midout[21] 
+ chany[1][1]_midout[22] 
+ chany[1][1]_midout[23] 
+ chany[1][1]_midout[24] 
+ chany[1][1]_midout[25] 
+ chany[1][1]_midout[26] 
+ chany[1][1]_midout[27] 
+ chany[1][1]_midout[28] 
+ chany[1][1]_midout[29] 
+ chany[1][1]_midout[30] 
+ chany[1][1]_midout[31] 
+ chany[1][1]_midout[32] 
+ chany[1][1]_midout[33] 
+ chany[1][1]_midout[34] 
+ chany[1][1]_midout[35] 
+ chany[1][1]_midout[36] 
+ chany[1][1]_midout[37] 
+ chany[1][1]_midout[38] 
+ chany[1][1]_midout[39] 
+ chany[1][1]_midout[40] 
+ chany[1][1]_midout[41] 
+ chany[1][1]_midout[42] 
+ chany[1][1]_midout[43] 
+ chany[1][1]_midout[44] 
+ chany[1][1]_midout[45] 
+ chany[1][1]_midout[46] 
+ chany[1][1]_midout[47] 
+ chany[1][1]_midout[48] 
+ chany[1][1]_midout[49] 
+ chany[1][1]_midout[50] 
+ chany[1][1]_midout[51] 
+ chany[1][1]_midout[52] 
+ chany[1][1]_midout[53] 
+ chany[1][1]_midout[54] 
+ chany[1][1]_midout[55] 
+ chany[1][1]_midout[56] 
+ chany[1][1]_midout[57] 
+ chany[1][1]_midout[58] 
+ chany[1][1]_midout[59] 
+ chany[1][1]_midout[60] 
+ chany[1][1]_midout[61] 
+ chany[1][1]_midout[62] 
+ chany[1][1]_midout[63] 
+ chany[1][1]_midout[64] 
+ chany[1][1]_midout[65] 
+ chany[1][1]_midout[66] 
+ chany[1][1]_midout[67] 
+ chany[1][1]_midout[68] 
+ chany[1][1]_midout[69] 
+ chany[1][1]_midout[70] 
+ chany[1][1]_midout[71] 
+ chany[1][1]_midout[72] 
+ chany[1][1]_midout[73] 
+ chany[1][1]_midout[74] 
+ chany[1][1]_midout[75] 
+ chany[1][1]_midout[76] 
+ chany[1][1]_midout[77] 
+ chany[1][1]_midout[78] 
+ chany[1][1]_midout[79] 
+ chany[1][1]_midout[80] 
+ chany[1][1]_midout[81] 
+ chany[1][1]_midout[82] 
+ chany[1][1]_midout[83] 
+ chany[1][1]_midout[84] 
+ chany[1][1]_midout[85] 
+ chany[1][1]_midout[86] 
+ chany[1][1]_midout[87] 
+ chany[1][1]_midout[88] 
+ chany[1][1]_midout[89] 
+ chany[1][1]_midout[90] 
+ chany[1][1]_midout[91] 
+ chany[1][1]_midout[92] 
+ chany[1][1]_midout[93] 
+ chany[1][1]_midout[94] 
+ chany[1][1]_midout[95] 
+ chany[1][1]_midout[96] 
+ chany[1][1]_midout[97] 
+ chany[1][1]_midout[98] 
+ chany[1][1]_midout[99] 
+ grid[2][1]_pin[0][3][0] 
+ grid[2][1]_pin[0][3][2] 
+ grid[2][1]_pin[0][3][4] 
+ grid[2][1]_pin[0][3][6] 
+ grid[2][1]_pin[0][3][8] 
+ grid[2][1]_pin[0][3][10] 
+ grid[2][1]_pin[0][3][12] 
+ grid[2][1]_pin[0][3][14] 
+ grid[1][1]_pin[0][1][1] 
+ grid[1][1]_pin[0][1][5] 
+ grid[1][1]_pin[0][1][9] 
+ grid[1][1]_pin[0][1][13] 
+ grid[1][1]_pin[0][1][17] 
+ grid[1][1]_pin[0][1][21] 
+ grid[1][1]_pin[0][1][25] 
+ grid[1][1]_pin[0][1][29] 
+ grid[1][1]_pin[0][1][33] 
+ grid[1][1]_pin[0][1][37] 
+ svdd sgnd
Xmux_2level_tapbuf_size16[54] chany[1][1]_midout[6] chany[1][1]_midout[7] chany[1][1]_midout[10] chany[1][1]_midout[11] chany[1][1]_midout[24] chany[1][1]_midout[25] chany[1][1]_midout[36] chany[1][1]_midout[37] chany[1][1]_midout[48] chany[1][1]_midout[49] chany[1][1]_midout[60] chany[1][1]_midout[61] chany[1][1]_midout[76] chany[1][1]_midout[77] chany[1][1]_midout[88] chany[1][1]_midout[89] grid[2][1]_pin[0][3][0] sram[2514]->outb sram[2514]->out sram[2515]->out sram[2515]->outb sram[2516]->out sram[2516]->outb sram[2517]->out sram[2517]->outb sram[2518]->outb sram[2518]->out sram[2519]->out sram[2519]->outb sram[2520]->out sram[2520]->outb sram[2521]->out sram[2521]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[54], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2514] sram->in sram[2514]->out sram[2514]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2514]->out) 0
.nodeset V(sram[2514]->outb) vsp
Xsram[2515] sram->in sram[2515]->out sram[2515]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2515]->out) 0
.nodeset V(sram[2515]->outb) vsp
Xsram[2516] sram->in sram[2516]->out sram[2516]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2516]->out) 0
.nodeset V(sram[2516]->outb) vsp
Xsram[2517] sram->in sram[2517]->out sram[2517]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2517]->out) 0
.nodeset V(sram[2517]->outb) vsp
Xsram[2518] sram->in sram[2518]->out sram[2518]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2518]->out) 0
.nodeset V(sram[2518]->outb) vsp
Xsram[2519] sram->in sram[2519]->out sram[2519]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2519]->out) 0
.nodeset V(sram[2519]->outb) vsp
Xsram[2520] sram->in sram[2520]->out sram[2520]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2520]->out) 0
.nodeset V(sram[2520]->outb) vsp
Xsram[2521] sram->in sram[2521]->out sram[2521]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2521]->out) 0
.nodeset V(sram[2521]->outb) vsp
Xmux_2level_tapbuf_size16[55] chany[1][1]_midout[0] chany[1][1]_midout[1] chany[1][1]_midout[12] chany[1][1]_midout[13] chany[1][1]_midout[24] chany[1][1]_midout[25] chany[1][1]_midout[42] chany[1][1]_midout[43] chany[1][1]_midout[54] chany[1][1]_midout[55] chany[1][1]_midout[66] chany[1][1]_midout[67] chany[1][1]_midout[76] chany[1][1]_midout[77] chany[1][1]_midout[90] chany[1][1]_midout[91] grid[2][1]_pin[0][3][2] sram[2522]->outb sram[2522]->out sram[2523]->out sram[2523]->outb sram[2524]->out sram[2524]->outb sram[2525]->out sram[2525]->outb sram[2526]->outb sram[2526]->out sram[2527]->out sram[2527]->outb sram[2528]->out sram[2528]->outb sram[2529]->out sram[2529]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[55], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2522] sram->in sram[2522]->out sram[2522]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2522]->out) 0
.nodeset V(sram[2522]->outb) vsp
Xsram[2523] sram->in sram[2523]->out sram[2523]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2523]->out) 0
.nodeset V(sram[2523]->outb) vsp
Xsram[2524] sram->in sram[2524]->out sram[2524]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2524]->out) 0
.nodeset V(sram[2524]->outb) vsp
Xsram[2525] sram->in sram[2525]->out sram[2525]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2525]->out) 0
.nodeset V(sram[2525]->outb) vsp
Xsram[2526] sram->in sram[2526]->out sram[2526]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2526]->out) 0
.nodeset V(sram[2526]->outb) vsp
Xsram[2527] sram->in sram[2527]->out sram[2527]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2527]->out) 0
.nodeset V(sram[2527]->outb) vsp
Xsram[2528] sram->in sram[2528]->out sram[2528]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2528]->out) 0
.nodeset V(sram[2528]->outb) vsp
Xsram[2529] sram->in sram[2529]->out sram[2529]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2529]->out) 0
.nodeset V(sram[2529]->outb) vsp
Xmux_2level_tapbuf_size16[56] chany[1][1]_midout[2] chany[1][1]_midout[3] chany[1][1]_midout[22] chany[1][1]_midout[23] chany[1][1]_midout[26] chany[1][1]_midout[27] chany[1][1]_midout[42] chany[1][1]_midout[43] chany[1][1]_midout[52] chany[1][1]_midout[53] chany[1][1]_midout[64] chany[1][1]_midout[65] chany[1][1]_midout[78] chany[1][1]_midout[79] chany[1][1]_midout[90] chany[1][1]_midout[91] grid[2][1]_pin[0][3][4] sram[2530]->outb sram[2530]->out sram[2531]->out sram[2531]->outb sram[2532]->out sram[2532]->outb sram[2533]->out sram[2533]->outb sram[2534]->outb sram[2534]->out sram[2535]->out sram[2535]->outb sram[2536]->out sram[2536]->outb sram[2537]->out sram[2537]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[56], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2530] sram->in sram[2530]->out sram[2530]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2530]->out) 0
.nodeset V(sram[2530]->outb) vsp
Xsram[2531] sram->in sram[2531]->out sram[2531]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2531]->out) 0
.nodeset V(sram[2531]->outb) vsp
Xsram[2532] sram->in sram[2532]->out sram[2532]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2532]->out) 0
.nodeset V(sram[2532]->outb) vsp
Xsram[2533] sram->in sram[2533]->out sram[2533]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2533]->out) 0
.nodeset V(sram[2533]->outb) vsp
Xsram[2534] sram->in sram[2534]->out sram[2534]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2534]->out) 0
.nodeset V(sram[2534]->outb) vsp
Xsram[2535] sram->in sram[2535]->out sram[2535]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2535]->out) 0
.nodeset V(sram[2535]->outb) vsp
Xsram[2536] sram->in sram[2536]->out sram[2536]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2536]->out) 0
.nodeset V(sram[2536]->outb) vsp
Xsram[2537] sram->in sram[2537]->out sram[2537]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2537]->out) 0
.nodeset V(sram[2537]->outb) vsp
Xmux_2level_tapbuf_size16[57] chany[1][1]_midout[2] chany[1][1]_midout[3] chany[1][1]_midout[16] chany[1][1]_midout[17] chany[1][1]_midout[28] chany[1][1]_midout[29] chany[1][1]_midout[40] chany[1][1]_midout[41] chany[1][1]_midout[52] chany[1][1]_midout[53] chany[1][1]_midout[68] chany[1][1]_midout[69] chany[1][1]_midout[80] chany[1][1]_midout[81] chany[1][1]_midout[92] chany[1][1]_midout[93] grid[2][1]_pin[0][3][6] sram[2538]->outb sram[2538]->out sram[2539]->out sram[2539]->outb sram[2540]->out sram[2540]->outb sram[2541]->out sram[2541]->outb sram[2542]->outb sram[2542]->out sram[2543]->out sram[2543]->outb sram[2544]->out sram[2544]->outb sram[2545]->out sram[2545]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[57], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2538] sram->in sram[2538]->out sram[2538]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2538]->out) 0
.nodeset V(sram[2538]->outb) vsp
Xsram[2539] sram->in sram[2539]->out sram[2539]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2539]->out) 0
.nodeset V(sram[2539]->outb) vsp
Xsram[2540] sram->in sram[2540]->out sram[2540]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2540]->out) 0
.nodeset V(sram[2540]->outb) vsp
Xsram[2541] sram->in sram[2541]->out sram[2541]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2541]->out) 0
.nodeset V(sram[2541]->outb) vsp
Xsram[2542] sram->in sram[2542]->out sram[2542]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2542]->out) 0
.nodeset V(sram[2542]->outb) vsp
Xsram[2543] sram->in sram[2543]->out sram[2543]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2543]->out) 0
.nodeset V(sram[2543]->outb) vsp
Xsram[2544] sram->in sram[2544]->out sram[2544]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2544]->out) 0
.nodeset V(sram[2544]->outb) vsp
Xsram[2545] sram->in sram[2545]->out sram[2545]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2545]->out) 0
.nodeset V(sram[2545]->outb) vsp
Xmux_2level_tapbuf_size16[58] chany[1][1]_midout[4] chany[1][1]_midout[5] chany[1][1]_midout[16] chany[1][1]_midout[17] chany[1][1]_midout[38] chany[1][1]_midout[39] chany[1][1]_midout[46] chany[1][1]_midout[47] chany[1][1]_midout[58] chany[1][1]_midout[59] chany[1][1]_midout[68] chany[1][1]_midout[69] chany[1][1]_midout[82] chany[1][1]_midout[83] chany[1][1]_midout[94] chany[1][1]_midout[95] grid[2][1]_pin[0][3][8] sram[2546]->outb sram[2546]->out sram[2547]->out sram[2547]->outb sram[2548]->out sram[2548]->outb sram[2549]->out sram[2549]->outb sram[2550]->outb sram[2550]->out sram[2551]->out sram[2551]->outb sram[2552]->out sram[2552]->outb sram[2553]->out sram[2553]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[58], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2546] sram->in sram[2546]->out sram[2546]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2546]->out) 0
.nodeset V(sram[2546]->outb) vsp
Xsram[2547] sram->in sram[2547]->out sram[2547]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2547]->out) 0
.nodeset V(sram[2547]->outb) vsp
Xsram[2548] sram->in sram[2548]->out sram[2548]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2548]->out) 0
.nodeset V(sram[2548]->outb) vsp
Xsram[2549] sram->in sram[2549]->out sram[2549]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2549]->out) 0
.nodeset V(sram[2549]->outb) vsp
Xsram[2550] sram->in sram[2550]->out sram[2550]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2550]->out) 0
.nodeset V(sram[2550]->outb) vsp
Xsram[2551] sram->in sram[2551]->out sram[2551]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2551]->out) 0
.nodeset V(sram[2551]->outb) vsp
Xsram[2552] sram->in sram[2552]->out sram[2552]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2552]->out) 0
.nodeset V(sram[2552]->outb) vsp
Xsram[2553] sram->in sram[2553]->out sram[2553]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2553]->out) 0
.nodeset V(sram[2553]->outb) vsp
Xmux_2level_tapbuf_size16[59] chany[1][1]_midout[14] chany[1][1]_midout[15] chany[1][1]_midout[18] chany[1][1]_midout[19] chany[1][1]_midout[38] chany[1][1]_midout[39] chany[1][1]_midout[44] chany[1][1]_midout[45] chany[1][1]_midout[56] chany[1][1]_midout[57] chany[1][1]_midout[70] chany[1][1]_midout[71] chany[1][1]_midout[82] chany[1][1]_midout[83] chany[1][1]_midout[96] chany[1][1]_midout[97] grid[2][1]_pin[0][3][10] sram[2554]->outb sram[2554]->out sram[2555]->out sram[2555]->outb sram[2556]->out sram[2556]->outb sram[2557]->out sram[2557]->outb sram[2558]->outb sram[2558]->out sram[2559]->out sram[2559]->outb sram[2560]->out sram[2560]->outb sram[2561]->out sram[2561]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[59], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2554] sram->in sram[2554]->out sram[2554]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2554]->out) 0
.nodeset V(sram[2554]->outb) vsp
Xsram[2555] sram->in sram[2555]->out sram[2555]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2555]->out) 0
.nodeset V(sram[2555]->outb) vsp
Xsram[2556] sram->in sram[2556]->out sram[2556]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2556]->out) 0
.nodeset V(sram[2556]->outb) vsp
Xsram[2557] sram->in sram[2557]->out sram[2557]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2557]->out) 0
.nodeset V(sram[2557]->outb) vsp
Xsram[2558] sram->in sram[2558]->out sram[2558]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2558]->out) 0
.nodeset V(sram[2558]->outb) vsp
Xsram[2559] sram->in sram[2559]->out sram[2559]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2559]->out) 0
.nodeset V(sram[2559]->outb) vsp
Xsram[2560] sram->in sram[2560]->out sram[2560]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2560]->out) 0
.nodeset V(sram[2560]->outb) vsp
Xsram[2561] sram->in sram[2561]->out sram[2561]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2561]->out) 0
.nodeset V(sram[2561]->outb) vsp
Xmux_2level_tapbuf_size16[60] chany[1][1]_midout[8] chany[1][1]_midout[9] chany[1][1]_midout[20] chany[1][1]_midout[21] chany[1][1]_midout[32] chany[1][1]_midout[33] chany[1][1]_midout[50] chany[1][1]_midout[51] chany[1][1]_midout[62] chany[1][1]_midout[63] chany[1][1]_midout[72] chany[1][1]_midout[73] chany[1][1]_midout[84] chany[1][1]_midout[85] chany[1][1]_midout[98] chany[1][1]_midout[99] grid[2][1]_pin[0][3][12] sram[2562]->outb sram[2562]->out sram[2563]->out sram[2563]->outb sram[2564]->out sram[2564]->outb sram[2565]->out sram[2565]->outb sram[2566]->outb sram[2566]->out sram[2567]->out sram[2567]->outb sram[2568]->out sram[2568]->outb sram[2569]->out sram[2569]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[60], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2562] sram->in sram[2562]->out sram[2562]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2562]->out) 0
.nodeset V(sram[2562]->outb) vsp
Xsram[2563] sram->in sram[2563]->out sram[2563]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2563]->out) 0
.nodeset V(sram[2563]->outb) vsp
Xsram[2564] sram->in sram[2564]->out sram[2564]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2564]->out) 0
.nodeset V(sram[2564]->outb) vsp
Xsram[2565] sram->in sram[2565]->out sram[2565]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2565]->out) 0
.nodeset V(sram[2565]->outb) vsp
Xsram[2566] sram->in sram[2566]->out sram[2566]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2566]->out) 0
.nodeset V(sram[2566]->outb) vsp
Xsram[2567] sram->in sram[2567]->out sram[2567]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2567]->out) 0
.nodeset V(sram[2567]->outb) vsp
Xsram[2568] sram->in sram[2568]->out sram[2568]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2568]->out) 0
.nodeset V(sram[2568]->outb) vsp
Xsram[2569] sram->in sram[2569]->out sram[2569]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2569]->out) 0
.nodeset V(sram[2569]->outb) vsp
Xmux_2level_tapbuf_size16[61] chany[1][1]_midout[10] chany[1][1]_midout[11] chany[1][1]_midout[30] chany[1][1]_midout[31] chany[1][1]_midout[34] chany[1][1]_midout[35] chany[1][1]_midout[50] chany[1][1]_midout[51] chany[1][1]_midout[60] chany[1][1]_midout[61] chany[1][1]_midout[74] chany[1][1]_midout[75] chany[1][1]_midout[86] chany[1][1]_midout[87] chany[1][1]_midout[98] chany[1][1]_midout[99] grid[2][1]_pin[0][3][14] sram[2570]->outb sram[2570]->out sram[2571]->out sram[2571]->outb sram[2572]->out sram[2572]->outb sram[2573]->out sram[2573]->outb sram[2574]->outb sram[2574]->out sram[2575]->out sram[2575]->outb sram[2576]->out sram[2576]->outb sram[2577]->out sram[2577]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[61], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2570] sram->in sram[2570]->out sram[2570]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2570]->out) 0
.nodeset V(sram[2570]->outb) vsp
Xsram[2571] sram->in sram[2571]->out sram[2571]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2571]->out) 0
.nodeset V(sram[2571]->outb) vsp
Xsram[2572] sram->in sram[2572]->out sram[2572]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2572]->out) 0
.nodeset V(sram[2572]->outb) vsp
Xsram[2573] sram->in sram[2573]->out sram[2573]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2573]->out) 0
.nodeset V(sram[2573]->outb) vsp
Xsram[2574] sram->in sram[2574]->out sram[2574]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2574]->out) 0
.nodeset V(sram[2574]->outb) vsp
Xsram[2575] sram->in sram[2575]->out sram[2575]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2575]->out) 0
.nodeset V(sram[2575]->outb) vsp
Xsram[2576] sram->in sram[2576]->out sram[2576]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2576]->out) 0
.nodeset V(sram[2576]->outb) vsp
Xsram[2577] sram->in sram[2577]->out sram[2577]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2577]->out) 0
.nodeset V(sram[2577]->outb) vsp
Xmux_2level_tapbuf_size16[62] chany[1][1]_midout[6] chany[1][1]_midout[7] chany[1][1]_midout[10] chany[1][1]_midout[11] chany[1][1]_midout[30] chany[1][1]_midout[31] chany[1][1]_midout[34] chany[1][1]_midout[35] chany[1][1]_midout[48] chany[1][1]_midout[49] chany[1][1]_midout[60] chany[1][1]_midout[61] chany[1][1]_midout[74] chany[1][1]_midout[75] chany[1][1]_midout[86] chany[1][1]_midout[87] grid[1][1]_pin[0][1][1] sram[2578]->outb sram[2578]->out sram[2579]->out sram[2579]->outb sram[2580]->out sram[2580]->outb sram[2581]->out sram[2581]->outb sram[2582]->outb sram[2582]->out sram[2583]->out sram[2583]->outb sram[2584]->out sram[2584]->outb sram[2585]->out sram[2585]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[62], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2578] sram->in sram[2578]->out sram[2578]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2578]->out) 0
.nodeset V(sram[2578]->outb) vsp
Xsram[2579] sram->in sram[2579]->out sram[2579]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2579]->out) 0
.nodeset V(sram[2579]->outb) vsp
Xsram[2580] sram->in sram[2580]->out sram[2580]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2580]->out) 0
.nodeset V(sram[2580]->outb) vsp
Xsram[2581] sram->in sram[2581]->out sram[2581]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2581]->out) 0
.nodeset V(sram[2581]->outb) vsp
Xsram[2582] sram->in sram[2582]->out sram[2582]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2582]->out) 0
.nodeset V(sram[2582]->outb) vsp
Xsram[2583] sram->in sram[2583]->out sram[2583]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2583]->out) 0
.nodeset V(sram[2583]->outb) vsp
Xsram[2584] sram->in sram[2584]->out sram[2584]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2584]->out) 0
.nodeset V(sram[2584]->outb) vsp
Xsram[2585] sram->in sram[2585]->out sram[2585]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2585]->out) 0
.nodeset V(sram[2585]->outb) vsp
Xmux_2level_tapbuf_size16[63] chany[1][1]_midout[6] chany[1][1]_midout[7] chany[1][1]_midout[12] chany[1][1]_midout[13] chany[1][1]_midout[24] chany[1][1]_midout[25] chany[1][1]_midout[36] chany[1][1]_midout[37] chany[1][1]_midout[48] chany[1][1]_midout[49] chany[1][1]_midout[66] chany[1][1]_midout[67] chany[1][1]_midout[76] chany[1][1]_midout[77] chany[1][1]_midout[88] chany[1][1]_midout[89] grid[1][1]_pin[0][1][5] sram[2586]->outb sram[2586]->out sram[2587]->out sram[2587]->outb sram[2588]->out sram[2588]->outb sram[2589]->out sram[2589]->outb sram[2590]->outb sram[2590]->out sram[2591]->out sram[2591]->outb sram[2592]->out sram[2592]->outb sram[2593]->out sram[2593]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[63], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2586] sram->in sram[2586]->out sram[2586]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2586]->out) 0
.nodeset V(sram[2586]->outb) vsp
Xsram[2587] sram->in sram[2587]->out sram[2587]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2587]->out) 0
.nodeset V(sram[2587]->outb) vsp
Xsram[2588] sram->in sram[2588]->out sram[2588]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2588]->out) 0
.nodeset V(sram[2588]->outb) vsp
Xsram[2589] sram->in sram[2589]->out sram[2589]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2589]->out) 0
.nodeset V(sram[2589]->outb) vsp
Xsram[2590] sram->in sram[2590]->out sram[2590]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2590]->out) 0
.nodeset V(sram[2590]->outb) vsp
Xsram[2591] sram->in sram[2591]->out sram[2591]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2591]->out) 0
.nodeset V(sram[2591]->outb) vsp
Xsram[2592] sram->in sram[2592]->out sram[2592]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2592]->out) 0
.nodeset V(sram[2592]->outb) vsp
Xsram[2593] sram->in sram[2593]->out sram[2593]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2593]->out) 0
.nodeset V(sram[2593]->outb) vsp
Xmux_2level_tapbuf_size16[64] chany[1][1]_midout[0] chany[1][1]_midout[1] chany[1][1]_midout[12] chany[1][1]_midout[13] chany[1][1]_midout[24] chany[1][1]_midout[25] chany[1][1]_midout[42] chany[1][1]_midout[43] chany[1][1]_midout[54] chany[1][1]_midout[55] chany[1][1]_midout[66] chany[1][1]_midout[67] chany[1][1]_midout[76] chany[1][1]_midout[77] chany[1][1]_midout[90] chany[1][1]_midout[91] grid[1][1]_pin[0][1][9] sram[2594]->outb sram[2594]->out sram[2595]->out sram[2595]->outb sram[2596]->out sram[2596]->outb sram[2597]->out sram[2597]->outb sram[2598]->outb sram[2598]->out sram[2599]->out sram[2599]->outb sram[2600]->out sram[2600]->outb sram[2601]->out sram[2601]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[64], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2594] sram->in sram[2594]->out sram[2594]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2594]->out) 0
.nodeset V(sram[2594]->outb) vsp
Xsram[2595] sram->in sram[2595]->out sram[2595]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2595]->out) 0
.nodeset V(sram[2595]->outb) vsp
Xsram[2596] sram->in sram[2596]->out sram[2596]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2596]->out) 0
.nodeset V(sram[2596]->outb) vsp
Xsram[2597] sram->in sram[2597]->out sram[2597]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2597]->out) 0
.nodeset V(sram[2597]->outb) vsp
Xsram[2598] sram->in sram[2598]->out sram[2598]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2598]->out) 0
.nodeset V(sram[2598]->outb) vsp
Xsram[2599] sram->in sram[2599]->out sram[2599]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2599]->out) 0
.nodeset V(sram[2599]->outb) vsp
Xsram[2600] sram->in sram[2600]->out sram[2600]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2600]->out) 0
.nodeset V(sram[2600]->outb) vsp
Xsram[2601] sram->in sram[2601]->out sram[2601]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2601]->out) 0
.nodeset V(sram[2601]->outb) vsp
Xmux_2level_tapbuf_size16[65] chany[1][1]_midout[2] chany[1][1]_midout[3] chany[1][1]_midout[22] chany[1][1]_midout[23] chany[1][1]_midout[26] chany[1][1]_midout[27] chany[1][1]_midout[42] chany[1][1]_midout[43] chany[1][1]_midout[52] chany[1][1]_midout[53] chany[1][1]_midout[64] chany[1][1]_midout[65] chany[1][1]_midout[78] chany[1][1]_midout[79] chany[1][1]_midout[90] chany[1][1]_midout[91] grid[1][1]_pin[0][1][13] sram[2602]->outb sram[2602]->out sram[2603]->out sram[2603]->outb sram[2604]->out sram[2604]->outb sram[2605]->out sram[2605]->outb sram[2606]->outb sram[2606]->out sram[2607]->out sram[2607]->outb sram[2608]->out sram[2608]->outb sram[2609]->out sram[2609]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[65], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2602] sram->in sram[2602]->out sram[2602]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2602]->out) 0
.nodeset V(sram[2602]->outb) vsp
Xsram[2603] sram->in sram[2603]->out sram[2603]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2603]->out) 0
.nodeset V(sram[2603]->outb) vsp
Xsram[2604] sram->in sram[2604]->out sram[2604]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2604]->out) 0
.nodeset V(sram[2604]->outb) vsp
Xsram[2605] sram->in sram[2605]->out sram[2605]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2605]->out) 0
.nodeset V(sram[2605]->outb) vsp
Xsram[2606] sram->in sram[2606]->out sram[2606]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2606]->out) 0
.nodeset V(sram[2606]->outb) vsp
Xsram[2607] sram->in sram[2607]->out sram[2607]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2607]->out) 0
.nodeset V(sram[2607]->outb) vsp
Xsram[2608] sram->in sram[2608]->out sram[2608]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2608]->out) 0
.nodeset V(sram[2608]->outb) vsp
Xsram[2609] sram->in sram[2609]->out sram[2609]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2609]->out) 0
.nodeset V(sram[2609]->outb) vsp
Xmux_2level_tapbuf_size16[66] chany[1][1]_midout[2] chany[1][1]_midout[3] chany[1][1]_midout[22] chany[1][1]_midout[23] chany[1][1]_midout[28] chany[1][1]_midout[29] chany[1][1]_midout[40] chany[1][1]_midout[41] chany[1][1]_midout[52] chany[1][1]_midout[53] chany[1][1]_midout[64] chany[1][1]_midout[65] chany[1][1]_midout[80] chany[1][1]_midout[81] chany[1][1]_midout[92] chany[1][1]_midout[93] grid[1][1]_pin[0][1][17] sram[2610]->outb sram[2610]->out sram[2611]->out sram[2611]->outb sram[2612]->out sram[2612]->outb sram[2613]->out sram[2613]->outb sram[2614]->outb sram[2614]->out sram[2615]->out sram[2615]->outb sram[2616]->out sram[2616]->outb sram[2617]->out sram[2617]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[66], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2610] sram->in sram[2610]->out sram[2610]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2610]->out) 0
.nodeset V(sram[2610]->outb) vsp
Xsram[2611] sram->in sram[2611]->out sram[2611]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2611]->out) 0
.nodeset V(sram[2611]->outb) vsp
Xsram[2612] sram->in sram[2612]->out sram[2612]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2612]->out) 0
.nodeset V(sram[2612]->outb) vsp
Xsram[2613] sram->in sram[2613]->out sram[2613]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2613]->out) 0
.nodeset V(sram[2613]->outb) vsp
Xsram[2614] sram->in sram[2614]->out sram[2614]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2614]->out) 0
.nodeset V(sram[2614]->outb) vsp
Xsram[2615] sram->in sram[2615]->out sram[2615]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2615]->out) 0
.nodeset V(sram[2615]->outb) vsp
Xsram[2616] sram->in sram[2616]->out sram[2616]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2616]->out) 0
.nodeset V(sram[2616]->outb) vsp
Xsram[2617] sram->in sram[2617]->out sram[2617]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2617]->out) 0
.nodeset V(sram[2617]->outb) vsp
Xmux_2level_tapbuf_size16[67] chany[1][1]_midout[4] chany[1][1]_midout[5] chany[1][1]_midout[16] chany[1][1]_midout[17] chany[1][1]_midout[28] chany[1][1]_midout[29] chany[1][1]_midout[46] chany[1][1]_midout[47] chany[1][1]_midout[58] chany[1][1]_midout[59] chany[1][1]_midout[68] chany[1][1]_midout[69] chany[1][1]_midout[80] chany[1][1]_midout[81] chany[1][1]_midout[94] chany[1][1]_midout[95] grid[1][1]_pin[0][1][21] sram[2618]->outb sram[2618]->out sram[2619]->out sram[2619]->outb sram[2620]->out sram[2620]->outb sram[2621]->out sram[2621]->outb sram[2622]->outb sram[2622]->out sram[2623]->out sram[2623]->outb sram[2624]->out sram[2624]->outb sram[2625]->out sram[2625]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[67], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2618] sram->in sram[2618]->out sram[2618]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2618]->out) 0
.nodeset V(sram[2618]->outb) vsp
Xsram[2619] sram->in sram[2619]->out sram[2619]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2619]->out) 0
.nodeset V(sram[2619]->outb) vsp
Xsram[2620] sram->in sram[2620]->out sram[2620]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2620]->out) 0
.nodeset V(sram[2620]->outb) vsp
Xsram[2621] sram->in sram[2621]->out sram[2621]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2621]->out) 0
.nodeset V(sram[2621]->outb) vsp
Xsram[2622] sram->in sram[2622]->out sram[2622]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2622]->out) 0
.nodeset V(sram[2622]->outb) vsp
Xsram[2623] sram->in sram[2623]->out sram[2623]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2623]->out) 0
.nodeset V(sram[2623]->outb) vsp
Xsram[2624] sram->in sram[2624]->out sram[2624]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2624]->out) 0
.nodeset V(sram[2624]->outb) vsp
Xsram[2625] sram->in sram[2625]->out sram[2625]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2625]->out) 0
.nodeset V(sram[2625]->outb) vsp
Xmux_2level_tapbuf_size16[68] chany[1][1]_midout[4] chany[1][1]_midout[5] chany[1][1]_midout[18] chany[1][1]_midout[19] chany[1][1]_midout[38] chany[1][1]_midout[39] chany[1][1]_midout[46] chany[1][1]_midout[47] chany[1][1]_midout[58] chany[1][1]_midout[59] chany[1][1]_midout[70] chany[1][1]_midout[71] chany[1][1]_midout[82] chany[1][1]_midout[83] chany[1][1]_midout[94] chany[1][1]_midout[95] grid[1][1]_pin[0][1][25] sram[2626]->outb sram[2626]->out sram[2627]->out sram[2627]->outb sram[2628]->out sram[2628]->outb sram[2629]->out sram[2629]->outb sram[2630]->outb sram[2630]->out sram[2631]->out sram[2631]->outb sram[2632]->out sram[2632]->outb sram[2633]->out sram[2633]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[68], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2626] sram->in sram[2626]->out sram[2626]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2626]->out) 0
.nodeset V(sram[2626]->outb) vsp
Xsram[2627] sram->in sram[2627]->out sram[2627]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2627]->out) 0
.nodeset V(sram[2627]->outb) vsp
Xsram[2628] sram->in sram[2628]->out sram[2628]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2628]->out) 0
.nodeset V(sram[2628]->outb) vsp
Xsram[2629] sram->in sram[2629]->out sram[2629]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2629]->out) 0
.nodeset V(sram[2629]->outb) vsp
Xsram[2630] sram->in sram[2630]->out sram[2630]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2630]->out) 0
.nodeset V(sram[2630]->outb) vsp
Xsram[2631] sram->in sram[2631]->out sram[2631]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2631]->out) 0
.nodeset V(sram[2631]->outb) vsp
Xsram[2632] sram->in sram[2632]->out sram[2632]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2632]->out) 0
.nodeset V(sram[2632]->outb) vsp
Xsram[2633] sram->in sram[2633]->out sram[2633]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2633]->out) 0
.nodeset V(sram[2633]->outb) vsp
Xmux_2level_tapbuf_size16[69] chany[1][1]_midout[14] chany[1][1]_midout[15] chany[1][1]_midout[18] chany[1][1]_midout[19] chany[1][1]_midout[32] chany[1][1]_midout[33] chany[1][1]_midout[44] chany[1][1]_midout[45] chany[1][1]_midout[56] chany[1][1]_midout[57] chany[1][1]_midout[70] chany[1][1]_midout[71] chany[1][1]_midout[84] chany[1][1]_midout[85] chany[1][1]_midout[96] chany[1][1]_midout[97] grid[1][1]_pin[0][1][29] sram[2634]->outb sram[2634]->out sram[2635]->out sram[2635]->outb sram[2636]->out sram[2636]->outb sram[2637]->out sram[2637]->outb sram[2638]->outb sram[2638]->out sram[2639]->out sram[2639]->outb sram[2640]->out sram[2640]->outb sram[2641]->out sram[2641]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[69], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2634] sram->in sram[2634]->out sram[2634]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2634]->out) 0
.nodeset V(sram[2634]->outb) vsp
Xsram[2635] sram->in sram[2635]->out sram[2635]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2635]->out) 0
.nodeset V(sram[2635]->outb) vsp
Xsram[2636] sram->in sram[2636]->out sram[2636]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2636]->out) 0
.nodeset V(sram[2636]->outb) vsp
Xsram[2637] sram->in sram[2637]->out sram[2637]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2637]->out) 0
.nodeset V(sram[2637]->outb) vsp
Xsram[2638] sram->in sram[2638]->out sram[2638]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2638]->out) 0
.nodeset V(sram[2638]->outb) vsp
Xsram[2639] sram->in sram[2639]->out sram[2639]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2639]->out) 0
.nodeset V(sram[2639]->outb) vsp
Xsram[2640] sram->in sram[2640]->out sram[2640]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2640]->out) 0
.nodeset V(sram[2640]->outb) vsp
Xsram[2641] sram->in sram[2641]->out sram[2641]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2641]->out) 0
.nodeset V(sram[2641]->outb) vsp
Xmux_2level_tapbuf_size16[70] chany[1][1]_midout[8] chany[1][1]_midout[9] chany[1][1]_midout[20] chany[1][1]_midout[21] chany[1][1]_midout[32] chany[1][1]_midout[33] chany[1][1]_midout[44] chany[1][1]_midout[45] chany[1][1]_midout[62] chany[1][1]_midout[63] chany[1][1]_midout[72] chany[1][1]_midout[73] chany[1][1]_midout[84] chany[1][1]_midout[85] chany[1][1]_midout[96] chany[1][1]_midout[97] grid[1][1]_pin[0][1][33] sram[2642]->outb sram[2642]->out sram[2643]->out sram[2643]->outb sram[2644]->out sram[2644]->outb sram[2645]->out sram[2645]->outb sram[2646]->outb sram[2646]->out sram[2647]->out sram[2647]->outb sram[2648]->out sram[2648]->outb sram[2649]->out sram[2649]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[70], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2642] sram->in sram[2642]->out sram[2642]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2642]->out) 0
.nodeset V(sram[2642]->outb) vsp
Xsram[2643] sram->in sram[2643]->out sram[2643]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2643]->out) 0
.nodeset V(sram[2643]->outb) vsp
Xsram[2644] sram->in sram[2644]->out sram[2644]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2644]->out) 0
.nodeset V(sram[2644]->outb) vsp
Xsram[2645] sram->in sram[2645]->out sram[2645]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2645]->out) 0
.nodeset V(sram[2645]->outb) vsp
Xsram[2646] sram->in sram[2646]->out sram[2646]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2646]->out) 0
.nodeset V(sram[2646]->outb) vsp
Xsram[2647] sram->in sram[2647]->out sram[2647]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2647]->out) 0
.nodeset V(sram[2647]->outb) vsp
Xsram[2648] sram->in sram[2648]->out sram[2648]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2648]->out) 0
.nodeset V(sram[2648]->outb) vsp
Xsram[2649] sram->in sram[2649]->out sram[2649]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2649]->out) 0
.nodeset V(sram[2649]->outb) vsp
Xmux_2level_tapbuf_size16[71] chany[1][1]_midout[8] chany[1][1]_midout[9] chany[1][1]_midout[30] chany[1][1]_midout[31] chany[1][1]_midout[34] chany[1][1]_midout[35] chany[1][1]_midout[50] chany[1][1]_midout[51] chany[1][1]_midout[62] chany[1][1]_midout[63] chany[1][1]_midout[74] chany[1][1]_midout[75] chany[1][1]_midout[86] chany[1][1]_midout[87] chany[1][1]_midout[98] chany[1][1]_midout[99] grid[1][1]_pin[0][1][37] sram[2650]->outb sram[2650]->out sram[2651]->out sram[2651]->outb sram[2652]->out sram[2652]->outb sram[2653]->out sram[2653]->outb sram[2654]->outb sram[2654]->out sram[2655]->out sram[2655]->outb sram[2656]->out sram[2656]->outb sram[2657]->out sram[2657]->outb svdd sgnd mux_2level_tapbuf_size16
***** SRAM bits for MUX[71], level=2, select_path_id=0. *****
*****10001000*****
Xsram[2650] sram->in sram[2650]->out sram[2650]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2650]->out) 0
.nodeset V(sram[2650]->outb) vsp
Xsram[2651] sram->in sram[2651]->out sram[2651]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2651]->out) 0
.nodeset V(sram[2651]->outb) vsp
Xsram[2652] sram->in sram[2652]->out sram[2652]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2652]->out) 0
.nodeset V(sram[2652]->outb) vsp
Xsram[2653] sram->in sram[2653]->out sram[2653]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2653]->out) 0
.nodeset V(sram[2653]->outb) vsp
Xsram[2654] sram->in sram[2654]->out sram[2654]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2654]->out) 0
.nodeset V(sram[2654]->outb) vsp
Xsram[2655] sram->in sram[2655]->out sram[2655]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2655]->out) 0
.nodeset V(sram[2655]->outb) vsp
Xsram[2656] sram->in sram[2656]->out sram[2656]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2656]->out) 0
.nodeset V(sram[2656]->outb) vsp
Xsram[2657] sram->in sram[2657]->out sram[2657]->outb gvdd_sram_cbs sgnd  sram6T
.nodeset V(sram[2657]->out) 0
.nodeset V(sram[2657]->outb) vsp
.eom
