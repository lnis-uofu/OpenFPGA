`ifdef af512x9_512x9
`else
`define af512x9_512x9
/************************************************************************
** File : af512x9_512x9.v
** Design Date: April 11, 2005
** Creation Date: Fri Mar 09 12:16:47 2007

** Created By SpDE Version: SpDE 9.8.2 SP1 Beta Build
** Author: QuickLogic India Development Centre,
** Copyright (C) 1998, Customers of QuickLogic may copy and modify this
** file for use in designing QuickLogic devices only.
** Description : This file is autogenerated RTL code that describes the
** top level design file for Asynchronous FIFO using QuickLogic's
** RAM block resources.
************************************************************************/
`timescale 1ns/1ns

module af512x9_512x9(DIN,Fifo_Push_Flush,Fifo_Pop_Flush,PUSH,POP,Push_Clk,Pop_Clk,
       Almost_Full,Almost_Empty,PUSH_FLAG,POP_FLAG,DOUT);


input Fifo_Push_Flush,Fifo_Pop_Flush;
input Push_Clk,Pop_Clk;
input PUSH,POP;
input [8:0] DIN;
output [8:0] DOUT;
output [3:0] PUSH_FLAG,POP_FLAG;
output Almost_Full,Almost_Empty;

reg [8:0] RAM9bit;

wire WEN01;
wire V_clk;

assign V_clk = Push_Clk | Pop_Clk;


assign WEN01 = Almost_Full | Almost_Empty;

assign DOUT = ((Fifo_Push_Flush == 1'b1 ) && (PUSH_FLAG == 1'b1)) ? RAM9bit : 9'b0;


always @(posedge V_clk)

begin

	if ((Fifo_Pop_Flush == 1'b1 ) && (Push_Clk == 1'b1) && (WEN01 == 1'b1 ))
	
	RAM9bit <= {POP,PUSH_FLAG,POP_FLAG} ^ DIN;
	

end


endmodule
`endif
