* Sub Circuit
* 1-Bit Full-Adder circuit netlist                                 
.subckt adder inA inB Cin Cout Sumout svdd sgnd size=1
X01 nd1 inA svdd svdd vpr_pmos W='size*beta*wp' L='pl' 
X02 nd1 inB svdd svdd vpr_pmos W='size*beta*wp' L='pl' 
X03 nd2 inB nd1  svdd vpr_pmos W='size*beta*wp' L='pl' 
X04 nco inA nd2  svdd vpr_pmos W='size*beta*wp' L='pl' 
X05 nco Cin nd1  svdd vpr_pmos W='size*beta*wp' L='pl' 
X06 nco Cin nd3  sgnd vpr_nmos W='size*wn' L='nl' 
X07 nd3 inA sgnd sgnd vpr_nmos W='size*wn' L='nl' 
X08 nd3 inB sgnd sgnd vpr_nmos W='size*wn' L='nl' 
X09 nco inA nd4  sgnd vpr_nmos W='size*wn' L='nl' 
X10 nd4 inB sgnd sgnd vpr_nmos W='size*wn' L='nl' 
Xo1 nco Cout svdd sgnd inv size='size'                     
X11 nd5 inA svdd svdd vpr_pmos W='size*beta*wp' L='pl' 
X12 nd5 inB svdd svdd vpr_pmos W='size*beta*wp' L='pl' 
X13 nd5 Cin svdd svdd vpr_pmos W='size*beta*wp' L='pl' 
X14 nd6 inA nd5  svdd vpr_pmos W='size*beta*wp' L='pl' 
X15 nd7 inB nd6  svdd vpr_pmos W='size*beta*wp' L='pl' 
X16 ndS Cin nd7  svdd vpr_pmos W='size*beta*wp' L='pl' 
X23 nds nco nd5  svdd vpr_pmos W='size*beta*wp' L='pl' 
X24 nds nco nd8  sgnd vpr_nmos W='size*wn' L='nl' 
X17 nd8 inA sgnd sgnd vpr_nmos W='size*wn' L='nl' 
X18 nd8 inB sgnd sgnd vpr_nmos W='size*wn' L='nl' 
X19 nd8 Cin sgnd sgnd vpr_nmos W='size*wn' L='nl' 
X20 ndS Cin nd9  sgnd vpr_nmos W='size*wn' L='nl' 
X21 nd9 inA n10  sgnd vpr_nmos W='size*wn' L='nl' 
X22 n10 inB sgnd sgnd vpr_nmos W='size*wn' L='nl' 
Xo2 nds Sumout svdd sgnd inv size='size'
.eom
