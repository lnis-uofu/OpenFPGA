// Benchmark "TOP" written by ABC on Mon Feb  4 17:33:45 2019

module seq ( 
    i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_,
    i_11_, i_12_, i_13_, i_14_, i_15_, i_16_, i_17_, i_18_, i_19_, i_20_,
    i_21_, i_22_, i_23_, i_24_, i_25_, i_26_, i_27_, i_28_, i_29_, i_30_,
    i_31_, i_32_, i_33_, i_34_, i_35_, i_36_, i_37_, i_38_, i_39_, i_40_,
    o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_,
    o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_,
    o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_,
    o_31_, o_32_, o_33_, o_34_  );
  input  i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_,
    i_10_, i_11_, i_12_, i_13_, i_14_, i_15_, i_16_, i_17_, i_18_, i_19_,
    i_20_, i_21_, i_22_, i_23_, i_24_, i_25_, i_26_, i_27_, i_28_, i_29_,
    i_30_, i_31_, i_32_, i_33_, i_34_, i_35_, i_36_, i_37_, i_38_, i_39_,
    i_40_;
  output o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_,
    o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_,
    o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_,
    o_31_, o_32_, o_33_, o_34_;
  wire n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
    n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
    n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
    n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
    n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
    n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
    n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
    n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
    n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
    n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
    n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
    n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
    n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
    n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
    n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
    n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
    n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
    n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
    n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
    n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
    n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
    n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
    n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
    n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
    n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
    n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
    n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
    n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
    n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
    n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
    n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
    n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
    n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
    n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
    n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
    n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
    n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
    n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
    n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
    n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
    n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
    n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
    n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
    n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
    n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
    n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
    n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
    n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
    n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
    n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
    n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
    n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
    n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
    n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
    n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
    n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
    n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
    n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
    n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
    n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
    n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
    n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
    n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
    n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
    n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
    n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
    n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
    n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
    n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
    n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
    n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
    n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
    n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
    n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095;
  assign o_0_ = ~n852;
  assign o_1_ = ~n754;
  assign o_2_ = ~n606;
  assign o_3_ = ~n488;
  assign o_4_ = ~n426;
  assign o_5_ = ~n986 | ~n990 | ~n980 | ~n982 | n191 | n192 | n189 | n190;
  assign o_6_ = ~n306;
  assign o_7_ = ~n188;
  assign o_8_ = ~n111;
  assign o_9_ = ~n185;
  assign o_10_ = ~n823 | ~n833 | n181 | ~n175 | n180;
  assign o_11_ = ~n179;
  assign o_12_ = ~n708 & ~n407 & i_8_ & n112;
  assign o_13_ = ~n174;
  assign o_14_ = ~n173;
  assign o_15_ = ~n149;
  assign o_16_ = ~n172;
  assign o_17_ = ~n1076 | ~n1078 | ~n437 | ~n812 | n165 | n166 | n163 | n164;
  assign o_18_ = ~n800;
  assign o_19_ = ~n162;
  assign o_20_ = ~n728;
  assign o_21_ = ~n161;
  assign o_22_ = n156 | n157 | n154 | n155 | n160 | ~n662 | n158 | n159;
  assign o_23_ = ~n153;
  assign o_24_ = ~n146;
  assign o_25_ = ~n138;
  assign o_26_ = ~n134;
  assign o_27_ = ~n131;
  assign o_28_ = ~n128;
  assign o_29_ = ~n617;
  assign o_30_ = ~n1029 | n122 | n123;
  assign o_31_ = ~n128 | n116 | n117 | n115 | n113 | n114;
  assign o_32_ = ~n1034;
  assign o_33_ = ~n576;
  assign o_34_ = ~n535;
  assign n111 = n223 & n149 & (n224 | n225);
  assign n112 = ~n1094 & (~i_37_ | (~n288 & ~n523));
  assign n113 = n200 & (~n715 | (~i_39_ & ~n277));
  assign n114 = ~n610 & n471 & n578;
  assign n115 = n579 & ~n222 & ~n257;
  assign n116 = n194 & n200;
  assign n117 = n385 & (~n387 | ~n715);
  assign n118 = ~n909 & ~n410 & ~n877;
  assign n119 = ~n906 & ~n410 & ~n877;
  assign n120 = ~n909 & ~n414 & ~n877;
  assign n121 = ~n906 & ~n414 & ~n877;
  assign n122 = ~n946 & (n582 | ~n701 | ~n864);
  assign n123 = n118 | n119 | n120 | n121;
  assign n124 = n355 | n911;
  assign n125 = n577 | n284 | n536;
  assign n126 = n515 | n284 | n577;
  assign n127 = n899 | n760 | n816;
  assign n128 = n127 & n126 & n124 & n125;
  assign n129 = ~n117 & n141 & (~n194 | n627);
  assign n130 = n954 & n953 & ~n622 & ~n619 & n618 & n328 & n312 & n319;
  assign n131 = n129 & n130;
  assign n132 = n630 | n476 | n360;
  assign n133 = ~n199 & n135 & ~n195;
  assign n134 = ~n203 & n132 & n133;
  assign n135 = n872 | n893 | ~i_34_ | n611;
  assign n136 = n607 & (n608 | n609);
  assign n137 = n130 & ~n201;
  assign n138 = n137 & n129 & n136 & n128 & n135;
  assign n139 = ~n594 & ~i_37_ & i_39_;
  assign n140 = ~n902 & (n139 | (~n307 & ~n594));
  assign n141 = n952 & ~n626 & ~n625 & n616 & n315 & ~n140 & ~n113 & ~n123;
  assign n142 = n631 & ~n203 & ~n117 & n124;
  assign n143 = n577 | n325 | i_39_;
  assign n144 = ~n194 | n627;
  assign n145 = n1034 & n126 & n127;
  assign n146 = n145 & n144 & n143 & n142 & n137 & n133 & n136 & n141;
  assign n147 = n407 | n644 | n284 | n462;
  assign n148 = i_35_ | i_34_ | n640 | n307;
  assign n149 = ~i_7_ | ~i_33_;
  assign n150 = n646 | ~i_37_ | n400;
  assign n151 = n646 | n515 | n645;
  assign n152 = n648 | n519 | n647;
  assign n153 = ~n1047 & ~n651 & n152 & n151 & n150 & n149 & n147 & n148;
  assign n154 = ~n666 & (~n231 | ~n355 | ~n647);
  assign n155 = ~i_40_ & (n667 | (~n338 & n663));
  assign n156 = ~n611 & n663;
  assign n157 = n673 & n671 & n672;
  assign n158 = ~n685 & (~n669 | (n674 & ~n920));
  assign n159 = n671 & ~i_7_ & i_32_;
  assign n160 = ~n708 & n670 & i_37_ & ~n333;
  assign n161 = n684 & i_33_ & (i_7_ | n680);
  assign n162 = n765 & n766 & (n767 | n267);
  assign n163 = n813 & ~n1093 & (~i_29_ | n814);
  assign n164 = ~n859 & n649 & n650;
  assign n165 = ~n926 & (~n514 | ~n675);
  assign n166 = ~n428 & (~n1075 | (n471 & ~n610));
  assign n167 = n338 | n820;
  assign n168 = n821 | n514;
  assign n169 = n630 | n476 | n815 | n816;
  assign n170 = n333 | n307 | n709 | n788;
  assign n171 = n451 | n817 | i_40_;
  assign n172 = ~n819 & n171 & n170 & n169 & n167 & n168;
  assign n173 = n492 & (~i_13_ | n407 | n822);
  assign n174 = n492 & (n536 | n333 | n537);
  assign n175 = n817 | n549;
  assign n176 = n918 | n405 | n917;
  assign n177 = n826 | n447 | n825;
  assign n178 = n823 & (n225 | n817);
  assign n179 = ~n828 & n178 & n177 & n175 & n176;
  assign n180 = i_15_ & n834 & i_20_ & i_21_;
  assign n181 = n578 & (n830 | (n561 & ~n585));
  assign n182 = n857 | n583 | n456 | n350;
  assign n183 = n222 | n221 | n220;
  assign n184 = n149 & ~n215 & (n210 | n216);
  assign n185 = n184 & n182 & n183;
  assign n186 = n240 & n239 & n238 & n182;
  assign n187 = n223 & (n869 | (n701 & n242));
  assign n188 = ~n245 & n187 & n184 & n186;
  assign n189 = n293 & (n378 | (~i_23_ & ~n377));
  assign n190 = ~n910 & (~n890 | (~i_37_ & ~n307));
  assign n191 = n385 & (n194 | ~n908);
  assign n192 = (n194 | n347) & (n384 | ~n951);
  assign n193 = i_1_ | i_4_ | i_2_ | i_3_;
  assign n194 = i_39_ & n653;
  assign n195 = n193 & ~n896 & (n194 | ~n280);
  assign n196 = ~n332 & (n628 | (i_0_ & i_4_));
  assign n197 = ~n333 & n629;
  assign n198 = ~n225 & ~n933;
  assign n199 = (n196 | n197) & (n198 | ~n955);
  assign n200 = ~n414 & ~i_24_ & ~n375;
  assign n201 = ~n593 & (~n609 | (~n489 & ~n900));
  assign n202 = i_2_ & ~n359;
  assign n203 = n202 & ~n333 & (n198 | ~n955);
  assign n204 = i_11_ | ~n861;
  assign n205 = ~i_17_ | n314;
  assign n206 = i_12_ | n413;
  assign n207 = (n204 | n205) & (n206 | ~n229);
  assign n208 = n211 & (~n729 | (n961 & n962));
  assign n209 = ~i_16_ | n314;
  assign n210 = n207 & n208 & (n204 | n209);
  assign n211 = i_12_ | ~i_15_ | ~i_17_ | ~n229;
  assign n212 = n962 & n961;
  assign n213 = n211 & (n212 | ~n729);
  assign n214 = n207 & (n204 | n209);
  assign n215 = ~n565 & ~n862 & (~n213 | ~n214);
  assign n216 = n565 | n318;
  assign n217 = ~i_18_ | n428;
  assign n218 = n217 & (~i_15_ | ~n963);
  assign n219 = n404 | ~n963;
  assign n220 = n219 & (~i_19_ | i_21_ | n218);
  assign n221 = ~i_23_ | n241;
  assign n222 = n864 | n333;
  assign n223 = n283 | n677 | n740 | ~n853;
  assign n224 = n841 | n500;
  assign n225 = ~i_38_ | n771;
  assign n226 = i_12_ & n861;
  assign n227 = i_22_ & (~n217 | (i_15_ & n226));
  assign n228 = i_15_ & i_22_;
  assign n229 = i_11_ & n861;
  assign n230 = i_19_ & (n227 | (n228 & n229));
  assign n231 = ~i_40_ | n440;
  assign n232 = ~i_38_ | i_39_;
  assign n233 = n231 & n232;
  assign n234 = n428 | n580 | n265 | n613;
  assign n235 = i_35_ | ~i_33_ | ~i_34_;
  assign n236 = n779 | i_32_ | n428;
  assign n237 = n234 & (~i_21_ | n235 | n236);
  assign n238 = n856 | n583 | n225 | n519;
  assign n239 = (~i_22_ | n237) & (n866 | ~n964);
  assign n240 = n965 & (n864 | n869);
  assign n241 = ~i_22_ | ~i_24_;
  assign n242 = n870 | n596;
  assign n243 = n242 | n241 | n218;
  assign n244 = ~n225 | ~n690;
  assign n245 = ~n333 & (~n243 | (n244 & ~n537));
  assign n246 = ~n872 & (~n966 | (~n225 & ~n875));
  assign n247 = n657 | n866 | ~n194 | ~n578;
  assign n248 = n767 | i_37_ | n350;
  assign n249 = n375 | n588 | ~i_24_ | ~n293;
  assign n250 = ~n246 & (n536 | n775 | n875);
  assign n251 = n250 & n249 & n247 & n248;
  assign n252 = ~i_18_ | n253;
  assign n253 = n314 & n310;
  assign n254 = n252 & (~i_19_ | n253);
  assign n255 = ~i_15_ | ~i_18_ | ~i_19_ | ~n293;
  assign n256 = ~i_9_ | n323;
  assign n257 = n255 & (n254 | n256);
  assign n258 = (~i_29_ & n825) | (n366 & (i_29_ | n825));
  assign n259 = i_29_ | n323;
  assign n260 = n258 & (~i_30_ | n259);
  assign n261 = ~n382 & (~n468 | (~n277 & ~n283));
  assign n262 = n644 | n256 | ~n624;
  assign n263 = n907 & n895;
  assign n264 = ~n261 & n262 & (n260 | n263);
  assign n265 = n859 | n400;
  assign n266 = (n476 | n875) & (n400 | n474);
  assign n267 = ~i_40_ | n876;
  assign n268 = ~i_34_ | n858;
  assign n269 = n265 & n266 & (n267 | n268);
  assign n270 = i_10_ & i_27_;
  assign n271 = n890 | n881 | n322;
  assign n272 = (n456 | n887) & (n817 | n338);
  assign n273 = n739 | n890 | n721;
  assign n274 = n271 & n272 & (~i_11_ | n273);
  assign n275 = n283 | n320;
  assign n276 = i_36_ | n307;
  assign n277 = i_36_ | n647;
  assign n278 = n275 & n276 & (~i_39_ | n277);
  assign n279 = n396 | ~n653;
  assign n280 = i_39_ | n456;
  assign n281 = n278 & n279 & n280;
  assign n282 = n536 | n500;
  assign n283 = ~i_39_ | ~i_40_;
  assign n284 = i_37_ | n858;
  assign n285 = n282 & (n283 | n284);
  assign n286 = (~i_40_ | n325) & (n284 | n440);
  assign n287 = n286 & n285;
  assign n288 = ~i_38_ | i_40_;
  assign n289 = ~n244 & (~i_37_ | n288);
  assign n290 = i_12_ | i_11_;
  assign n291 = n290 & n228 & ~n256;
  assign n292 = i_18_ & n228;
  assign n293 = ~n410 | ~n414;
  assign n294 = ~n613 & (n291 | (n292 & n293));
  assign n295 = ~i_37_ & ~n558 & (n294 | ~n775);
  assign n296 = ~n400 & (n295 | (~n474 & ~n775));
  assign n297 = ~n887 & (n194 | ~n611);
  assign n298 = n256 | n504 | ~n624 | n878;
  assign n299 = i_32_ | i_13_ | n877 | n382;
  assign n300 = n880 | n771 | n875;
  assign n301 = n967 & (n263 | n857 | n365);
  assign n302 = ~n296 & n970 & (n289 | n337);
  assign n303 = (n281 | n889) & (~i_40_ | n274);
  assign n304 = n971 & (n269 | n888);
  assign n305 = n251 & n973 & (n897 | n702);
  assign n306 = n305 & n304 & n303 & n302 & n301 & n300 & n298 & n299;
  assign n307 = i_38_ | ~i_40_;
  assign n308 = n310 | n901;
  assign n309 = n307 | n594;
  assign n310 = ~i_11_ | ~i_15_;
  assign n311 = n903 | n462 | n881;
  assign n312 = (n310 | n311) & (n308 | n309);
  assign n313 = ~n835 & ~n881 & (~n451 | ~n690);
  assign n314 = ~i_12_ | ~i_15_;
  assign n315 = ~n116 & ~n313 & (n311 | n314);
  assign n316 = n903 | n253 | n216;
  assign n317 = n902 & n308;
  assign n318 = n594 | n863;
  assign n319 = n316 & (n317 | n318);
  assign n320 = i_36_ | i_37_;
  assign n321 = n276 & n280 & (~i_39_ | n320);
  assign n322 = i_15_ | n323;
  assign n323 = i_7_ | i_5_;
  assign n324 = n322 & (i_12_ | n323);
  assign n325 = i_38_ | n858;
  assign n326 = (~i_40_ | n325) & (~i_39_ | n284);
  assign n327 = ~n376 & ~n881 & (~n324 | ~n411);
  assign n328 = ~n139 | n308;
  assign n329 = n974 & (n321 | n889);
  assign n330 = (~n194 | n975) & (n318 | ~n1095);
  assign n331 = n330 & n329 & n328 & n319 & n315 & n312 & ~n140 & ~n195;
  assign n332 = i_7_ | n333;
  assign n333 = i_34_ | n407;
  assign n334 = (n333 | ~n914) & (n332 | ~n976);
  assign n335 = (n334 | n916) & (n273 | ~n290);
  assign n336 = n978 & (n821 | (n451 & n549));
  assign n337 = n767 | n463;
  assign n338 = ~i_37_ | n232;
  assign n339 = n335 & n336 & (n337 | n338);
  assign n340 = n835 | ~i_15_ | ~n290;
  assign n341 = n340 & (~i_15_ | i_18_ | ~n293);
  assign n342 = n314 | n913;
  assign n343 = n310 | n913;
  assign n344 = i_21_ | n407;
  assign n345 = i_19_ | n341;
  assign n346 = n342 & n343 & (n344 | n345);
  assign n347 = ~i_40_ & ~n908;
  assign n348 = n790 | i_34_ | n898;
  assign n349 = (n523 | n890) & (n400 | n912);
  assign n350 = ~i_39_ | i_40_;
  assign n351 = n463 | n645;
  assign n352 = n348 & n349 & (n350 | n351);
  assign n353 = n322 | n565 | n231;
  assign n354 = i_38_ | n577;
  assign n355 = ~i_38_ | n396;
  assign n356 = n353 & n354 & (n317 | n355);
  assign n357 = ~i_25_ & i_26_;
  assign n358 = i_4_ & i_1_;
  assign n359 = ~i_0_ | i_7_;
  assign n360 = ~n914 & (n358 | n359);
  assign n361 = n975 | n908;
  assign n362 = n915 | n360 | n333;
  assign n363 = n519 | n878 | n879 | n549;
  assign n364 = n175 & n363 & n361 & n362;
  assign n365 = ~i_29_ | n323;
  assign n366 = ~i_28_ | n323;
  assign n367 = n365 & n366 & (~i_30_ | n323);
  assign n368 = n284 | n596;
  assign n369 = n368 & n318;
  assign n370 = i_14_ | n369 | n314 | n410;
  assign n371 = i_34_ | n477;
  assign n372 = n370 & (n367 | n350 | n371);
  assign n373 = ~i_15_ | i_21_;
  assign n374 = n333 | n536 | n439;
  assign n375 = n657 | n874;
  assign n376 = i_40_ | n859;
  assign n377 = (n375 | n376) & (n373 | n374);
  assign n378 = ~n235 & ~n779 & (~n906 | ~n909);
  assign n379 = n721 | ~i_0_ | n657;
  assign n380 = n350 | n379 | i_36_ | ~i_37_;
  assign n381 = n279 | n693;
  assign n382 = i_12_ | n411;
  assign n383 = n381 | n382 | ~i_13_ | i_31_;
  assign n384 = ~n909 & ~n410 & ~n657;
  assign n385 = ~n410 & ~i_24_ & ~n375;
  assign n386 = n260 & (i_30_ | n365);
  assign n387 = ~n194 & (i_39_ | n277);
  assign n388 = n956 | n919;
  assign n389 = n451 | i_40_ | n821;
  assign n390 = ~i_13_ | n886;
  assign n391 = n388 & n389 & (n387 | n390);
  assign n392 = i_13_ | n277 | n283 | ~n853;
  assign n393 = n407 | n514 | ~i_40_ | n400;
  assign n394 = n235 | n456 | i_32_ | ~i_39_;
  assign n395 = n392 & n393 & (~i_13_ | n394);
  assign n396 = i_39_ | i_40_;
  assign n397 = n267 & (~i_37_ | n396);
  assign n398 = n871 | i_34_ | n225;
  assign n399 = (n523 | n376) & (n351 | n690);
  assign n400 = i_36_ | n868;
  assign n401 = n398 & n399 & (n397 | n400);
  assign n402 = n322 & (~i_24_ | n323);
  assign n403 = n373 | n256 | ~n290;
  assign n404 = ~i_18_ | n373;
  assign n405 = n403 & (~n293 | n404);
  assign n406 = ~i_17_ | n407;
  assign n407 = i_32_ | ~i_33_;
  assign n408 = n406 & (~i_16_ | n407);
  assign n409 = (i_11_ | n314) & (i_12_ | n310);
  assign n410 = ~i_11_ | n323;
  assign n411 = i_11_ | n323;
  assign n412 = (n209 | n411) & (n206 | n410);
  assign n413 = ~i_15_ | ~i_16_;
  assign n414 = ~i_12_ | n323;
  assign n415 = n412 & (i_14_ | n413 | n414);
  assign n416 = (n406 | n415) & (n256 | ~n992);
  assign n417 = ~n323 & ~n333 & (~n958 | ~n991);
  assign n418 = ~i_39_ & (~n892 | ~n979);
  assign n419 = ~n1089 & (i_40_ | (n175 & n957));
  assign n420 = n1004 & (n910 | n790);
  assign n421 = (n267 | n821) & (n401 | n872);
  assign n422 = n1003 & (n695 | n416);
  assign n423 = ~n418 & (n474 | (n919 & n1002));
  assign n424 = n1000 & (~i_31_ | (~n417 & n1001));
  assign n425 = n998 & n135 & n176 & n997 & n995 & n996;
  assign n426 = n425 & n424 & n423 & n422 & n421 & n420 & n419 & n391;
  assign n427 = n929 | n428 | n400;
  assign n428 = n854 & (i_5_ | n310);
  assign n429 = n427 & (n428 | n400 | n344);
  assign n430 = ~i_3_ | n432;
  assign n431 = ~i_2_ | n432;
  assign n432 = ~i_0_ | i_32_;
  assign n433 = n430 & n431 & (n358 | n432);
  assign n434 = ~n270 | n396 | n756 | ~n853;
  assign n435 = n863 | ~n649 | ~n650;
  assign n436 = (n859 | n926) & (n925 | ~n1014);
  assign n437 = n436 & n435 & n434 & n149;
  assign n438 = n858 | i_5_ | ~i_31_;
  assign n439 = ~i_37_ | ~i_35_ | i_36_;
  assign n440 = i_38_ | ~i_39_;
  assign n441 = (n439 | n440) & (~n314 | n438);
  assign n442 = ~i_39_ & n307;
  assign n443 = ~i_35_ | n898;
  assign n444 = ~i_36_ | n923;
  assign n445 = (n283 | n444) & (n396 | n443);
  assign n446 = ~n350 & (~n915 | (~n452 & ~n803));
  assign n447 = i_29_ | i_30_;
  assign n448 = ~i_5_ & ~n907 & (i_28_ | n447);
  assign n449 = n542 | n806 | ~i_15_ | i_17_;
  assign n450 = ~n448 & (~i_36_ | n231 | n740);
  assign n451 = ~i_37_ | n462;
  assign n452 = i_9_ | i_5_;
  assign n453 = n449 & n450 & (n451 | n452);
  assign n454 = (~i_4_ | n432) & (i_32_ | ~n628);
  assign n455 = n454 & n430 & n431;
  assign n456 = i_36_ | n477;
  assign n457 = n456 & (i_36_ | ~i_39_);
  assign n458 = i_11_ & ~n452;
  assign n459 = ~n928 & (~n1010 | (n458 & ~n867));
  assign n460 = n932 | i_36_ | ~n863;
  assign n461 = ~n459 & n460 & (~i_40_ | ~n1009);
  assign n462 = ~i_38_ | ~i_39_;
  assign n463 = ~i_0_ | n884;
  assign n464 = n288 & n462 & (n463 | n396);
  assign n465 = ~i_9_ | ~i_14_ | ~n644 | n737;
  assign n466 = ~i_14_ | ~n644;
  assign n467 = n465 & (n466 | ~n729);
  assign n468 = n456 | n771;
  assign n469 = (i_13_ | n468) & (~i_15_ | ~n624);
  assign n470 = n150 & (i_5_ | n407 | n371);
  assign n471 = ~i_23_ & ~n407;
  assign n472 = ~n690 & ~n875 & (~n344 | n471);
  assign n473 = n929 & n344;
  assign n474 = ~i_37_ | n307;
  assign n475 = ~n472 & (n268 | n473 | n474);
  assign n476 = i_40_ | n536;
  assign n477 = ~i_37_ | i_38_;
  assign n478 = n476 & n477;
  assign n479 = n928 | n519 | n763;
  assign n480 = n479 & (i_18_ | n373 | ~n829);
  assign n481 = ~n693 & (~n1008 | (~n467 & ~n702));
  assign n482 = ~n333 & (~n441 | ~n1012 | ~n1013);
  assign n483 = (n536 | n926) & (n453 | ~n853);
  assign n484 = (n675 | n224) & (n464 | n761);
  assign n485 = (n461 | n504) & (n859 | n427);
  assign n486 = n1019 & n1020 & (n428 | n475);
  assign n487 = n1017 & n1018 & (n927 | ~n1006);
  assign n488 = n487 & n486 & n485 & n484 & n483 & ~n482 & n437 & ~n481;
  assign n489 = i_31_ | n333;
  assign n490 = (n368 | n489) & (n216 | ~n466);
  assign n491 = n333 | n870;
  assign n492 = n149 & (n491 | (n231 & n355));
  assign n493 = ~n904 & (i_9_ | ~n672);
  assign n494 = ~i_31_ & ~n290 & (~n279 | ~n287);
  assign n495 = n858 | ~i_5_ | n493;
  assign n496 = (n788 | n690) & (n476 | n933);
  assign n497 = n496 & ~n494 & n495;
  assign n498 = ~i_34_ & ~n320 & (~n462 | ~n536);
  assign n499 = (n400 | n675) & (n594 | ~n863);
  assign n500 = ~i_37_ | n858;
  assign n501 = ~n498 & n499 & (n231 | n500);
  assign n502 = n763 | n718;
  assign n503 = n504 | n280;
  assign n504 = i_35_ | n855;
  assign n505 = n502 & n503 & (n278 | n504);
  assign n506 = ~n284 & ~i_15_ & i_39_;
  assign n507 = ~n690 & ~i_35_ & ~i_37_;
  assign n508 = ~n489 & (n506 | (n507 & ~n644));
  assign n509 = n815 | n739 | n935;
  assign n510 = i_2_ | ~i_0_ | i_1_;
  assign n511 = n657 | n444;
  assign n512 = ~n283 | n235 | n277;
  assign n513 = n509 & (n510 | (n511 & n512));
  assign n514 = i_37_ | n536;
  assign n515 = i_38_ | i_40_;
  assign n516 = n514 & (i_37_ | n515);
  assign n517 = n511 & (~i_40_ | n338 | n739);
  assign n518 = (n504 | n859) & (n690 | n718);
  assign n519 = ~i_33_ | n858;
  assign n520 = n517 & n518 & (n516 | n519);
  assign n521 = n451 | ~i_40_ | n268;
  assign n522 = n860 & n882;
  assign n523 = ~i_36_ | n868;
  assign n524 = n521 & (n522 | n523);
  assign n525 = ~n510 & ~i_3_ & ~i_4_;
  assign n526 = n525 & (~n706 | (i_39_ & ~n756));
  assign n527 = ~n526 & (~i_5_ | i_36_ | ~n674);
  assign n528 = i_9_ & (n508 | (~n490 & ~n904));
  assign n529 = (n490 | n672) & (n497 | n333);
  assign n530 = (n505 | n878) & (n224 | n355);
  assign n531 = n501 | n936;
  assign n532 = (n513 | n925) & (n520 | n648);
  assign n533 = (n527 | ~n853) & (n524 | n934);
  assign n534 = n749 & (~i_11_ | n550 | n741);
  assign n535 = n534 & n533 & n532 & n531 & n530 & n529 & n492 & ~n528;
  assign n536 = i_38_ | i_39_;
  assign n537 = ~i_35_ | n871;
  assign n538 = ~i_17_ | n539;
  assign n539 = i_32_ | i_31_;
  assign n540 = n538 & (~i_16_ | n539);
  assign n541 = ~n540 & (~n503 | (~n504 & ~n542));
  assign n542 = i_36_ | n462;
  assign n543 = n503 & (~i_40_ | n504 | n542);
  assign n544 = n543 | i_14_ | n540;
  assign n545 = (i_12_ | n1022) & (i_15_ | n940);
  assign n546 = n462 | n500;
  assign n547 = n544 & n545 & (n489 | n546);
  assign n548 = n756 | n771 | n333;
  assign n549 = i_37_ | n232;
  assign n550 = n407 | n894;
  assign n551 = n548 & (n270 | n549 | n550);
  assign n552 = n1023 & (n218 | n241 | n941);
  assign n553 = n1024 & (n350 | n756);
  assign n554 = i_31_ | i_15_ | i_5_;
  assign n555 = n552 & n553 & (n287 | n554);
  assign n556 = n511 & (n235 | n277);
  assign n557 = ~n815 & ~n657 & i_36_ & ~n476;
  assign n558 = ~i_38_ | ~i_40_;
  assign n559 = (n474 | n523) & (n558 | ~n959);
  assign n560 = ~i_13_ & ~n407;
  assign n561 = ~n231 & ~n268;
  assign n562 = n560 & (n561 | (~n476 & ~n875));
  assign n563 = ~n863 | ~n890;
  assign n564 = ~n881 & (~n307 | n563 | ~n770);
  assign n565 = i_31_ | n407;
  assign n566 = n284 | n355;
  assign n567 = ~n562 & ~n564 & (n565 | n566);
  assign n568 = ~n869 & (~n941 | ~n942);
  assign n569 = ~n925 & (n557 | (~n510 & ~n556));
  assign n570 = (n204 | n1022) & (~i_32_ | i_33_);
  assign n571 = (n333 | n555) & (n801 | ~n943);
  assign n572 = (n381 | n554) & (n547 | ~n861);
  assign n573 = ~n568 & (n931 | (n222 & n937));
  assign n574 = n1025 & (~n290 | n550 | n741);
  assign n575 = ~n569 & n1026 & (n935 | n939);
  assign n576 = n575 & n574 & n573 & n572 & n571 & n570 & n551 & n186;
  assign n577 = n899 | n841 | n816;
  assign n578 = n293 & n873;
  assign n579 = ~i_23_ & n921;
  assign n580 = ~i_21_ | ~i_23_;
  assign n581 = ~n870 & n580 & ~n690;
  assign n582 = ~n462 & ~n870;
  assign n583 = i_28_ | i_5_ | i_29_;
  assign n584 = n583 & (i_5_ | ~n960);
  assign n585 = ~i_25_ | n407;
  assign n586 = n585 & (~i_26_ | n407);
  assign n587 = n841 | n566;
  assign n588 = i_37_ | n771;
  assign n589 = n400 | n613;
  assign n590 = n587 & (n428 | n588 | n589);
  assign n591 = ~i_22_ | n373;
  assign n592 = (n217 | ~n921) & (n591 | ~n963);
  assign n593 = n500 | n790;
  assign n594 = i_34_ | n858;
  assign n595 = n593 & (n594 | n225);
  assign n596 = ~i_38_ | n283;
  assign n597 = n596 & n476;
  assign n598 = n1030 & (n771 | n870 | n931);
  assign n599 = (n537 | n690) & (n1031 | n933);
  assign n600 = n598 & n599 & (n597 | n439);
  assign n601 = (n801 | n939) & (n588 | ~n943);
  assign n602 = (n586 | n822) & (n600 | n333);
  assign n603 = n224 | n790;
  assign n604 = n1032 & (n592 | n596 | n589);
  assign n605 = n374 | n220 | n221;
  assign n606 = n605 & n604 & n603 & n602 & n184 & n601 & n590 & n551;
  assign n607 = n900 | n608 | n489;
  assign n608 = n771 | n803;
  assign n609 = n447 | n366 | n489;
  assign n610 = n400 | n376;
  assign n611 = i_40_ | n514;
  assign n612 = n610 & (n400 | n611);
  assign n613 = ~i_24_ | n407;
  assign n614 = (n612 | n613) & (n224 | n231);
  assign n615 = n614 | ~n293 | n591;
  assign n616 = n767 | n895;
  assign n617 = n616 & n615 & n136 & ~n201;
  assign n618 = i_23_ | n222 | ~n293 | n373;
  assign n619 = ~n265 & (~n342 | ~n343);
  assign n620 = ~n410 & n905;
  assign n621 = ~n414 & n905;
  assign n622 = ~n318 & (n620 | n621);
  assign n623 = ~n375 & ~i_23_ & n293;
  assign n624 = ~n350 & n653;
  assign n625 = n624 & (n384 | n623 | ~n951);
  assign n626 = ~n950 & (n194 | ~n949);
  assign n627 = n906 | n657 | n410;
  assign n628 = i_0_ & i_1_;
  assign n629 = i_3_ & ~n359;
  assign n630 = n333 | n443;
  assign n631 = n515 | n630 | n360;
  assign n632 = (i_37_ | n690) & (n463 | n923);
  assign n633 = n632 & n588 & n514;
  assign n634 = n290 & (i_9_ | i_16_);
  assign n635 = i_9_ | i_16_ | i_36_ | ~i_39_;
  assign n636 = n867 | n290;
  assign n637 = n635 & n636 & (n307 | n634);
  assign n638 = n1090 & (~i_37_ | n648 | n855);
  assign n639 = n1035 & n1036 & (n894 | n646);
  assign n640 = i_15_ | n407;
  assign n641 = n638 & n639 & (n284 | n640);
  assign n642 = i_3_ | n899;
  assign n643 = n642 | i_38_;
  assign n644 = i_11_ & i_12_;
  assign n645 = ~i_37_ | n868;
  assign n646 = ~i_0_ | n407;
  assign n647 = i_38_ | i_37_;
  assign n648 = i_32_ | i_0_ | ~i_5_;
  assign n649 = ~n268 & ~n407;
  assign n650 = n884 | i_2_ | i_3_;
  assign n651 = n649 & (~n643 | (~n477 & n650));
  assign n652 = ~n841 & (~n1037 | (n283 & ~n803));
  assign n653 = i_38_ & ~n320;
  assign n654 = ~n693 & (~n1038 | (i_40_ & n653));
  assign n655 = ~n594 & (~n922 | ~n936 | ~n1040);
  assign n656 = ~n333 & (~n1043 | ~n1044 | ~n1045);
  assign n657 = ~i_35_ | n855;
  assign n658 = (n267 | n519) & (~n194 | n657);
  assign n659 = ~n708 & (~n1049 | (~n333 & ~n955));
  assign n660 = ~i_5_ | n721;
  assign n661 = (n514 | n718) & (n657 | n715);
  assign n662 = ~n659 & (n660 | (n658 & n661));
  assign n663 = ~i_7_ & n792;
  assign n664 = n663 & (~n1048 | (i_9_ & ~n314));
  assign n665 = ~i_11_ | i_7_ | ~i_9_;
  assign n666 = ~n664 & (~i_15_ | n665 | ~n792);
  assign n667 = ~n920 & ~n665 & ~n314 & ~i_31_ & ~i_37_;
  assign n668 = n923 & ~n904 & n440 & n232 & n288;
  assign n669 = n668 | ~i_33_ | n594;
  assign n670 = (i_35_ & ~n690) | (~n225 & (~i_35_ | ~n690));
  assign n671 = i_33_ & ~n594;
  assign n672 = ~i_16_ | ~i_17_;
  assign n673 = ~i_9_ & ~n685;
  assign n674 = ~i_15_ | n466;
  assign n675 = i_38_ | n771;
  assign n676 = (n675 | n443) & (n596 | n537);
  assign n677 = ~i_36_ | n647;
  assign n678 = n268 & (i_35_ | n677 | n396);
  assign n679 = n500 | n596 | i_6_ | ~i_34_;
  assign n680 = n679 & ~n1091 & (~i_32_ | n678);
  assign n681 = n1050 & (n523 | n923);
  assign n682 = (n645 | n690) & (n860 | n894);
  assign n683 = n681 & n682 & (n516 | n268);
  assign n684 = n323 | i_0_ | n683;
  assign n685 = ~i_5_ | i_7_;
  assign n686 = i_17_ | n407;
  assign n687 = (n685 | n686) & (n407 | ~n673);
  assign n688 = (~n673 | n686) & (i_16_ | n687);
  assign n689 = ~n408 & (~n318 | (~n594 & ~n859));
  assign n690 = ~i_38_ | n350;
  assign n691 = ~n689 & (n284 | n333 | n690);
  assign n692 = n456 | n283;
  assign n693 = i_35_ | n407;
  assign n694 = ~n829 & (n692 | n693);
  assign n695 = n318 & n862;
  assign n696 = n408 | n695 | i_14_;
  assign n697 = i_9_ & (~n696 | (~i_12_ & ~n691));
  assign n698 = ~i_16_ | n406 | ~n466 | n695;
  assign n699 = n594 | n922;
  assign n700 = ~n697 & n698 & (n493 | n699);
  assign n701 = n870 | n476;
  assign n702 = n283 | ~n653;
  assign n703 = (n440 | n284) & (n771 | n325);
  assign n704 = n468 & (~i_13_ | i_36_ | n675);
  assign n705 = n704 & n703 & n702 & n701 & n566 & n282;
  assign n706 = n771 | n444;
  assign n707 = n706 & (i_40_ | n542);
  assign n708 = i_0_ | n685;
  assign n709 = i_7_ | n290;
  assign n710 = (n705 | n709) & (n707 | n708);
  assign n711 = n785 & n867 & n780;
  assign n712 = n711 & (i_36_ | n288);
  assign n713 = ~i_31_ | n721;
  assign n714 = (n711 | n660) & (n712 | n713);
  assign n715 = ~i_40_ | n908;
  assign n716 = n279 & n715 & (~i_39_ | n277);
  assign n717 = n1053 & n503 & (n716 | n504);
  assign n718 = i_36_ | n855;
  assign n719 = n658 & n717 & (n522 | n718);
  assign n720 = (~i_13_ | n715) & (~i_9_ | ~n194);
  assign n721 = i_7_ | i_32_;
  assign n722 = (n719 | n721) & (n720 | n332);
  assign n723 = i_11_ | n691 | i_7_ | ~i_9_;
  assign n724 = (i_7_ | n700) & (n710 | n333);
  assign n725 = n694 | n709;
  assign n726 = (n714 | n504) & (i_15_ | n722);
  assign n727 = n1054 & n1055 & (n688 | n594);
  assign n728 = n727 & n726 & n725 & n724 & n662 & n723;
  assign n729 = i_15_ & ~n672;
  assign n730 = n729 & ~i_5_ & i_12_;
  assign n731 = ~i_14_ & (n730 | (n226 & ~n737));
  assign n732 = ~n282 & (~n213 | ~n214 | n731);
  assign n733 = n1058 & (n931 | (n1057 & n285));
  assign n734 = ~n732 & (n439 | (n283 & n355));
  assign n735 = n1030 & (n537 | (n350 & n440));
  assign n736 = n735 & n734 & n733 & n441;
  assign n737 = ~i_15_ | n904;
  assign n738 = (n428 | n672) & (n737 | ~n963);
  assign n739 = ~i_36_ | n855;
  assign n740 = i_11_ | ~i_12_;
  assign n741 = ~i_40_ | n890;
  assign n742 = n741 | n739 | n740;
  assign n743 = ~n563 & (i_37_ | ~i_40_ | ~n232);
  assign n744 = n560 & n938;
  assign n745 = n744 & (~n1056 | (~n594 & ~n743));
  assign n746 = ~n931 & (~n381 | ~n694 | ~n883);
  assign n747 = ~n504 & ~n702;
  assign n748 = ~i_32_ & (~n742 | (~n738 & n747));
  assign n749 = n368 | n467 | n333;
  assign n750 = n1059 & (n586 | n647 | n523);
  assign n751 = n1060 & (~n863 | n920 | n932);
  assign n752 = (n860 | n939) & (n736 | n333);
  assign n753 = ~n746 & (~n943 | (n474 & n956));
  assign n754 = n753 & n752 & n751 & n750 & n749 & ~n748 & n149 & n590;
  assign n755 = ~i_36_ | n477;
  assign n756 = ~i_38_ | n871;
  assign n757 = (~i_40_ | n755) & (n283 | n756);
  assign n758 = n924 | n283 | n235;
  assign n759 = n758 & (n757 | n657);
  assign n760 = ~i_38_ | n630;
  assign n761 = n841 | n284;
  assign n762 = n760 & (n761 | (n536 & n515));
  assign n763 = i_40_ | n549;
  assign n764 = n741 & n763;
  assign n765 = (n821 | n935) & (n764 | n944);
  assign n766 = n1062 & (n456 | n396 | n897);
  assign n767 = n872 | n523;
  assign n768 = ~i_15_ | i_40_ | ~n644 | n803;
  assign n769 = n546 & n768;
  assign n770 = i_37_ | n283;
  assign n771 = i_39_ | ~i_40_;
  assign n772 = n288 & n770 & (~i_37_ | n771);
  assign n773 = (i_11_ | n307) & (n270 | n288);
  assign n774 = ~n872 & (~n338 | ~n912);
  assign n775 = ~n873 | ~n293 | n613;
  assign n776 = ~n774 & (n775 | (n477 & n558));
  assign n777 = ~i_37_ | ~i_39_;
  assign n778 = n675 & n690 & n777 & n588;
  assign n779 = ~i_40_ | n867;
  assign n780 = i_36_ | n232;
  assign n781 = n779 & n277 & (i_40_ | n780);
  assign n782 = n729 & ~i_7_ & ~n466;
  assign n783 = (n253 | n256) & (~n293 | n413);
  assign n784 = n333 | n816 | n915 | n815;
  assign n785 = n924 & n277;
  assign n786 = i_31_ | n504;
  assign n787 = n784 & (n785 | n323 | n786);
  assign n788 = i_37_ | n893;
  assign n789 = (n476 | n788) & (~i_38_ | n351);
  assign n790 = i_38_ | n350;
  assign n791 = n790 & (i_39_ | i_37_);
  assign n792 = ~i_31_ & n671;
  assign n793 = ~n386 & n792 & (~n225 | ~n895);
  assign n794 = ~n817 & (~n232 | (i_37_ & ~n350));
  assign n795 = n1092 & (~i_36_ | n773 | n891);
  assign n796 = n1071 & (n588 | n887);
  assign n797 = (n820 | n923) & (n855 | ~n1064);
  assign n798 = n1069 & n1070 & (n787 | n396);
  assign n799 = n1068 & n1067 & n1066 & n957 & n823 & ~n794 & ~n159 & ~n793;
  assign n800 = n799 & n798 & n797 & n796 & n795 & n251;
  assign n801 = n882 & n859;
  assign n802 = n801 & n611;
  assign n803 = ~i_38_ | n858;
  assign n804 = n282 & (~i_39_ | n803);
  assign n805 = n326 & n804 & (n284 | n288);
  assign n806 = ~i_12_ | n452;
  assign n807 = ~n458 & n806;
  assign n808 = n546 & (n350 | n803);
  assign n809 = n804 | n807 | ~i_15_ | i_17_;
  assign n810 = n805 | n807 | ~i_15_ | i_16_;
  assign n811 = n809 & n810 & (n808 | n452);
  assign n812 = n433 | i_40_ | n755 | n657;
  assign n813 = ~i_5_ & (~n907 | (~n350 & ~n456));
  assign n814 = n853 & ~i_31_ & ~i_28_ & i_30_;
  assign n815 = i_2_ | ~n628;
  assign n816 = i_7_ | i_3_ | ~i_4_;
  assign n817 = n872 | n268;
  assign n818 = ~n332 & n525;
  assign n819 = n818 & (~n955 | (~n232 & ~n933));
  assign n820 = (i_40_ & n944) | (n821 & (~i_40_ | n944));
  assign n821 = n872 | n894;
  assign n822 = n523 | n514;
  assign n823 = n817 | n741;
  assign n824 = ~n540 & ~n256 & ~n409;
  assign n825 = i_28_ | n323;
  assign n826 = n907 | i_31_ | n693;
  assign n827 = ~n503 | n747;
  assign n828 = n827 & (n824 | (~n412 & ~n538));
  assign n829 = ~n333 & n582;
  assign n830 = i_24_ & i_23_ & i_25_ & n829;
  assign n831 = n1053 & ~n865 & n917;
  assign n832 = ~i_24_ | i_32_;
  assign n833 = n831 | ~i_25_ | ~n293 | n832 | ~n873;
  assign n834 = n293 & (~n1080 | (~n221 & n829));
  assign n835 = i_9_ | n323;
  assign n836 = n252 | n832 | n835 | ~n865;
  assign n837 = n863 | n400;
  assign n838 = n256 | ~i_40_ | n254 | n613 | n837;
  assign n839 = n928 | n786 | n410 | i_12_ | i_17_;
  assign n840 = n839 & (~i_21_ | ~n293 | n375);
  assign n841 = ~i_34_ | n407;
  assign n842 = n325 | n283 | n841;
  assign n843 = ~i_18_ & ~n340 & (~n222 | n829);
  assign n844 = n293 & ~n927 & (n561 | ~n612);
  assign n845 = ~n826 & (~n900 | (~n366 & ~n447));
  assign n846 = n579 & (~n836 | ~n838);
  assign n847 = n331 & n1088 & (n350 | n957);
  assign n848 = n1087 & n1086 & (n675 | n919);
  assign n849 = ~n845 & n1084 & (n842 | n879);
  assign n850 = n1083 & n1082 & (n222 | n345);
  assign n851 = n1081 & n1054 & n953 & ~n843 & n616 & ~n201 & ~n113 & ~n199;
  assign n852 = n851 & n850 & n849 & n848 & n847 & n178 & n142 & n391;
  assign n853 = ~i_32_ & ~n504;
  assign n854 = i_5_ | n314;
  assign n855 = ~i_33_ | i_34_;
  assign n856 = i_30_ | n539;
  assign n857 = n856 | n504;
  assign n858 = i_36_ | i_35_;
  assign n859 = i_37_ | n462;
  assign n860 = ~i_40_ | n859;
  assign n861 = ~i_5_ & i_9_;
  assign n862 = n860 | n594;
  assign n863 = ~i_37_ | n536;
  assign n864 = n439 | n675;
  assign n865 = ~n468 & ~n657;
  assign n866 = ~i_23_ | n832;
  assign n867 = i_36_ | n440;
  assign n868 = i_34_ | ~i_35_;
  assign n869 = n333 | n428 | ~i_21_ | n241;
  assign n870 = ~i_35_ | n320;
  assign n871 = ~i_36_ | i_37_;
  assign n872 = i_7_ | n407;
  assign n873 = n228 & i_21_;
  assign n874 = ~i_15_ | i_32_;
  assign n875 = i_37_ | n868;
  assign n876 = ~i_37_ | n440;
  assign n877 = n235 | n692;
  assign n878 = i_15_ | n539;
  assign n879 = ~i_13_ | n323;
  assign n880 = n879 | n640;
  assign n881 = n594 | n565;
  assign n882 = ~i_40_ | n863;
  assign n883 = n333 | n307 | n439;
  assign n884 = i_4_ | i_1_;
  assign n885 = n489 | ~i_13_ | n382;
  assign n886 = n382 | i_32_ | n657;
  assign n887 = i_13_ | n886;
  assign n888 = n640 | i_13_ | n323;
  assign n889 = n879 | n504 | n878;
  assign n890 = i_37_ | n440;
  assign n891 = i_7_ | ~n853;
  assign n892 = n756 | n270 | n891;
  assign n893 = i_35_ | ~i_36_;
  assign n894 = i_34_ | n893;
  assign n895 = i_40_ | n876;
  assign n896 = n235 | n721;
  assign n897 = n650 | n896;
  assign n898 = ~i_36_ | ~i_37_;
  assign n899 = ~i_2_ | ~i_0_ | i_1_;
  assign n900 = n825 | ~i_29_ | ~i_30_;
  assign n901 = n835 | i_16_ | n565;
  assign n902 = n314 | n901;
  assign n903 = i_17_ | n835;
  assign n904 = ~i_16_ & ~i_17_;
  assign n905 = n904 & i_15_ & ~n565;
  assign n906 = i_22_ | n874;
  assign n907 = ~i_40_ | n780;
  assign n908 = i_36_ | n536;
  assign n909 = i_32_ | n373;
  assign n910 = n463 | n817;
  assign n911 = n788 | ~n270 | n332;
  assign n912 = ~i_37_ | n515;
  assign n913 = n344 | i_18_ | n835;
  assign n914 = n629 | n202;
  assign n915 = ~i_35_ | n477;
  assign n916 = ~i_38_ | n893;
  assign n917 = n657 | n702;
  assign n918 = i_32_ | n241;
  assign n919 = n400 | n880;
  assign n920 = i_36_ | n504;
  assign n921 = ~i_21_ & i_22_;
  assign n922 = ~i_31_ | n407;
  assign n923 = ~i_37_ | ~i_38_;
  assign n924 = i_36_ | n923;
  assign n925 = i_32_ | i_3_ | ~i_4_;
  assign n926 = i_24_ | n428 | n407 | n400;
  assign n927 = ~i_15_ | n407;
  assign n928 = i_16_ | n874;
  assign n929 = i_22_ | n407;
  assign n930 = i_40_ | n235 | n899 | n925;
  assign n931 = i_13_ | i_15_ | i_5_;
  assign n932 = i_32_ | i_5_ | ~i_31_;
  assign n933 = ~i_37_ | n893;
  assign n934 = ~i_6_ | n407;
  assign n935 = i_40_ | n863;
  assign n936 = ~i_5_ | n407;
  assign n937 = ~n829 & n842;
  assign n938 = ~i_5_ & ~n290;
  assign n939 = ~n649 | n650;
  assign n940 = n565 | i_34_ | ~n507;
  assign n941 = n283 | n870;
  assign n942 = n647 | ~i_35_ | n396;
  assign n943 = ~n400 & n744;
  assign n944 = n400 | n872;
  assign n945 = n333 | ~i_15_ | ~i_24_;
  assign n946 = n945 | i_22_ | ~n293;
  assign n947 = n277 | n396;
  assign n948 = n400 | n882;
  assign n949 = n947 & n468;
  assign n950 = n906 | n657 | n414;
  assign n951 = n909 | n657 | n414;
  assign n952 = (n949 | n627) & (n947 | n951);
  assign n953 = i_37_ | n317 | n594 | n288;
  assign n954 = n1033 & (n346 | n948);
  assign n955 = n596 | n788;
  assign n956 = n514 & n859;
  assign n957 = n379 | n924;
  assign n958 = (i_38_ & n500) | (n284 & (~i_38_ | n500));
  assign n959 = (~i_37_ & ~n523) | (~n268 & (i_37_ | ~n523));
  assign n960 = (i_28_ & (i_29_ | i_30_)) | (i_29_ & ~i_30_);
  assign n961 = i_5_ | n740;
  assign n962 = i_12_ | i_5_ | ~i_11_;
  assign n963 = n226 | n229;
  assign n964 = n865 & (n230 | (n292 & n963));
  assign n965 = (n841 | n608) & (n233 | n761);
  assign n966 = (n400 | n876) & (n647 | n523);
  assign n967 = ~n578 | n224 | n231;
  assign n968 = n882 | n881 | n322;
  assign n969 = n968 & (i_31_ | n264 | ~n853);
  assign n970 = n969 & (n257 | n221 | n883);
  assign n971 = ~n297 & (n885 | (n287 & n566));
  assign n972 = (n821 | n895) & (n396 | n892);
  assign n973 = n972 & (n588 | n390);
  assign n974 = ~n327 & (n885 | (n282 & n326));
  assign n975 = n950 & n627;
  assign n976 = n884 & i_0_;
  assign n977 = n539 | n519 | n382 | n890;
  assign n978 = n977 & (n400 | n514 | n888);
  assign n979 = n357 | n677 | n657 | n721;
  assign n980 = n248 & n607 & n127 & n383 & n979 & n380;
  assign n981 = n907 | n857 | n259;
  assign n982 = n981 & (n771 | n277 | n887);
  assign n983 = (n232 | n911) & (n372 | n565);
  assign n984 = n983 & (n817 | n770);
  assign n985 = (n352 | n872) & (n356 | n284);
  assign n986 = n984 & n985 & (n368 | ~n1095);
  assign n987 = (n346 | n837) & (n975 | n280);
  assign n988 = (~i_40_ & n364) | (n339 & (i_40_ | n364));
  assign n989 = n331 & n988 & (~n200 | n908);
  assign n990 = n987 & n989 & (n882 | n821);
  assign n991 = (~n283 | n803) & (~i_39_ | n325);
  assign n992 = ~n408 & (~n409 | (~i_14_ & ~n314));
  assign n993 = n890 | n594 | n888;
  assign n994 = n993 & (n456 | n390);
  assign n995 = n447 | n825 | ~n853 | n907;
  assign n996 = i_5_ | n713 | ~n904 | n920;
  assign n997 = n268 | n876 | n880;
  assign n998 = n893 | n332 | n283 | i_38_ | n740;
  assign n999 = n491 | n402 | n675;
  assign n1000 = n999 & (n386 | n407 | n593);
  assign n1001 = i_36_ | ~n672 | n835 | ~n853;
  assign n1002 = ~i_23_ | n257 | n589 | ~n921;
  assign n1003 = (n395 | n382) & (n324 | n699);
  assign n1004 = (n225 | n337) & (n817 | n895);
  assign n1005 = ~i_32_ & (~n503 | (~n519 & ~n860));
  assign n1006 = ~n212 & (~n318 | (~n284 & ~n462));
  assign n1007 = n469 | i_12_ | i_5_;
  assign n1008 = n1007 & (n931 | (n468 & ~n624));
  assign n1009 = ~n455 & (~n898 | (i_36_ & ~n462));
  assign n1010 = (n807 | n276) & (n457 | n806);
  assign n1011 = (n442 | n933) & (n445 | n463);
  assign n1012 = ~n446 & n1011 & (i_14_ | n438);
  assign n1013 = (n439 | n515) & (~n244 | n537);
  assign n1014 = ~n899 & (~n511 | (~n235 & ~n908));
  assign n1015 = i_17_ | n874 | n503 | n806;
  assign n1016 = n1015 & (n854 | ~n904 | ~n1005);
  assign n1017 = n1016 & (i_25_ | n407 | n822);
  assign n1018 = n912 | n433 | n657;
  assign n1019 = (n429 | n478) & (n807 | n480);
  assign n1020 = (n320 | n930) & (n470 | n350);
  assign n1021 = n827 & ~i_5_ & n466;
  assign n1022 = ~n541 & n940;
  assign n1023 = n931 | n942;
  assign n1024 = (n476 | n933) & (n231 | n443);
  assign n1025 = n174 & (~i_16_ | n538 | ~n1021);
  assign n1026 = (n559 | n934) & (n567 | ~n938);
  assign n1027 = n293 & (n581 | (~i_21_ & ~n701));
  assign n1028 = ~i_24_ | i_21_ | i_23_ | n222 | n257;
  assign n1029 = n124 & n1028 & (n945 | ~n1027);
  assign n1030 = n225 | ~i_35_ | i_37_;
  assign n1031 = n307 & n440;
  assign n1032 = n565 | n584 | n595;
  assign n1033 = (~n384 | n947) & (n862 | ~n1095);
  assign n1034 = n944 | i_40_ | n338;
  assign n1035 = n936 | i_34_ | i_35_;
  assign n1036 = n642 | n407 | n645;
  assign n1037 = (n284 | n463) & (n1031 | n500);
  assign n1038 = n907 & (n677 | n396);
  assign n1039 = n462 | i_9_ | n407;
  assign n1040 = n1039 & (n440 | n640);
  assign n1041 = (~i_35_ | n633) & (n307 | n893);
  assign n1042 = (n232 | n788) & (n350 | n915);
  assign n1043 = n1041 & n1042 & (i_40_ | n916);
  assign n1044 = (i_38_ | n537) & (n439 | ~n690);
  assign n1045 = (~n283 | n456) & (~i_39_ | n933);
  assign n1046 = (~i_38_ | n641) & (n637 | ~n853);
  assign n1047 = n655 | n652 | n654 | ~n1046 | n656 | ~n937;
  assign n1048 = n209 & (~i_16_ | n310);
  assign n1049 = n760 & (n277 | ~n283 | n693);
  assign n1050 = n898 | i_34_ | n225;
  assign n1051 = n443 | i_0_ | n476;
  assign n1052 = n1051 & (i_6_ | n676);
  assign n1053 = n657 | n947;
  assign n1054 = n677 | n891 | ~i_11_ | n283;
  assign n1055 = n660 | n376 | n718;
  assign n1056 = n566 & (n500 | n231);
  assign n1057 = (n536 | n870) & (n1031 | n284);
  assign n1058 = n596 | n933;
  assign n1059 = n699 | i_5_ | n493;
  assign n1060 = ~n745 & (n476 | n788 | n841);
  assign n1061 = n759 | ~i_6_ | n721;
  assign n1062 = n1061 & (n762 | n816 | n510);
  assign n1063 = i_14_ & (~n209 | (i_17_ & ~n314));
  assign n1064 = ~n1074 & (n782 | (~n665 & n1063));
  assign n1065 = i_31_ | n769 | n855 | n256;
  assign n1066 = n1065 & (n781 | n783 | n786);
  assign n1067 = (n789 | n872) & (n791 | n910);
  assign n1068 = n916 | ~i_40_ | ~n818;
  assign n1069 = n888 | n771 | n875;
  assign n1070 = ~n578 | n842;
  assign n1071 = (n776 | n400) & (n778 | n821);
  assign n1072 = ~n455 & (~n706 | (~n283 & ~n756));
  assign n1073 = n268 | n473 | n267;
  assign n1074 = n282 & n368;
  assign n1075 = n1073 & (n489 | ~n904 | n1074);
  assign n1076 = (n489 | n811) & (n504 | ~n1072);
  assign n1077 = (n277 | n930) & (n429 | n802);
  assign n1078 = n1077 & (n630 | n790);
  assign n1079 = ~n649 | ~i_22_ | n231;
  assign n1080 = n1079 & (n831 | n918);
  assign n1081 = n537 | n332 | n536 | i_25_ | i_26_;
  assign n1082 = ~n844 & (n556 | n642 | n721);
  assign n1083 = n885 | n284 | n288;
  assign n1084 = n889 | i_40_ | ~n653;
  assign n1085 = (n390 | n715) & (n337 | n923);
  assign n1086 = ~n846 & n1085 & (~n194 | n840);
  assign n1087 = (n775 | n948) & (n864 | n946);
  assign n1088 = (~n621 | n862) & (n647 | n910);
  assign n1089 = i_40_ & (~n994 | (~n514 & ~n910));
  assign n1090 = n519 | i_37_ | i_32_ | n634;
  assign n1091 = ~i_34_ & (~n1052 | (i_32_ & n858));
  assign n1092 = i_36_ | n772 | n897;
  assign n1093 = ~i_29_ & (~i_28_ | n857);
  assign n1094 = ~i_37_ & (n268 | n515);
  assign n1095 = n620 | n621;
endmodule


