// Benchmark "top" written by ABC on Mon Feb  4 17:32:32 2019

module frisc (  
    tin_pdata_8_8_, tin_pdata_0_0_, tin_pdata_7_7_, preset_0_0_,
    tin_pdata_2_2_, tin_pdata_9_9_, tin_pdata_1_1_, tin_pdata_4_4_, pclk,
    pirq_0_0_, tin_pdata_10_10_, tin_pdata_3_3_, tin_pdata_6_6_,
    tin_pdata_15_15_, tin_pdata_11_11_, tin_pdata_14_14_, tin_pdata_12_12_,
    tin_pdata_5_5_, preset, tin_pdata_13_13_,
    ppeakb_7_7_, ppeakp_12_12_, ppeakp_0_0_, ppeaka_7_7_, ppeaki_15_15_,
    ppeaki_11_11_, ppeaki_3_3_, paddress_3_3_, pdata_8_8_, pdata_0_0_,
    ppeakb_14_14_, ppeakb_10_10_, ppeakb_8_8_, ppeakp_1_1_, ppeaka_14_14_,
    ppeaka_10_10_, ppeaka_8_8_, ppeaki_4_4_, paddress_15_15_,
    paddress_11_11_, paddress_2_2_, ppeakb_9_9_, ppeakp_2_2_, ppeaka_9_9_,
    ppeaks_12_12_, ppeaks_0_0_, ppeaki_5_5_, paddress_5_5_, pdata_7_7_,
    ppeakb_15_15_, ppeakp_3_3_, pwr_0_0_, ppeaks_1_1_, ppeaki_6_6_,
    paddress_4_4_, piack_0_0_, ppeakp_13_13_, ppeakp_4_4_, ppeaka_15_15_,
    ppeaka_11_11_, ppeaks_2_2_, ppeaki_7_7_, paddress_10_10_,
    paddress_7_7_, pdata_2_2_, ppeakp_5_5_, ppeaks_13_13_, ppeaks_3_3_,
    ppeaki_14_14_, ppeaki_10_10_, ppeaki_8_8_, paddress_6_6_, ppeakp_6_6_,
    ppeaks_4_4_, ppeaki_9_9_, paddress_9_9_, pdata_9_9_, pdata_1_1_,
    ppeakb_11_11_, ppeakp_7_7_, ppeaks_5_5_, paddress_13_13_,
    paddress_8_8_, ppeakp_14_14_, ppeakp_10_10_, ppeakp_8_8_, ppeaks_6_6_,
    ppeaki_13_13_, pdata_4_4_, ppeakb_0_0_, ppeakp_9_9_, ppeaka_0_0_,
    ppeaks_7_7_, ppeakb_1_1_, ppeaka_1_1_, ppeaks_10_10_, ppeaks_8_8_,
    pdata_10_10_, pdata_3_3_, ppeakb_12_12_, ppeakb_2_2_, ppeaka_12_12_,
    ppeaka_2_2_, ppeaks_15_15_, ppeaks_9_9_, ppeakb_3_3_, ppeakp_15_15_,
    ppeakp_11_11_, ppeaka_13_13_, ppeaka_3_3_, paddress_14_14_,
    paddress_12_12_, pdata_6_6_, ppeakb_13_13_, ppeakb_4_4_, pdn,
    ppeaka_4_4_, ppeaki_0_0_, prd_0_0_, pdata_15_15_, pdata_11_11_,
    ppeakb_5_5_, ppeaka_5_5_, ppeaks_14_14_, ppeaki_1_1_, paddress_1_1_,
    pdata_14_14_, pdata_12_12_, pdata_5_5_, ppeakb_6_6_, ppeaka_6_6_,
    ppeaks_11_11_, ppeaki_12_12_, ppeaki_2_2_, paddress_0_0_, pdata_13_13_  );
  input  tin_pdata_8_8_, tin_pdata_0_0_, tin_pdata_7_7_, preset_0_0_,
    tin_pdata_2_2_, tin_pdata_9_9_, tin_pdata_1_1_, tin_pdata_4_4_, pclk,
    pirq_0_0_, tin_pdata_10_10_, tin_pdata_3_3_, tin_pdata_6_6_,
    tin_pdata_15_15_, tin_pdata_11_11_, tin_pdata_14_14_, tin_pdata_12_12_,
    tin_pdata_5_5_, preset, tin_pdata_13_13_;
  output ppeakb_7_7_, ppeakp_12_12_, ppeakp_0_0_, ppeaka_7_7_, ppeaki_15_15_,
    ppeaki_11_11_, ppeaki_3_3_, paddress_3_3_, pdata_8_8_, pdata_0_0_,
    ppeakb_14_14_, ppeakb_10_10_, ppeakb_8_8_, ppeakp_1_1_, ppeaka_14_14_,
    ppeaka_10_10_, ppeaka_8_8_, ppeaki_4_4_, paddress_15_15_,
    paddress_11_11_, paddress_2_2_, ppeakb_9_9_, ppeakp_2_2_, ppeaka_9_9_,
    ppeaks_12_12_, ppeaks_0_0_, ppeaki_5_5_, paddress_5_5_, pdata_7_7_,
    ppeakb_15_15_, ppeakp_3_3_, pwr_0_0_, ppeaks_1_1_, ppeaki_6_6_,
    paddress_4_4_, piack_0_0_, ppeakp_13_13_, ppeakp_4_4_, ppeaka_15_15_,
    ppeaka_11_11_, ppeaks_2_2_, ppeaki_7_7_, paddress_10_10_,
    paddress_7_7_, pdata_2_2_, ppeakp_5_5_, ppeaks_13_13_, ppeaks_3_3_,
    ppeaki_14_14_, ppeaki_10_10_, ppeaki_8_8_, paddress_6_6_, ppeakp_6_6_,
    ppeaks_4_4_, ppeaki_9_9_, paddress_9_9_, pdata_9_9_, pdata_1_1_,
    ppeakb_11_11_, ppeakp_7_7_, ppeaks_5_5_, paddress_13_13_,
    paddress_8_8_, ppeakp_14_14_, ppeakp_10_10_, ppeakp_8_8_, ppeaks_6_6_,
    ppeaki_13_13_, pdata_4_4_, ppeakb_0_0_, ppeakp_9_9_, ppeaka_0_0_,
    ppeaks_7_7_, ppeakb_1_1_, ppeaka_1_1_, ppeaks_10_10_, ppeaks_8_8_,
    pdata_10_10_, pdata_3_3_, ppeakb_12_12_, ppeakb_2_2_, ppeaka_12_12_,
    ppeaka_2_2_, ppeaks_15_15_, ppeaks_9_9_, ppeakb_3_3_, ppeakp_15_15_,
    ppeakp_11_11_, ppeaka_13_13_, ppeaka_3_3_, paddress_14_14_,
    paddress_12_12_, pdata_6_6_, ppeakb_13_13_, ppeakb_4_4_, pdn,
    ppeaka_4_4_, ppeaki_0_0_, prd_0_0_, pdata_15_15_, pdata_11_11_,
    ppeakb_5_5_, ppeaka_5_5_, ppeaks_14_14_, ppeaki_1_1_, paddress_1_1_,
    pdata_14_14_, pdata_12_12_, pdata_5_5_, ppeakb_6_6_, ppeaka_6_6_,
    ppeaks_11_11_, ppeaki_12_12_, ppeaki_2_2_, paddress_0_0_, pdata_13_13_;
  reg ndout, ppeakb_12_12_, ppeakb_1_1_, ppeaka_6_6_, \[4295] , \[4310] ,
    ppeaks_5_5_, ppeakp_10_10_, \[4355] , \[4370] , \[4385] , \[4400] ,
    \[4415] , \[4430] , \[4445] , \[4460] , \[4475] , \[4490] , \[4505] ,
    \[4520] , \[4535] , \[4550] , \[4565] , \[4580] , \[4595] , \[4610] ,
    \[4625] , \[4640] , \[4655] , \[4670] , \[4700] , \[4715] , \[4730] ,
    \[4745] , \[4760] , \[4775] , \[4790] , \[4805] , \[4820] , \[4835] ,
    \[4850] , \[4865] , \[4880] , \[4895] , \[4910] , \[4925] , \[4940] ,
    \[4955] , \[4970] , ppeakb_0_0_, ppeaka_7_7_, \[5015] , \[5030] ,
    ppeaks_4_4_, ppeakp_11_11_, \[5075] , \[5090] , \[5105] , \[5120] ,
    \[5135] , \[5150] , \[5165] , \[5180] , \[5195] , \[5210] , \[5225] ,
    \[5240] , \[5255] , \[5270] , \[5285] , \[5300] , \[5315] , \[5330] ,
    \[5345] , \[5360] , \[5375] , \[5390] , \[5405] , \[5420] , \[5435] ,
    \[5450] , \[5465] , \[5480] , \[5495] , \[5510] , \[5525] , \[5540] ,
    \[5555] , \[5570] , \[5600] , \[5615] , \[5630] , \[5645] , \[5660] ,
    \[5675] , ppeakb_10_10_, ppeaka_8_8_, \[5720] , ppeaks_14_14_,
    ppeaks_7_7_, ppeakp_12_12_, \[5780] , \[5795] , \[5810] , \[5825] ,
    \[5840] , \[5855] , \[5870] , \[5885] , \[5900] , \[5915] , \[5930] ,
    \[5945] , \[5960] , \[5975] , \[5990] , \[6005] , \[6020] , \[6035] ,
    \[6050] , \[6065] , \[6080] , \[6095] , \[6110] , \[6125] , \[6140] ,
    \[6155] , \[6170] , \[6185] , \[6200] , \[6215] , \[6230] , \[6245] ,
    \[6260] , \[6275] , \[6290] , \[6305] , \[6320] , \[6335] , \[6350] ,
    \[6365] , ppeakb_11_11_, ppeakb_2_2_, \[6410] , ppeaks_15_15_,
    ppeaks_6_6_, ppeakp_13_13_, \[6470] , \[6485] , \[6500] , \[6515] ,
    \[6530] , \[6545] , \[6560] , \[6575] , \[6590] , \[6605] , \[6620] ,
    \[6635] , \[6650] , \[6665] , \[6680] , \[6695] , \[6710] , \[6725] ,
    \[6740] , \[6755] , \[6770] , \[6785] , \[6815] , \[6830] , \[6845] ,
    \[6860] , \[6875] , \[6890] , \[6905] , \[6920] , \[6935] , \[6950] ,
    \[6965] , \[6980] , \[6995] , \[7010] , \[7025] , \[7055] ,
    ppeaks_12_12_, ppeaks_1_1_, ppeakp_3_3_, \[7115] , \[7130] , \[7145] ,
    \[7160] , \[7175] , \[7190] , \[7205] , \[7220] , \[7235] , \[7250] ,
    \[7265] , \[7280] , \[7295] , \[7310] , \[7325] , \[7340] , \[7355] ,
    \[7370] , \[7385] , \[7400] , \[7415] , \[7430] , \[7445] , \[7460] ,
    \[7475] , \[7490] , \[7505] , \[7520] , \[7535] , \[7550] , \[7565] ,
    \[7580] , \[7595] , \[7625] , \[7640] , \[7655] , \[7670] , \[7685] ,
    ppeaks_13_13_, ppeakp_7_7_, ppeakp_2_2_, \[7745] , \[7760] , \[7775] ,
    \[7790] , \[7805] , \[7820] , \[7835] , \[7850] , \[7865] , \[7880] ,
    \[7895] , \[7910] , \[7925] , \[7940] , \[7955] , \[7970] , \[8000] ,
    \[8015] , \[8030] , \[8045] , \[8060] , \[8075] , \[8090] , \[8105] ,
    \[8120] , \[8135] , \[8150] , \[8165] , \[8180] , \[8195] , \[8210] ,
    \[8225] , \[8240] , \[8255] , \[8285] , \[8300] , \[8315] , \[8330] ,
    ppeaks_3_3_, ppeakp_8_8_, ppeakp_1_1_, \[8390] , \[8405] , \[8420] ,
    \[8435] , \[8450] , \[8465] , \[8480] , \[8495] , \[8510] , \[8525] ,
    \[8540] , \[8555] , \[8570] , \[8585] , \[8600] , \[8615] , \[8630] ,
    \[8645] , \[8660] , \[8675] , \[8690] , \[8705] , \[8720] , \[8735] ,
    \[8750] , \[8765] , \[8780] , \[8810] , \[8825] , \[8840] , \[8855] ,
    \[8870] , \[8885] , \[8900] , \[8915] , \[8930] , \[8945] , \[8960] ,
    \[8975] , ppeaks_11_11_, ppeaks_2_2_, ppeakp_9_9_, ppeakp_0_0_,
    \[9050] , \[9065] , \[9080] , \[9095] , \[9110] , \[9125] , \[9140] ,
    \[9155] , \[9170] , \[9185] , \[9200] , \[9215] , \[9230] , \[9245] ,
    \[9260] , \[9275] , \[9290] , \[9305] , \[9320] , \[9335] , \[9350] ,
    \[9365] , \[9380] , \[9395] , \[9410] , \[9440] , \[9455] , \[9470] ,
    \[9485] , \[9500] , \[9515] , \[9530] , \[9545] , \[9560] , \[9575] ,
    \[9590] , \[9605] , \[9620] , \[9635] , \[9650] , \[9665] , \[9680] ,
    ppeaki_6_6_, \[9710] , \[9725] , \[9740] , \[9770] , \[9785] ,
    \[9800] , \[9815] , \[9830] , \[9845] , \[9860] , \[9875] , \[9890] ,
    \[9905] , \[9920] , \[9935] , \[9950] , \[9980] , \[9995] , \[10010] ,
    \[10025] , \[10040] , \[10055] , \[10070] , \[10085] , \[10100] ,
    \[10115] , \[10130] , \[10145] , \[10175] , \[10190] , \[10205] ,
    \[10220] , ppeaki_15_15_, ppeaki_4_4_, \[10265] , \[10280] , \[10310] ,
    \[10325] , \[10340] , \[10355] , \[10370] , \[10400] , \[10415] ,
    \[10430] , \[10445] , \[10460] , \[10475] , \[10490] , \[10505] ,
    ppeaki_14_14_, ppeaki_5_5_, \[10550] , \[10565] , \[10580] , \[10595] ,
    \[10610] , \[10625] , \[10655] , \[10670] , \[10685] , \[10700] ,
    \[10715] , \[10730] , \[10745] , \[10760] , \[10775] , \[10790] ,
    \[10805] , \[10820] , \[10850] , \[10865] , \[10880] , \[10895] ,
    \[10925] , \[10940] , \[10955] , \[10970] , \[10985] , \[11015] ,
    \[11030] , \[11045] , \[11060] , \[11075] , \[11090] , \[11120] ,
    \[11135] , \[11150] , \[11165] , \[11180] , \[11195] , \[11210] ,
    \[11225] , \[11240] , \[11255] , \[11270] , \[11285] , \[11300] ,
    \[11315] , \[11330] , \[11345] , \[11375] , \[11390] , \[11405] ,
    \[11420] , \[11435] , \[11450] , \[11465] , \[11480] , \[11495] ,
    \[11510] , \[11525] , \[11540] , \[11555] , \[11570] , \[11585] ,
    \[11600] , \[11615] , \[11630] , \[11645] , \[11660] , \[11675] ,
    \[11690] , \[11705] , \[11720] , \[11735] , \[11750] , \[11765] ,
    \[11780] , \[11795] , \[11810] , ppeaki_9_9_, ppeakb_14_14_, \[11885] ,
    \[11900] , \[11915] , \[11930] , ppeaki_8_8_, ppeakb_15_15_, \[12005] ,
    \[12020] , \[12035] , \[12050] , \[12065] , \[12080] , ppeaki_7_7_,
    \[12125] , \[12140] , \[12155] , \[12170] , \[12185] , \[12200] ,
    ppeakb_13_13_, \[12245] , \[12260] , \[12275] , ppeaki_13_13_,
    ppeaki_2_2_, \[12335] , \[12350] , \[12365] , \[12380] , \[12395] ,
    \[12410] , \[12425] , \[12440] , \[12455] , \[12470] , \[12485] ,
    ppeaki_12_12_, ppeaki_3_3_, \[12545] , \[12560] , \[12575] , \[12590] ,
    \[12605] , \[12620] , \[12635] , \[12650] , \[12665] , \[12680] ,
    \[12695] , ppeaki_11_11_, ppeaki_0_0_, \[12770] , \[12800] , \[12815] ,
    \[12830] , \[12845] , \[12860] , \[12875] , \[12890] , \[12905] ,
    \[12920] , \[12935] , ppeaki_10_10_, ppeaki_1_1_, \[13010] , \[13025] ,
    \[13040] , \[13055] , \[13070] , \[13085] , \[13100] , \[13115] ,
    \[13130] , \[13160] , \[13175] , ppeakb_4_4_, ppeaka_9_9_, \[13220] ,
    \[13235] , \[13250] , \[13265] , \[13280] , \[13295] , \[13310] ,
    \[13325] , \[13340] , \[13355] , \[13370] , \[13385] , \[13400] ,
    \[13415] , \[13430] , \[13445] , \[13460] , \[13475] , \[13490] ,
    \[13505] , ppeakb_5_5_, \[13550] , ppeakp_6_6_, \[13580] , \[13595] ,
    \[13610] , \[13625] , \[13640] , \[13655] , \[13670] , \[13685] ,
    \[13700] , \[13715] , \[13730] , \[13745] , \[13775] , \[13790] ,
    \[13805] , \[13820] , \[13835] , \[13850] , \[13865] , \[13880] ,
    \[13895] , ppeaka_11_11_, ppeaka_0_0_, ppeakp_5_5_, \[13955] ,
    \[13970] , \[13985] , \[14000] , \[14015] , \[14030] , \[14045] ,
    \[14060] , \[14075] , \[14090] , \[14105] , \[14120] , \[14135] ,
    \[14150] , \[14165] , \[14180] , \[14210] , \[14225] , \[14240] ,
    \[14255] , \[14270] , \[14285] , ppeakb_3_3_, ppeaka_10_10_,
    ppeaka_1_1_, ppeakp_4_4_, \[14360] , \[14375] , \[14390] , \[14405] ,
    \[14420] , \[14435] , \[14450] , \[14465] , \[14480] , \[14495] ,
    \[14510] , \[14525] , \[14540] , \[14555] , \[14570] , \[14585] ,
    \[14600] , \[14615] , \[14630] , \[14660] , \[14675] , \[14690] ,
    \[14705] , ppeakb_8_8_, ppeaka_13_13_, ppeaka_2_2_, \[14765] ,
    ppeaks_9_9_, ppeakp_14_14_, \[14810] , \[14825] , \[14840] , \[14855] ,
    \[14870] , \[14885] , \[14900] , \[14915] , \[14930] , \[14960] ,
    \[14975] , \[14990] , \[15005] , \[15020] , \[15035] , \[15050] ,
    \[15065] , \[15080] , ppeakb_9_9_, ppeaka_12_12_, ppeaka_3_3_,
    \[15140] , ppeaks_8_8_, ppeakp_15_15_, \[15185] , \[15200] , \[15215] ,
    \[15230] , \[15245] , \[15260] , \[15275] , \[15290] , \[15305] ,
    \[15320] , \[15335] , \[15350] , \[15365] , \[15380] , \[15395] ,
    \[15410] , \[15425] , \[15440] , ppeakb_6_6_, ppeaka_15_15_,
    ppeaka_4_4_, \[15500] , \[15515] , ppeaks_0_0_, \[15545] , \[15560] ,
    \[15575] , \[15590] , \[15605] , \[15620] , \[15635] , \[15650] ,
    \[15665] , \[15680] , \[15695] , \[15710] , \[15725] , \[15755] ,
    \[15770] , \[15785] , ppeakb_7_7_, ppeaka_14_14_, ppeaka_5_5_,
    \[15845] , \[15860] , ppeaks_10_10_, \[15890] , \[15905] , \[15920] ,
    \[15935] , \[15950] , \[15965] , \[15980] , \[15995] , \[16010] ,
    \[16025] , \[16040] , \[16055] , \[16070] , \[16085] , \[16100] ,
    paddress_8_8_, \[16907] , \[16920] , \[16933] , paddress_9_9_,
    \[16959] , \[16972] , \[16985] , \[16998] , \[17011] , \[17024] ,
    \[17037] , \[17050] , \[17063] , \[17076] , \[17089] , \[17102] ,
    \[17115] , \[17128] , \[17141] , \[17154] , \[17167] , \[17180] ,
    \[17193] , \[17206] , \[17219] , \[17232] , \[17245] , \[17258] ,
    \[17271] , \[17284] , \[17297] , \[17310] , \[17323] , \[17336] ,
    \[17349] , \[17362] , \[17375] , \[17388] , paddress_11_11_, \[17414] ,
    \[17427] , \[17453] , paddress_10_10_, \[17479] , \[17492] , \[17505] ,
    \[17518] , \[17531] , \[17544] , paddress_13_13_, \[17570] , \[17583] ,
    \[17596] , \[17609] , paddress_12_12_, \[17635] , \[17648] , \[17661] ,
    \[17674] , paddress_15_15_, \[17700] , \[17713] , paddress_14_14_,
    \[17739] , \[17752] , \[17765] , \[17778] , \[17791] , \[17804] ,
    \[17817] , pwr_0_0_, \[17843] , \[17856] , \[17869] , \[17882] ,
    prd_0_0_, \[17908] , \[17921] , \[17934] , \[17947] , \[17960] ,
    \[17973] , \[17986] , \[17999] , \[18012] , \[18025] , \[18038] , pdn,
    \[18064] , \[18077] , \[18090] , \[18103] , \[18116] , \[18129] ,
    \[18142] , \[18155] , \[18168] , \[18181] , \[18194] , \[18207] ,
    \[18220] , \[18233] , \[18246] , paddress_0_0_, piack_0_0_, \[18285] ,
    \[18298] , \[18311] , paddress_1_1_, \[18337] , \[18350] , \[18363] ,
    \[18376] , \[18389] , paddress_2_2_, \[18415] , \[18428] , \[18441] ,
    paddress_3_3_, \[18467] , \[18480] , \[18493] , \[18506] ,
    paddress_4_4_, paddress_5_5_, \[18545] , paddress_6_6_, \[18571] ,
    \[18584] , \[18597] , \[18610] , paddress_7_7_, \[18636] ;
  wire n3696_1, n3697, n3698, n3699, n3700, n3701_1, n3702, n3703, n3704,
    n3705, n3706_1, n3707, n3708, n3709, n3710, n3711_1, n3712, n3713,
    n3714, n3715, n3716_1, n3717, n3718, n3719, n3720, n3721_1, n3722,
    n3723, n3724, n3725, n3726_1, n3727, n3728, n3729, n3730, n3731_1,
    n3732, n3733, n3734, n3735, n3736_1, n3737, n3738, n3739, n3740,
    n3741_1, n3742, n3743, n3744, n3745, n3746_1, n3747, n3748, n3749,
    n3750_1, n3751, n3752, n3753, n3754_1, n3755, n3756, n3757, n3758_1,
    n3759, n3760, n3761, n3762, n3763_1, n3764, n3765, n3766, n3767,
    n3768_1, n3769, n3770, n3771, n3772_1, n3773, n3774, n3775, n3776,
    n3777_1, n3778, n3779, n3780, n3781, n3782_1, n3783, n3784, n3785,
    n3786, n3787_1, n3788, n3789, n3790, n3791, n3792_1, n3793, n3794,
    n3795, n3796, n3797_1, n3798, n3799, n3800, n3801, n3802_1, n3803,
    n3804, n3805, n3806, n3807_1, n3808, n3809, n3810, n3811, n3812_1,
    n3813, n3814, n3815, n3816, n3817_1, n3818, n3819, n3820, n3821,
    n3822_1, n3823, n3824, n3825, n3826, n3827_1, n3828, n3829, n3830,
    n3831, n3832_1, n3833, n3834, n3835, n3836, n3837_1, n3838, n3839,
    n3840, n3841, n3842_1, n3843, n3844, n3845, n3846, n3847_1, n3848,
    n3849, n3850, n3851, n3852_1, n3853, n3854, n3855, n3856_1, n3857,
    n3858, n3859, n3860_1, n3861, n3862, n3863, n3864_1, n3865, n3866,
    n3867, n3868, n3869_1, n3870, n3871, n3872, n3873, n3874_1, n3875,
    n3876, n3877, n3878_1, n3879, n3880, n3881, n3882, n3883_1, n3884,
    n3885, n3886, n3887, n3888_1, n3889, n3890, n3891, n3892, n3893_1,
    n3894, n3895, n3896, n3897, n3898_1, n3899, n3900, n3901, n3902,
    n3903_1, n3904, n3905, n3906, n3907, n3908_1, n3909, n3910, n3911,
    n3912, n3913_1, n3914, n3915, n3916, n3917, n3918_1, n3919, n3920,
    n3921, n3922, n3923_1, n3924, n3925, n3926, n3927, n3928_1, n3929,
    n3930, n3931, n3932, n3933_1, n3934, n3935, n3936, n3937, n3938_1,
    n3939, n3940, n3941, n3942, n3943_1, n3944, n3945, n3946, n3947,
    n3948_1, n3949, n3950, n3951, n3952, n3953_1, n3954, n3955, n3956,
    n3957_1, n3958, n3959, n3960, n3961, n3962_1, n3963, n3964, n3965,
    n3966, n3967_1, n3968, n3969, n3970, n3971, n3972_1, n3973, n3974,
    n3975, n3976_1, n3977, n3978, n3979, n3980, n3981_1, n3982, n3983,
    n3984, n3985, n3986_1, n3987, n3988, n3989, n3990, n3991_1, n3992,
    n3993, n3994, n3995, n3996_1, n3997, n3998, n3999, n4000, n4001_1,
    n4002, n4003, n4004, n4005, n4006_1, n4007, n4008, n4009, n4010,
    n4011_1, n4012, n4013, n4014, n4015, n4016_1, n4017, n4018, n4019,
    n4020, n4021_1, n4022, n4023, n4024, n4025, n4026_1, n4027, n4028,
    n4029, n4030, n4031_1, n4032, n4033, n4034, n4035, n4036_1, n4037,
    n4038, n4039, n4040, n4041_1, n4042, n4043, n4044, n4045, n4046_1,
    n4047, n4048, n4049, n4050, n4051_1, n4052, n4053, n4054, n4055,
    n4056_1, n4057, n4058, n4059, n4060, n4061_1, n4062, n4063, n4064,
    n4065, n4066_1, n4067, n4068, n4069, n4070, n4071_1, n4072, n4073,
    n4074, n4075, n4076_1, n4077, n4078, n4079, n4080, n4081_1, n4082,
    n4083, n4084, n4085, n4086_1, n4087, n4088, n4089, n4090, n4091_1,
    n4092, n4093, n4094, n4095, n4096_1, n4097, n4098, n4099, n4100,
    n4101_1, n4102, n4103, n4104, n4105, n4106_1, n4107, n4108, n4109,
    n4110, n4111_1, n4112, n4113, n4114, n4115, n4116_1, n4117, n4118,
    n4119, n4120, n4121_1, n4122, n4123, n4124, n4125, n4126_1, n4127,
    n4128, n4129, n4130, n4131_1, n4132, n4133, n4134, n4135, n4136_1,
    n4137, n4138, n4139, n4140, n4141_1, n4142, n4143, n4144, n4145,
    n4146_1, n4147, n4148, n4149, n4150_1, n4151, n4152, n4153, n4154,
    n4155_1, n4156, n4157, n4158, n4159, n4160_1, n4161, n4162, n4163,
    n4164, n4165_1, n4166, n4167, n4168, n4169_1, n4170, n4171, n4172,
    n4173, n4174_1, n4175, n4176, n4177, n4178, n4179_1, n4180, n4181,
    n4182, n4183, n4184_1, n4185, n4186, n4187, n4188, n4189_1, n4190,
    n4191, n4192, n4193, n4194_1, n4195, n4196, n4197, n4198, n4199_1,
    n4200, n4201, n4202, n4203_1, n4204, n4205, n4206, n4207, n4208_1,
    n4209, n4210, n4211, n4212, n4213_1, n4214, n4215, n4216, n4217,
    n4218_1, n4219, n4220, n4221, n4222, n4223_1, n4224, n4225, n4226,
    n4227_1, n4228, n4229, n4230, n4231, n4232_1, n4233, n4234, n4235,
    n4236, n4237_1, n4238, n4239, n4240, n4241, n4242_1, n4243, n4244,
    n4245, n4246, n4247_1, n4248, n4249, n4250, n4251_1, n4252, n4253,
    n4254, n4255, n4256_1, n4257, n4258, n4259, n4260, n4261_1, n4262,
    n4263, n4264, n4265_1, n4266, n4267, n4268, n4269, n4270_1, n4271,
    n4272, n4273, n4274, n4275_1, n4276, n4277, n4278, n4279, n4280_1,
    n4281, n4282, n4283, n4284, n4285_1, n4286, n4287, n4288, n4289,
    n4290_1, n4291, n4292, n4293, n4294, n4295_1, n4296, n4297, n4298,
    n4299, n4300_1, n4301, n4302, n4303, n4304_1, n4305, n4306, n4307,
    n4308, n4309_1, n4310, n4311, n4312, n4313, n4314_1, n4315, n4316,
    n4317, n4318, n4319_1, n4320, n4321, n4322, n4323, n4324_1, n4325,
    n4326, n4327, n4328_1, n4329, n4330, n4331, n4332, n4333_1, n4334,
    n4335, n4336, n4337, n4338_1, n4339, n4340, n4341, n4342, n4343_1,
    n4344, n4345, n4346, n4347, n4348_1, n4349, n4350, n4351, n4352,
    n4353_1, n4354, n4355, n4356, n4357, n4358_1, n4359, n4360, n4361,
    n4362, n4363_1, n4364, n4365, n4366, n4367, n4368_1, n4369, n4370,
    n4371, n4372, n4373_1, n4374, n4375, n4376, n4377, n4378_1, n4379,
    n4380, n4381, n4382, n4383_1, n4384, n4385, n4386, n4387_1, n4388,
    n4389, n4390, n4391, n4392_1, n4393, n4394, n4395, n4396, n4397_1,
    n4398, n4399, n4400, n4401, n4402_1, n4403, n4404, n4405, n4406,
    n4407_1, n4408, n4409, n4410, n4411, n4412_1, n4413, n4414, n4415,
    n4416, n4417_1, n4418, n4419, n4420, n4421, n4422_1, n4423, n4424,
    n4425, n4426, n4427_1, n4428, n4429, n4430, n4431, n4432_1, n4433,
    n4434, n4435, n4436, n4437_1, n4438, n4439, n4440, n4441, n4442_1,
    n4443, n4444, n4445, n4446, n4447_1, n4448, n4449, n4450, n4451,
    n4452_1, n4453, n4454, n4455, n4456, n4457_1, n4458, n4459, n4460,
    n4461, n4462_1, n4463, n4464, n4465, n4466_1, n4467, n4468, n4469,
    n4470_1, n4471, n4472, n4473, n4474, n4475_1, n4476, n4477, n4478,
    n4479, n4480_1, n4481, n4482, n4483, n4484, n4485_1, n4486, n4487,
    n4488, n4489_1, n4490, n4491, n4492, n4493, n4494_1, n4495, n4496,
    n4497, n4498, n4499_1, n4500, n4501, n4502, n4503, n4504_1, n4505,
    n4506, n4507, n4508, n4509_1, n4510, n4511, n4512, n4513, n4514_1,
    n4515, n4516, n4517, n4518_1, n4519, n4520, n4521, n4522, n4523_1,
    n4524, n4525, n4526, n4527, n4528_1, n4529, n4530, n4531, n4532,
    n4533_1, n4534, n4535, n4536, n4537_1, n4538, n4539, n4540, n4541,
    n4542_1, n4543, n4544, n4545, n4546, n4547_1, n4548, n4549, n4550,
    n4551, n4552_1, n4553, n4554, n4555, n4556, n4557_1, n4558, n4559,
    n4560, n4561_1, n4562, n4563, n4564, n4565_1, n4566, n4567, n4568,
    n4569, n4570_1, n4571, n4572, n4573, n4574_1, n4575, n4576, n4577,
    n4578, n4579_1, n4580, n4581, n4582, n4583, n4584_1, n4585, n4586,
    n4587, n4588, n4589_1, n4590, n4591, n4592, n4593, n4594_1, n4595,
    n4596, n4597, n4598_1, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
    n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
    n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
    n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
    n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
    n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
    n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
    n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
    n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
    n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
    n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
    n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
    n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
    n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
    n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
    n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
    n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
    n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
    n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
    n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
    n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
    n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
    n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
    n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
    n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
    n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
    n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
    n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
    n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
    n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
    n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
    n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
    n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
    n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
    n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
    n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
    n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
    n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
    n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
    n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
    n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
    n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
    n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
    n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
    n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
    n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
    n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
    n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
    n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
    n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
    n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
    n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
    n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
    n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
    n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
    n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
    n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
    n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
    n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
    n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
    n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
    n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
    n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
    n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
    n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
    n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
    n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
    n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
    n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
    n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
    n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
    n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
    n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
    n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
    n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
    n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
    n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
    n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
    n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
    n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
    n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
    n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
    n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
    n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
    n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
    n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
    n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
    n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
    n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
    n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
    n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
    n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
    n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
    n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
    n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
    n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
    n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
    n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
    n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
    n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
    n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
    n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
    n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
    n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
    n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
    n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
    n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
    n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
    n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
    n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
    n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
    n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
    n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
    n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
    n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
    n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
    n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
    n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
    n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
    n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
    n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
    n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
    n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
    n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
    n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
    n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
    n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
    n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
    n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
    n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
    n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
    n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
    n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
    n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
    n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
    n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
    n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
    n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
    n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
    n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
    n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
    n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
    n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
    n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
    n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
    n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
    n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
    n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
    n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
    n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
    n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
    n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
    n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
    n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
    n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
    n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
    n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
    n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
    n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
    n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
    n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
    n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
    n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
    n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
    n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
    n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
    n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
    n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
    n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
    n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
    n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
    n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
    n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
    n6326, n6327, n6328, n6329, n6330, n6331, n6332, n273, n278, n282,
    n286, n290, n295, n300, n304, n308, n313, n318, n323, n328, n333, n338,
    n343, n348, n353, n358, n363, n368, n373, n378, n383, n388, n393, n398,
    n403, n408, n413, n418, n423, n428, n433, n438, n443, n448, n453, n458,
    n463, n468, n473, n478, n483, n488, n493, n498, n503, n508, n513, n517,
    n521, n526, n531, n535, n539, n544, n549, n554, n559, n564, n569, n574,
    n579, n584, n589, n594, n599, n604, n609, n614, n619, n624, n629, n634,
    n639, n644, n649, n654, n659, n664, n669, n674, n679, n684, n689, n694,
    n699, n704, n709, n714, n719, n724, n729, n734, n739, n743, n747, n752,
    n756, n760, n764, n769, n774, n779, n784, n789, n794, n799, n804, n809,
    n814, n819, n824, n829, n834, n839, n844, n849, n854, n859, n864, n869,
    n874, n879, n884, n889, n894, n899, n904, n909, n914, n919, n924, n929,
    n934, n939, n944, n949, n954, n959, n964, n968, n972, n977, n981, n985,
    n989, n994, n999, n1004, n1009, n1014, n1019, n1024, n1029, n1034,
    n1039, n1044, n1049, n1054, n1059, n1064, n1069, n1074, n1079, n1084,
    n1089, n1094, n1099, n1104, n1109, n1114, n1119, n1124, n1129, n1134,
    n1139, n1144, n1149, n1154, n1159, n1164, n1169, n1174, n1179, n1183,
    n1187, n1191, n1196, n1201, n1206, n1211, n1216, n1221, n1226, n1231,
    n1236, n1241, n1246, n1251, n1256, n1261, n1266, n1271, n1276, n1281,
    n1286, n1291, n1296, n1301, n1306, n1311, n1316, n1321, n1326, n1331,
    n1336, n1341, n1346, n1351, n1356, n1361, n1366, n1371, n1376, n1381,
    n1385, n1389, n1393, n1398, n1403, n1408, n1413, n1418, n1423, n1428,
    n1433, n1438, n1443, n1448, n1453, n1458, n1463, n1468, n1473, n1478,
    n1483, n1488, n1493, n1498, n1503, n1508, n1513, n1518, n1523, n1528,
    n1533, n1538, n1543, n1548, n1553, n1558, n1563, n1568, n1573, n1578,
    n1583, n1587, n1591, n1595, n1600, n1605, n1610, n1615, n1620, n1625,
    n1630, n1635, n1640, n1645, n1650, n1655, n1660, n1665, n1670, n1675,
    n1680, n1685, n1690, n1695, n1700, n1705, n1710, n1715, n1720, n1725,
    n1730, n1735, n1740, n1745, n1750, n1755, n1760, n1765, n1770, n1775,
    n1780, n1785, n1790, n1794, n1798, n1802, n1806, n1811, n1816, n1821,
    n1826, n1831, n1836, n1841, n1846, n1851, n1856, n1861, n1866, n1871,
    n1876, n1881, n1886, n1891, n1896, n1901, n1906, n1911, n1916, n1921,
    n1926, n1931, n1936, n1941, n1946, n1951, n1956, n1961, n1966, n1971,
    n1976, n1981, n1986, n1991, n1996, n2001, n2006, n2011, n2016, n2020,
    n2025, n2030, n2035, n2040, n2045, n2050, n2055, n2060, n2065, n2070,
    n2075, n2080, n2085, n2090, n2095, n2100, n2105, n2110, n2115, n2120,
    n2125, n2130, n2135, n2140, n2145, n2150, n2155, n2160, n2165, n2170,
    n2175, n2180, n2184, n2188, n2193, n2198, n2203, n2208, n2213, n2218,
    n2223, n2228, n2233, n2238, n2243, n2248, n2253, n2258, n2263, n2267,
    n2271, n2276, n2281, n2286, n2291, n2296, n2301, n2306, n2311, n2316,
    n2321, n2326, n2331, n2336, n2341, n2346, n2351, n2356, n2361, n2366,
    n2371, n2376, n2381, n2386, n2391, n2396, n2401, n2406, n2411, n2416,
    n2421, n2426, n2431, n2436, n2441, n2446, n2451, n2456, n2461, n2466,
    n2471, n2476, n2481, n2486, n2491, n2496, n2501, n2506, n2511, n2516,
    n2521, n2526, n2531, n2536, n2541, n2546, n2551, n2556, n2561, n2566,
    n2571, n2576, n2581, n2586, n2591, n2596, n2601, n2606, n2611, n2616,
    n2621, n2626, n2631, n2636, n2641, n2646, n2651, n2656, n2661, n2666,
    n2670, n2674, n2679, n2684, n2689, n2694, n2698, n2702, n2707, n2712,
    n2717, n2722, n2727, n2732, n2736, n2741, n2746, n2751, n2756, n2761,
    n2766, n2770, n2775, n2780, n2785, n2789, n2793, n2798, n2803, n2808,
    n2813, n2818, n2823, n2828, n2833, n2838, n2843, n2848, n2852, n2856,
    n2861, n2866, n2871, n2876, n2881, n2886, n2891, n2896, n2901, n2906,
    n2911, n2915, n2919, n2924, n2929, n2934, n2939, n2944, n2949, n2954,
    n2959, n2964, n2969, n2974, n2978, n2982, n2987, n2992, n2997, n3002,
    n3007, n3012, n3017, n3022, n3027, n3032, n3037, n3041, n3045, n3050,
    n3055, n3060, n3065, n3070, n3075, n3080, n3085, n3090, n3095, n3100,
    n3105, n3110, n3115, n3120, n3125, n3130, n3135, n3140, n3145, n3149,
    n3154, n3158, n3163, n3168, n3173, n3178, n3183, n3188, n3193, n3198,
    n3203, n3208, n3213, n3218, n3223, n3228, n3233, n3238, n3243, n3248,
    n3253, n3258, n3263, n3267, n3271, n3275, n3280, n3285, n3290, n3295,
    n3300, n3305, n3310, n3315, n3320, n3325, n3330, n3335, n3340, n3345,
    n3350, n3355, n3360, n3365, n3370, n3375, n3380, n3385, n3389, n3393,
    n3397, n3401, n3406, n3411, n3416, n3421, n3426, n3431, n3436, n3441,
    n3446, n3451, n3456, n3461, n3466, n3471, n3476, n3481, n3486, n3491,
    n3496, n3501, n3506, n3511, n3516, n3520, n3524, n3528, n3533, n3537,
    n3541, n3546, n3551, n3556, n3561, n3566, n3571, n3576, n3581, n3586,
    n3591, n3596, n3601, n3606, n3611, n3616, n3621, n3626, n3631, n3635,
    n3639, n3643, n3648, n3652, n3656, n3661, n3666, n3671, n3676, n3681,
    n3686, n3691, n3696, n3701, n3706, n3711, n3716, n3721, n3726, n3731,
    n3736, n3741, n3746, n3750, n3754, n3758, n3763, n3768, n3772, n3777,
    n3782, n3787, n3792, n3797, n3802, n3807, n3812, n3817, n3822, n3827,
    n3832, n3837, n3842, n3847, n3852, n3856, n3860, n3864, n3869, n3874,
    n3878, n3883, n3888, n3893, n3898, n3903, n3908, n3913, n3918, n3923,
    n3928, n3933, n3938, n3943, n3948, n3953, n3957, n3962, n3967, n3972,
    n3976, n3981, n3986, n3991, n3996, n4001, n4006, n4011, n4016, n4021,
    n4026, n4031, n4036, n4041, n4046, n4051, n4056, n4061, n4066, n4071,
    n4076, n4081, n4086, n4091, n4096, n4101, n4106, n4111, n4116, n4121,
    n4126, n4131, n4136, n4141, n4146, n4150, n4155, n4160, n4165, n4169,
    n4174, n4179, n4184, n4189, n4194, n4199, n4203, n4208, n4213, n4218,
    n4223, n4227, n4232, n4237, n4242, n4247, n4251, n4256, n4261, n4265,
    n4270, n4275, n4280, n4285, n4290, n4295, n4300, n4304, n4309, n4314,
    n4319, n4324, n4328, n4333, n4338, n4343, n4348, n4353, n4358, n4363,
    n4368, n4373, n4378, n4383, n4387, n4392, n4397, n4402, n4407, n4412,
    n4417, n4422, n4427, n4432, n4437, n4442, n4447, n4452, n4457, n4462,
    n4466, n4470, n4475, n4480, n4485, n4489, n4494, n4499, n4504, n4509,
    n4514, n4518, n4523, n4528, n4533, n4537, n4542, n4547, n4552, n4557,
    n4561, n4565, n4570, n4574, n4579, n4584, n4589, n4594, n4598;
  assign pdata_8_8_ = \[17882]  ? \[16959]  : tin_pdata_8_8_;
  assign pdata_0_0_ = \[17479]  ? \[18337]  : tin_pdata_0_0_;
  assign pdata_7_7_ = \[17869]  ? \[16907]  : tin_pdata_7_7_;
  assign pdata_2_2_ = \[18181]  ? \[17323]  : tin_pdata_2_2_;
  assign pdata_9_9_ = \[18571]  ? \[17765]  : tin_pdata_9_9_;
  assign pdata_1_1_ = \[18116]  ? \[17258]  : tin_pdata_1_1_;
  assign pdata_4_4_ = \[18038]  ? \[17193]  : tin_pdata_4_4_;
  assign pdata_10_10_ = \[17011]  ? \[17921]  : tin_pdata_10_10_;
  assign pdata_3_3_ = \[17960]  ? \[17128]  : tin_pdata_3_3_;
  assign pdata_6_6_ = \[17934]  ? \[17063]  : tin_pdata_6_6_;
  assign pdata_15_15_ = \[17947]  ? \[17076]  : tin_pdata_15_15_;
  assign pdata_11_11_ = \[17336]  ? \[18194]  : tin_pdata_11_11_;
  assign pdata_14_14_ = \[18584]  ? \[17778]  : tin_pdata_14_14_;
  assign pdata_12_12_ = \[17141]  ? \[17973]  : tin_pdata_12_12_;
  assign pdata_5_5_ = \[17908]  ? \[16998]  : tin_pdata_5_5_;
  assign pdata_13_13_ = \[18350]  ? \[17492]  : tin_pdata_13_13_;
  assign n273 = n5632 | (pdata_2_2_ & n3696_1);
  assign n278 = n5690 | n5687 | n5688;
  assign n282 = n5694 | n5691 | n5692;
  assign n286 = n5700 | n5698 | n5699;
  assign n290 = n5703 | n5596 | n5597;
  assign n295 = n5704 | n5593 | n5594;
  assign n300 = n5715 | n5713 | n5714;
  assign n304 = n5573 | n5575 | n5576 | n5727;
  assign n308 = n5572 | (pdata_0_0_ & n3703);
  assign n313 = n5571 | (pdata_11_11_ & n3703);
  assign n318 = ~preset & (n3792_1 ? pdata_6_6_ : \[4385] );
  assign n323 = n5570 | (pdata_1_1_ & n3705);
  assign n328 = n5569 | (pdata_12_12_ & n3705);
  assign n333 = ~preset & (n3817_1 ? pdata_7_7_ : \[4430] );
  assign n338 = ~preset & (n3817_1 ? pdata_2_2_ : \[4445] );
  assign n343 = ~preset & (n3817_1 ? pdata_13_13_ : \[4460] );
  assign n348 = n5568 | (pdata_8_8_ & n3708);
  assign n353 = n5567 | (pdata_3_3_ & n4504);
  assign n358 = n5566 | (pdata_14_14_ & n4504);
  assign n363 = n5564 | n5565;
  assign n368 = n5562 | n5563;
  assign n373 = n5560 | n5561;
  assign n378 = ~preset & (n3813 ? pdata_5_5_ : \[4565] );
  assign n383 = ~preset & (n3813 ? pdata_0_0_ : \[4580] );
  assign n388 = ~preset & (n3813 ? pdata_11_11_ : \[4595] );
  assign n393 = n5559 | (pdata_6_6_ & n3711_1);
  assign n398 = (n4160 & n3712) | (\[4625]  & n3713);
  assign n403 = (n4160 & n3714) | (\[4640]  & n3713);
  assign n408 = n5481 | n5482;
  assign n413 = n5480 | (\[4670]  & n3707);
  assign n418 = n5478 | n5479;
  assign n423 = n5477 | (\[4715]  & n3717);
  assign n428 = (\[4730]  & n3717) | (n3718 & n3719);
  assign n433 = n5461 | (n4547 & n3720);
  assign n438 = n5460 | (\[4760]  & n3710);
  assign n443 = n5459 | (\[4775]  & n3710);
  assign n448 = n5457 | n5458;
  assign n453 = (n3712 & n3723) | (\[4805]  & n3722);
  assign n458 = (n3714 & n3723) | (\[4820]  & n3722);
  assign n463 = ~preset & (n3825 ? n3724 : \[4835] );
  assign n468 = n5378 | (n3726_1 & n3727);
  assign n473 = (n3728 & n3730) | (\[4865]  & n3729);
  assign n478 = n5342 | (n3730 & (~n3930 ^ n3931));
  assign n483 = n5341 | (n3731_1 & n3732);
  assign n488 = (n3733 & n3735) | (\[4910]  & n3734);
  assign n493 = (\[4925]  & n3722) | (n3723 & n3736_1);
  assign n498 = (\[4940]  & n3722) | (n3723 & n3737);
  assign n503 = (n3724 & n3739) | (\[4955]  & n3738);
  assign n508 = n5340 | (pdata_1_1_ & n3696_1);
  assign n513 = n5862 | n5859 | n5860;
  assign n517 = n5868 | n5866 | n5867;
  assign n521 = n5869 | n5319 | n5320;
  assign n526 = n5870 | n5316 | n5317;
  assign n531 = n5876 | n5874 | n5875;
  assign n535 = n5298 | n5300 | n5301 | n5878;
  assign n539 = n5297 | (pdata_1_1_ & n3703);
  assign n544 = n5296 | (pdata_10_10_ & n3703);
  assign n549 = n5295 | (pdata_2_2_ & n3705);
  assign n554 = n5294 | (pdata_11_11_ & n3705);
  assign n559 = ~preset & (n3817_1 ? pdata_8_8_ : \[5135] );
  assign n564 = ~preset & (n3817_1 ? pdata_1_1_ : \[5150] );
  assign n569 = ~preset & (n3817_1 ? pdata_14_14_ : \[5165] );
  assign n574 = n5293 | (pdata_7_7_ & n3708);
  assign n579 = n5292 | (pdata_4_4_ & n4504);
  assign n584 = n5291 | (pdata_13_13_ & n4504);
  assign n589 = n5289 | n5290;
  assign n594 = n5287 | n5288;
  assign n599 = n5285 | n5286;
  assign n604 = ~preset & (n3813 ? pdata_4_4_ : \[5270] );
  assign n609 = ~preset & (n3813 ? pdata_1_1_ : \[5285] );
  assign n614 = ~preset & (n3813 ? pdata_10_10_ : \[5300] );
  assign n619 = n5284 | (pdata_7_7_ & n3711_1);
  assign n624 = n5283 | (n4160 & (n3893_1 ^ n3894));
  assign n629 = n5282 | (\[5345]  & n3713);
  assign n634 = n5281 | (n3714 & n3715);
  assign n639 = n5280 | (\[5375]  & n3707);
  assign n644 = n5279 | (n3716_1 & (n3893_1 ^ n3894));
  assign n649 = n5278 | (n3716_1 & n3720);
  assign n654 = n5277 | (\[5420]  & n3717);
  assign n659 = (\[5435]  & n3717) | (n3718 & n3740);
  assign n664 = n5275 | n5276;
  assign n669 = n5274 | (n4106 & n3720);
  assign n674 = (n3709 & n3740) | (\[5480]  & n3710);
  assign n679 = n5273 | (n3721_1 & n3741_1);
  assign n684 = n5272 | (\[5510]  & n3722);
  assign n689 = n5271 | (\[5525]  & n3722);
  assign n694 = ~preset & (n3825 ? n3742 : \[5540] );
  assign n699 = n5270 | (n3727 & n3743);
  assign n704 = (\[5570]  & n3729) | (n3730 & n3733);
  assign n709 = n5269 | (n3732 & n3744);
  assign n714 = (n3728 & n3735) | (\[5615]  & n3734);
  assign n719 = n5268 | (n4081 & n3744);
  assign n724 = (\[5645]  & n3722) | (n3723 & n3745);
  assign n729 = (\[5660]  & n3738) | (n3739 & n3746_1);
  assign n734 = n5267 | (pdata_0_0_ & n3696_1);
  assign n739 = n5882 | n5879 | n5880;
  assign n743 = n5888 | n5886 | n5887;
  assign n747 = n5889 | n5246 | n5247;
  assign n752 = n5895 | n5893 | n5894;
  assign n756 = n5901 | n5899 | n5900;
  assign n760 = n5214 | n5216 | n5217 | n5903;
  assign n764 = n5213 | (pdata_2_2_ & n3703);
  assign n769 = ~preset & (n3792_1 ? pdata_4_4_ : \[5795] );
  assign n774 = ~preset & (n3792_1 ? pdata_8_8_ : \[5810] );
  assign n779 = ~preset & (n3817_1 ? pdata_9_9_ : \[5825] );
  assign n784 = ~preset & (n3817_1 ? pdata_4_4_ : \[5840] );
  assign n789 = ~preset & (n3817_1 ? pdata_11_11_ : \[5855] );
  assign n794 = n5212 | (pdata_6_6_ & n3708);
  assign n799 = n5211 | (pdata_5_5_ & n4504);
  assign n804 = n5209 | n5210;
  assign n809 = n5207 | n5208;
  assign n814 = n5205 | n5206;
  assign n819 = n5203 | n5204;
  assign n824 = ~preset & (n3813 ? pdata_7_7_ : \[5960] );
  assign n829 = ~preset & (n3813 ? pdata_14_14_ : \[5975] );
  assign n834 = ~preset & (n3813 ? pdata_9_9_ : \[5990] );
  assign n839 = n5202 | (pdata_8_8_ & n3711_1);
  assign n844 = (n4160 & n3747) | (\[6020]  & n3713);
  assign n849 = n5201 | (\[6035]  & n3713);
  assign n854 = n5199 | n5200;
  assign n859 = n5198 | (\[6065]  & n3707);
  assign n864 = (n3706_1 & n3740) | (\[6080]  & n3707);
  assign n869 = n5196 | n5197;
  assign n874 = (\[6110]  & n3717) | (n3718 & n3741_1);
  assign n879 = n5195 | (n4547 & (n3893_1 ^ n3894));
  assign n884 = n5193 | n5194;
  assign n889 = n5191 | n5192;
  assign n894 = n5190 | (\[6170]  & n3710);
  assign n899 = n5188 | n5189;
  assign n904 = (\[6200]  & n3722) | (n3723 & n3747);
  assign n909 = (\[6215]  & n3722) | (n3723 & n3740);
  assign n914 = ~preset & (n3825 ? n3728 : \[6230] );
  assign n919 = n5187 | (n3742 & n3748);
  assign n924 = n5186 | (n3727 & n3736_1);
  assign n929 = n5185 | (n3732 & n3749);
  assign n934 = n5184 | (n3732 & n3743);
  assign n939 = (\[6305]  & n3734) | (n3735 & n3736_1);
  assign n944 = n5183 | (n3750_1 & (~n3930 ^ n3931));
  assign n949 = (\[6335]  & n3722) | (n3723 & n3752);
  assign n954 = (\[6350]  & n3738) | (n3739 & n3744);
  assign n959 = n5182 | (n3739 & (~n3930 ^ n3931));
  assign n964 = n5907 | n5904 | n5905;
  assign n968 = n5911 | n5908 | n5909;
  assign n972 = n5912 | n5159 | n5160;
  assign n977 = n5918 | n5916 | n5917;
  assign n981 = n5924 | n5922 | n5923;
  assign n985 = n5127 | n5129 | n5130 | n5926;
  assign n989 = n5126 | (pdata_12_12_ & n3703);
  assign n994 = ~preset & (n3792_1 ? pdata_5_5_ : \[6485] );
  assign n999 = ~preset & (n3792_1 ? pdata_7_7_ : \[6500] );
  assign n1004 = ~preset & (n3817_1 ? pdata_10_10_ : \[6515] );
  assign n1009 = ~preset & (n3817_1 ? pdata_3_3_ : \[6530] );
  assign n1014 = ~preset & (n3817_1 ? pdata_12_12_ : \[6545] );
  assign n1019 = n5125 | (pdata_5_5_ & n3708);
  assign n1024 = n5124 | (pdata_6_6_ & n4504);
  assign n1029 = n5123 | (pdata_15_15_ & n4504);
  assign n1034 = n5121 | n5122;
  assign n1039 = n5119 | n5120;
  assign n1044 = ~preset & (n3813 ? pdata_6_6_ : \[6635] );
  assign n1049 = ~preset & (n3813 ? pdata_15_15_ : \[6650] );
  assign n1054 = ~preset & (n3813 ? pdata_8_8_ : \[6665] );
  assign n1059 = n5118 | (pdata_9_9_ & n3711_1);
  assign n1064 = n5117 | (\[6695]  & n3713);
  assign n1069 = n5116 | (\[6710]  & n3713);
  assign n1074 = n5115 | (n3715 & n3740);
  assign n1079 = (n3706_1 & n3741_1) | (\[6740]  & n3707);
  assign n1084 = (n3706_1 & n3719) | (\[6755]  & n3707);
  assign n1089 = n5113 | n5114;
  assign n1094 = n5112 | (\[6785]  & n3717);
  assign n1099 = n5110 | n5111;
  assign n1104 = n5108 | n5109;
  assign n1109 = (n3709 & n3747) | (\[6845]  & n3710);
  assign n1114 = (n3709 & n3714) | (\[6860]  & n3710);
  assign n1119 = n5107 | (\[6875]  & n3722);
  assign n1124 = n5106 | (\[6890]  & n3722);
  assign n1129 = ~preset & (n3825 ? n3746_1 : \[6905] );
  assign n1134 = n5105 | (n3744 & n3748);
  assign n1139 = n5104 | (n3727 & n3749);
  assign n1144 = n5103 | (n3732 & n3736_1);
  assign n1149 = n5102 | (n3726_1 & n3732);
  assign n1154 = (\[6980]  & n3734) | (n3735 & n3753);
  assign n1159 = (n3746_1 & n3750_1) | (\[6995]  & n3751);
  assign n1164 = n5101 | (n3723 & (~n3930 ^ n3931));
  assign n1169 = (\[7025]  & n3738) | (n3739 & n3742);
  assign n1174 = n5927 | n5098 | n5099;
  assign n1179 = n5933 | n5931 | n5932;
  assign n1183 = n5939 | n5937 | n5938;
  assign n1187 = n5066 | n5068 | n5069 | n5941;
  assign n1191 = n5065 | (pdata_7_7_ & n3703);
  assign n1196 = ~preset & (n3792_1 ? pdata_2_2_ : \[7130] );
  assign n1201 = ~preset & (n3817_1 ? pdata_11_11_ : \[7145] );
  assign n1206 = ~preset & (n3817_1 ? pdata_6_6_ : \[7160] );
  assign n1211 = n5064 | (pdata_1_1_ & n3708);
  assign n1216 = n5063 | (pdata_12_12_ & n3708);
  assign n1221 = n5062 | (pdata_15_15_ & n3708);
  assign n1226 = n5061 | (pdata_10_10_ & n4504);
  assign n1231 = n5059 | n5060;
  assign n1236 = n5057 | n5058;
  assign n1241 = ~preset & (n3813 ? pdata_9_9_ : \[7265] );
  assign n1246 = ~preset & (n3813 ? pdata_4_4_ : \[7280] );
  assign n1251 = ~preset & (n3813 ? pdata_15_15_ : \[7295] );
  assign n1256 = n5056 | (pdata_2_2_ & n3711_1);
  assign n1261 = n5055 | (pdata_13_13_ & n3711_1);
  assign n1266 = n5054 | (\[7340]  & n3713);
  assign n1271 = n5053 | (n3715 & n3719);
  assign n1276 = (n3706_1 & n3720) | (\[7370]  & n3707);
  assign n1281 = n5052 | (n3716_1 & n3747);
  assign n1286 = n5051 | (n3716_1 & n3740);
  assign n1291 = n5050 | (n3718 & (n3893_1 ^ n3894));
  assign n1296 = n5049 | (\[7430]  & n3717);
  assign n1301 = n5047 | n5048;
  assign n1306 = n5046 | (n4106 & n3714);
  assign n1311 = (n3709 & n3741_1) | (\[7475]  & n3710);
  assign n1316 = n5045 | (n3721_1 & (n3893_1 ^ n3894));
  assign n1321 = n5043 | n5044;
  assign n1326 = n5042 | (\[7520]  & n3722);
  assign n1331 = ~preset & (n3825 ? n3753 : \[7535] );
  assign n1336 = n5041 | (n3731_1 & n3748);
  assign n1341 = n5040 | (n3727 & n3733);
  assign n1346 = n5039 | (n3727 & n3752);
  assign n1351 = (\[7595]  & n3729) | (n3730 & n3744);
  assign n1356 = (n3724 & n3750_1) | (\[7625]  & n3751);
  assign n1361 = n5038 | (n4081 & n3749);
  assign n1366 = n5037 | (n4081 & n3743);
  assign n1371 = (\[7670]  & n3722) | (n3723 & n3746_1);
  assign n1376 = n5942 | n5034 | n5035;
  assign n1381 = n5948 | n5946 | n5947;
  assign n1385 = n5016 | n5018 | n5019 | n5950;
  assign n1389 = n5012 | n5014 | n5015 | n5952;
  assign n1393 = n5011 | (pdata_6_6_ & n3703);
  assign n1398 = ~preset & (n3792_1 ? pdata_3_3_ : \[7760] );
  assign n1403 = ~preset & (n3817_1 ? pdata_12_12_ : \[7775] );
  assign n1408 = ~preset & (n3817_1 ? pdata_5_5_ : \[7790] );
  assign n1413 = n5010 | (pdata_2_2_ & n3708);
  assign n1418 = n5009 | (pdata_11_11_ & n3708);
  assign n1423 = n5008 | (pdata_0_0_ & n4504);
  assign n1428 = n5007 | (pdata_9_9_ & n4504);
  assign n1433 = n5005 | n5006;
  assign n1438 = n5003 | n5004;
  assign n1443 = ~preset & (n3813 ? pdata_8_8_ : \[7895] );
  assign n1448 = ~preset & (n3813 ? pdata_5_5_ : \[7910] );
  assign n1453 = ~preset & (n3813 ? pdata_14_14_ : \[7925] );
  assign n1458 = n5002 | (pdata_3_3_ & n3711_1);
  assign n1463 = n5001 | (pdata_12_12_ & n3711_1);
  assign n1468 = (n4160 & n3720) | (\[7970]  & n3713);
  assign n1473 = n5000 | (\[8000]  & n3707);
  assign n1478 = n4998 | n4999;
  assign n1483 = n4996 | n4997;
  assign n1488 = (n3712 & n3718) | (\[8045]  & n3717);
  assign n1493 = n4995 | (\[8060]  & n3717);
  assign n1498 = n4994 | (n4547 & n3741_1);
  assign n1503 = n4992 | n4993;
  assign n1508 = n4991 | (\[8105]  & n3710);
  assign n1513 = n4990 | (n3712 & n3721_1);
  assign n1518 = n4988 | n4989;
  assign n1523 = n4987 | (n3719 & n3721_1);
  assign n1528 = ~preset & (n3825 ? n3733 : \[8165] );
  assign n1533 = n4986 | (n3726_1 & n3748);
  assign n1538 = n4985 | (n3727 & n3753);
  assign n1543 = n4984 | (n3727 & (~n3930 ^ n3931));
  assign n1548 = (\[8225]  & n3729) | (n3730 & n3742);
  assign n1553 = (\[8240]  & n3734) | (n3735 & n3749);
  assign n1558 = (n3742 & n3750_1) | (\[8255]  & n3751);
  assign n1563 = n4983 | (n4081 & n3737);
  assign n1568 = (\[8300]  & n3722) | (n3723 & n3728);
  assign n1573 = (\[8315]  & n3738) | (n3739 & n3752);
  assign n1578 = n5953 | n4980 | n4981;
  assign n1583 = n5959 | n5957 | n5958;
  assign n1587 = n4962 | n4964 | n4965 | n5961;
  assign n1591 = n4958 | n4960 | n4961 | n5963;
  assign n1595 = n4957 | (pdata_9_9_ & n3703);
  assign n1600 = ~preset & (n3792_1 ? pdata_0_0_ : \[8405] );
  assign n1605 = ~preset & (n3817_1 ? pdata_13_13_ : \[8420] );
  assign n1610 = ~preset & (n3817_1 ? pdata_8_8_ : \[8435] );
  assign n1615 = ~preset & (n3817_1 ? pdata_15_15_ : \[8450] );
  assign n1620 = n4956 | (pdata_10_10_ & n3708);
  assign n1625 = n4955 | (pdata_1_1_ & n4504);
  assign n1630 = n4954 | (pdata_12_12_ & n4504);
  assign n1635 = n4952 | n4953;
  assign n1640 = ~preset & (n3813 ? pdata_0_0_ : \[8525] );
  assign n1645 = ~preset & (n3813 ? pdata_11_11_ : \[8540] );
  assign n1650 = ~preset & (n3813 ? pdata_2_2_ : \[8555] );
  assign n1655 = ~preset & (n3813 ? pdata_13_13_ : \[8570] );
  assign n1660 = n4951 | (pdata_4_4_ & n3711_1);
  assign n1665 = n4950 | (pdata_15_15_ & n3711_1);
  assign n1670 = (n4160 & n3741_1) | (\[8615]  & n3713);
  assign n1675 = n4949 | (n3706_1 & (n3893_1 ^ n3894));
  assign n1680 = n4948 | (\[8645]  & n3707);
  assign n1685 = n4947 | (n3712 & n3716_1);
  assign n1690 = n4946 | (n3714 & n3716_1);
  assign n1695 = n4945 | (\[8690]  & n3717);
  assign n1700 = n4944 | (\[8705]  & n3717);
  assign n1705 = n4943 | (n4547 & n3747);
  assign n1710 = n4942 | (n4106 & n3740);
  assign n1715 = n4941 | (\[8750]  & n3710);
  assign n1720 = (n3709 & n3719) | (\[8765]  & n3710);
  assign n1725 = n4940 | (n3720 & n3721_1);
  assign n1730 = n4939 | (\[8810]  & n3722);
  assign n1735 = n4938 | (n3743 & n3748);
  assign n1740 = n4937 | (n3727 & n3746_1);
  assign n1745 = n4936 | (n3727 & n3737);
  assign n1750 = (n3724 & n3730) | (\[8870]  & n3729);
  assign n1755 = (\[8885]  & n3729) | (n3730 & n3745);
  assign n1760 = n4935 | (n3732 & n3742);
  assign n1765 = (n3744 & n3750_1) | (\[8915]  & n3751);
  assign n1770 = n4934 | (n4081 & n3753);
  assign n1775 = n4933 | (n4081 & n3731_1);
  assign n1780 = (\[8960]  & n3722) | (n3723 & n3733);
  assign n1785 = (n3728 & n3739) | (\[8975]  & n3738);
  assign n1790 = n5969 | n5967 | n5968;
  assign n1794 = n5975 | n5973 | n5974;
  assign n1798 = n4901 | n4903 | n4904 | n5977;
  assign n1802 = n4897 | n4899 | n4900 | n5979;
  assign n1806 = n4896 | (pdata_8_8_ & n3703);
  assign n1811 = ~preset & (n3792_1 ? pdata_1_1_ : \[9065] );
  assign n1816 = ~preset & (n3817_1 ? pdata_14_14_ : \[9080] );
  assign n1821 = ~preset & (n3817_1 ? pdata_7_7_ : \[9095] );
  assign n1826 = n4895 | (pdata_0_0_ & n3708);
  assign n1831 = n4894 | (pdata_9_9_ & n3708);
  assign n1836 = n4893 | (pdata_2_2_ & n4504);
  assign n1841 = n4892 | (pdata_11_11_ & n4504);
  assign n1846 = n4890 | n4891;
  assign n1851 = ~preset & (n3813 ? pdata_1_1_ : \[9185] );
  assign n1856 = ~preset & (n3813 ? pdata_10_10_ : \[9200] );
  assign n1861 = ~preset & (n3813 ? pdata_3_3_ : \[9215] );
  assign n1866 = ~preset & (n3813 ? pdata_12_12_ : \[9230] );
  assign n1871 = n4889 | (pdata_5_5_ & n3711_1);
  assign n1876 = n4888 | (pdata_14_14_ & n3711_1);
  assign n1881 = n4887 | (\[9275]  & n3713);
  assign n1886 = (n3706_1 & n3712) | (\[9290]  & n3707);
  assign n1891 = n4886 | (\[9305]  & n3707);
  assign n1896 = n4884 | n4885;
  assign n1901 = n4882 | n4883;
  assign n1906 = (\[9350]  & n3717) | (n3718 & n3747);
  assign n1911 = (n3714 & n3718) | (\[9365]  & n3717);
  assign n1916 = n4880 | n4881;
  assign n1921 = n4879 | (n4106 & n3719);
  assign n1926 = n4878 | (\[9410]  & n3710);
  assign n1931 = n4876 | n4877;
  assign n1936 = n4875 | (n3723 & (n3893_1 ^ n3894));
  assign n1941 = (n3720 & n3723) | (\[9470]  & n3722);
  assign n1946 = ~preset & (n3825 ? n3736_1 : \[9485] );
  assign n1951 = n4874 | (n3737 & n3748);
  assign n1956 = n4873 | (n3727 & n3728);
  assign n1961 = n4872 | (n3727 & n3745);
  assign n1966 = (\[9545]  & n3729) | (n3730 & n3746_1);
  assign n1971 = (\[9560]  & n3729) | (n3730 & n3752);
  assign n1976 = n4871 | (n3724 & n3732);
  assign n1981 = (n3731_1 & n3750_1) | (\[9590]  & n3751);
  assign n1986 = n4870 | (n4081 & n3736_1);
  assign n1991 = n4869 | (n4081 & n3726_1);
  assign n1996 = (\[9635]  & n3722) | (n3723 & n3753);
  assign n2001 = (\[9650]  & n3722) | (n3723 & n3743);
  assign n2006 = n4868 | (pdata_1_1_ & n3754_1);
  assign n2011 = n4867 | (pdata_12_12_ & n3754_1);
  assign n2016 = n4865 | (n3755 & n3756) | n4866;
  assign n2020 = ~preset & (n3813 ? pdata_2_2_ : \[9710] );
  assign n2025 = n4864 | (\[9725]  & n3707);
  assign n2030 = n4863 | (\[9740]  & n3707);
  assign n2035 = n4862 | (\[9770]  & n3710);
  assign n2040 = n4860 | n4861;
  assign n2045 = n4859 | (n3745 & n3748);
  assign n2050 = n4858 | (n3727 & n3742);
  assign n2055 = (\[9830]  & n3729) | (n3730 & n3736_1);
  assign n2060 = (\[9845]  & n3729) | (n3730 & n3737);
  assign n2065 = (n3726_1 & n3750_1) | (\[9860]  & n3751);
  assign n2070 = n4857 | (n4081 & n3728);
  assign n2075 = n4856 | (n4081 & (~n3930 ^ n3931));
  assign n2080 = (\[9905]  & n3722) | (n3723 & n3731_1);
  assign n2085 = (n3733 & n3739) | (\[9920]  & n3738);
  assign n2090 = n4855 | (pdata_0_0_ & n3754_1);
  assign n2095 = n4854 | (pdata_6_6_ & n3757);
  assign n2100 = ~preset & (n3813 ? pdata_12_12_ : \[9980] );
  assign n2105 = (n3706_1 & n3747) | (\[9995]  & n3707);
  assign n2110 = (n3706_1 & n3714) | (\[10010]  & n3707);
  assign n2115 = n4853 | (n3709 & (n3893_1 ^ n3894));
  assign n2120 = (n3709 & n3720) | (\[10040]  & n3710);
  assign n2125 = n4852 | (n3721_1 & n3740);
  assign n2130 = n4851 | (n3748 & n3752);
  assign n2135 = n4850 | (n3724 & n3727);
  assign n2140 = (\[10100]  & n3729) | (n3730 & n3753);
  assign n2145 = (\[10115]  & n3729) | (n3730 & n3743);
  assign n2150 = (n3743 & n3750_1) | (\[10130]  & n3751);
  assign n2155 = n4849 | (n4081 & n3733);
  assign n2160 = (\[10175]  & n3722) | (n3723 & n3744);
  assign n2165 = (\[10190]  & n3738) | (n3739 & n3745);
  assign n2170 = n4848 | (pdata_10_10_ & n3754_1);
  assign n2175 = n4847 | (pdata_5_5_ & n3757);
  assign n2180 = n4846 | (\[12200]  & (n5627 | n5628));
  assign n2184 = n4844 | (n3756 & n3758_1) | n4845;
  assign n2188 = ~preset & (n3813 ? pdata_6_6_ : \[10265] );
  assign n2193 = n4842 | n4843;
  assign n2198 = (n3709 & n3712) | (\[10310]  & n3710);
  assign n2203 = n4840 | n4841;
  assign n2208 = n4838 | n4839;
  assign n2213 = n4837 | (n3748 & (~n3930 ^ n3931));
  assign n2218 = n4836 | (n3727 & n3731_1);
  assign n2223 = (n3726_1 & n3730) | (\[10400]  & n3729);
  assign n2228 = (n3737 & n3750_1) | (\[10415]  & n3751);
  assign n2233 = n4835 | (n4081 & n3724);
  assign n2238 = n4834 | (n4081 & n3745);
  assign n2243 = (\[10460]  & n3722) | (n3723 & n3742);
  assign n2248 = n4833 | (pdata_2_2_ & n3754_1);
  assign n2253 = n4832 | (pdata_11_11_ & n3754_1);
  assign n2258 = n4831 | (pdata_4_4_ & n3757);
  assign n2263 = n4830 | (\[12080]  & (n5627 | n5628));
  assign n2267 = n4828 | (n3756 & n3759) | n4829;
  assign n2271 = n4827 | (pdata_0_0_ & n3711_1);
  assign n2276 = n4826 | (n3716_1 & n3741_1);
  assign n2281 = n4825 | (n3716_1 & n3719);
  assign n2286 = n4824 | (\[10595]  & n3710);
  assign n2291 = n4823 | (n3721_1 & n3747);
  assign n2296 = n4822 | (n3714 & n3721_1);
  assign n2301 = n4821 | (n3727 & n3744);
  assign n2306 = (\[10670]  & n3729) | (n3730 & n3749);
  assign n2311 = (\[10685]  & n3729) | (n3730 & n3731_1);
  assign n2316 = (n3745 & n3750_1) | (\[10700]  & n3751);
  assign n2321 = n4820 | (n4081 & n3746_1);
  assign n2326 = n4819 | (n4081 & n3752);
  assign n2331 = (\[10745]  & n3722) | (n3723 & n3724);
  assign n2336 = n4818 | (pdata_13_13_ & n3696_1);
  assign n2341 = n4817 | (pdata_8_8_ & n3754_1);
  assign n2346 = n4816 | (pdata_3_3_ & n3757);
  assign n2351 = n4815 | (pdata_1_1_ & n3760);
  assign n2356 = n4814 | (pdata_12_12_ & n3760);
  assign n2361 = n4813 | (pdata_10_10_ & n3711_1);
  assign n2366 = n4812 | (\[10865]  & n3717);
  assign n2371 = n4810 | n4811;
  assign n2376 = n4809 | (\[10895]  & n3722);
  assign n2381 = ~preset & (n3825 ? n3726_1 : \[10925] );
  assign n2386 = n4808 | (n3732 & n3753);
  assign n2391 = n4807 | (n3732 & n3745);
  assign n2396 = (\[10970]  & n3734) | (n3735 & n3742);
  assign n2401 = (n3750_1 & n3752) | (\[10985]  & n3751);
  assign n2406 = (n3726_1 & n3739) | (\[11015]  & n3738);
  assign n2411 = n4806 | (pdata_12_12_ & n3696_1);
  assign n2416 = n4805 | (pdata_9_9_ & n3754_1);
  assign n2421 = n4804 | (pdata_2_2_ & n3757);
  assign n2426 = n4803 | (pdata_7_7_ & n3757);
  assign n2431 = n4802 | (pdata_13_13_ & n3760);
  assign n2436 = n4801 | (\[11120]  & n3713);
  assign n2441 = (\[11135]  & n3717) | (n3718 & n3720);
  assign n2446 = n4800 | (n4547 & n3712);
  assign n2451 = (\[11165]  & n3722) | (n3723 & n3741_1);
  assign n2456 = (n3719 & n3723) | (\[11180]  & n3722);
  assign n2461 = n4799 | (n3732 & n3733);
  assign n2466 = n4798 | (n3732 & n3737);
  assign n2471 = (\[11225]  & n3734) | (n3735 & n3744);
  assign n2476 = n4797 | (n4081 & n3742);
  assign n2481 = (\[11255]  & n3738) | (n3739 & n3749);
  assign n2486 = (n3731_1 & n3739) | (\[11270]  & n3738);
  assign n2491 = n4796 | (pdata_15_15_ & n3696_1);
  assign n2496 = n4795 | (pdata_6_6_ & n3754_1);
  assign n2501 = n4794 | (pdata_1_1_ & n3757);
  assign n2506 = n4793 | (pdata_8_8_ & n3757);
  assign n2511 = n4792 | (pdata_3_3_ & n3760);
  assign n2516 = (n4160 & n3740) | (\[11375]  & n3713);
  assign n2521 = n4790 | n4791;
  assign n2526 = n4789 | (\[11405]  & n3722);
  assign n2531 = ~preset & (n3825 ? n3744 : \[11420] );
  assign n2536 = n4788 | (n3728 & n3732);
  assign n2541 = n4787 | (n3732 & (~n3930 ^ n3931));
  assign n2546 = (\[11465]  & n3734) | (n3735 & n3746_1);
  assign n2551 = (\[11480]  & n3722) | (n3723 & n3749);
  assign n2556 = (n3736_1 & n3739) | (\[11495]  & n3738);
  assign n2561 = (n3737 & n3739) | (\[11510]  & n3738);
  assign n2566 = n4786 | (pdata_14_14_ & n3696_1);
  assign n2571 = n4785 | (pdata_7_7_ & n3754_1);
  assign n2576 = n4784 | (pdata_0_0_ & n3757);
  assign n2581 = n4783 | (pdata_9_9_ & n3757);
  assign n2586 = n4782 | (pdata_2_2_ & n3760);
  assign n2591 = n4781 | (pdata_11_11_ & n3760);
  assign n2596 = n4780 | (n4547 & n3714);
  assign n2601 = ~preset & (n3825 ? n3749 : \[11630] );
  assign n2606 = ~preset & (n3825 ? n3731_1 : \[11645] );
  assign n2611 = n4779 | (n3732 & n3746_1);
  assign n2616 = n4778 | (n3732 & n3752);
  assign n2621 = (n3724 & n3735) | (\[11690]  & n3734);
  assign n2626 = (\[11705]  & n3722) | (n3723 & n3726_1);
  assign n2631 = (\[11720]  & n3738) | (n3739 & n3753);
  assign n2636 = (\[11735]  & n3738) | (n3739 & n3743);
  assign n2641 = n4777 | (pdata_9_9_ & n3696_1);
  assign n2646 = n4776 | (pdata_4_4_ & n3754_1);
  assign n2651 = n4775 | (pdata_15_15_ & n3754_1);
  assign n2656 = n4774 | (pdata_10_10_ & n3757);
  assign n2661 = n4773 | (pdata_5_5_ & n3760);
  assign n2666 = n4771 | (n3756 & n3761) | n4772;
  assign n2670 = n5983 | n5980 | n5981;
  assign n2674 = n4760 | (pdata_5_5_ & n3754_1);
  assign n2679 = n4759 | (pdata_14_14_ & n3754_1);
  assign n2684 = n4758 | (pdata_11_11_ & n3757);
  assign n2689 = n4757 | (pdata_4_4_ & n3760);
  assign n2694 = n4755 | (n3756 & n3762) | n4756;
  assign n2698 = n4753 | n5985 | n5986 | n5987;
  assign n2702 = (n3736_1 & n3764) | (\[12005]  & n3763_1);
  assign n2707 = n4743 | (pdata_11_11_ & n3696_1);
  assign n2712 = n4742 | (pdata_13_13_ & n3754_1);
  assign n2717 = n4741 | (pdata_12_12_ & n3757);
  assign n2722 = n4740 | (pdata_7_7_ & n3760);
  assign n2727 = n4739 | (pdata_14_14_ & n3760);
  assign n2732 = n4737 | (n3756 & n3765) | n4738;
  assign n2736 = (n3743 & n3764) | (\[12125]  & n3763_1);
  assign n2741 = n4736 | (pdata_10_10_ & n3696_1);
  assign n2746 = n4735 | (pdata_3_3_ & n3754_1);
  assign n2751 = n4734 | (pdata_13_13_ & n3757);
  assign n2756 = n4733 | (pdata_6_6_ & n3760);
  assign n2761 = n4732 | (pdata_15_15_ & n3760);
  assign n2766 = n4730 | n5989 | n5990 | n5991;
  assign n2770 = (n3728 & n3750_1) | (\[12245]  & n3751);
  assign n2775 = n4720 | (pdata_14_14_ & n3757);
  assign n2780 = n4719 | (pdata_9_9_ & n3760);
  assign n2785 = n4718 | (\[11090]  & (n5627 | n5628));
  assign n2789 = n4716 | (n3756 & n3766) | n4717;
  assign n2793 = n4715 | (\[12335]  & n3704);
  assign n2798 = n4713 | n4714;
  assign n2803 = n4712 | (n3962 & n3719);
  assign n2808 = n4711 | (n3736_1 & n3767);
  assign n2813 = n4710 | (n3737 & n3767);
  assign n2818 = n4709 | (n3724 & n3748);
  assign n2823 = n4708 | (n3735 & (~n3930 ^ n3931));
  assign n2828 = (n3731_1 & n3764) | (\[12440]  & n3763_1);
  assign n2833 = (n3733 & n3750_1) | (\[12455]  & n3751);
  assign n2838 = n4707 | (pdata_15_15_ & n3757);
  assign n2843 = n4706 | (pdata_8_8_ & n3760);
  assign n2848 = n4705 | (\[10820]  & (n5627 | n5628));
  assign n2852 = n4703 | (n3756 & n3768_1) | n4704;
  assign n2856 = n4701 | n4702;
  assign n2861 = (n4427 & n3741_1) | (\[12560]  & n3704);
  assign n2866 = n4700 | (n3962 & n3747);
  assign n2871 = n4698 | n4699;
  assign n2876 = n4697 | (n3749 & n3767);
  assign n2881 = n4696 | (n3745 & n3767);
  assign n2886 = n4695 | (n3746_1 & n3748);
  assign n2891 = (\[12650]  & n3734) | (n3735 & n3752);
  assign n2896 = (n3726_1 & n3764) | (\[12665]  & n3763_1);
  assign n2901 = (n3750_1 & n3753) | (\[12680]  & n3751);
  assign n2906 = n4694 | (pdata_0_0_ & n3760);
  assign n2911 = n4692 | (n3756 & n3769) | n4693;
  assign n2915 = n4690 | (n3756 & n3770) | n4691;
  assign n2919 = n4688 | n4689;
  assign n2924 = n4686 | n4687;
  assign n2929 = n4684 | n4685;
  assign n2934 = n4682 | n4683;
  assign n2939 = n4681 | (n3733 & n3767);
  assign n2944 = n4680 | (n3726_1 & n3767);
  assign n2949 = n4679 | (n3728 & n3748);
  assign n2954 = (n3749 & n3764) | (\[12890]  & n3763_1);
  assign n2959 = (n3742 & n3764) | (\[12905]  & n3763_1);
  assign n2964 = (n3736_1 & n3750_1) | (\[12920]  & n3751);
  assign n2969 = n4678 | (pdata_10_10_ & n3760);
  assign n2974 = n4676 | (n3756 & n3771) | n4677;
  assign n2978 = n4674 | (n3756 & n3772_1) | n4675;
  assign n2982 = n4672 | n4673;
  assign n2987 = n4671 | (n3715 & (n3893_1 ^ n3894));
  assign n2992 = n4670 | (n3715 & n3720);
  assign n2997 = n4668 | n4669;
  assign n3002 = n4667 | (n3962 & n3740);
  assign n3007 = n4666 | (n4106 & n3741_1);
  assign n3012 = n4665 | (n3753 & n3767);
  assign n3017 = n4664 | (n3743 & n3767);
  assign n3022 = n4663 | (n3733 & n3748);
  assign n3027 = (n3744 & n3764) | (\[13160]  & n3763_1);
  assign n3032 = (n3749 & n3750_1) | (\[13175]  & n3751);
  assign n3037 = n5995 | n5992 | n5993;
  assign n3041 = n6001 | n5999 | n6000;
  assign n3045 = n4644 | (pdata_3_3_ & n3703);
  assign n3050 = n4643 | (pdata_14_14_ & n3703);
  assign n3055 = ~preset & (n3792_1 ? pdata_14_14_ : \[13250] );
  assign n3060 = n4642 | (pdata_9_9_ & n3705);
  assign n3065 = ~preset & (n3817_1 ? pdata_4_4_ : \[13280] );
  assign n3070 = n4640 | n4641;
  assign n3075 = n4638 | n4639;
  assign n3080 = n4636 | n4637;
  assign n3085 = n4634 | n4635;
  assign n3090 = (n4427 & n3747) | (\[13355]  & n3704);
  assign n3095 = (n4427 & n3740) | (\[13370]  & n3704);
  assign n3100 = n4632 | n4633;
  assign n3105 = n4631 | (n3962 & (n3893_1 ^ n3894));
  assign n3110 = n4629 | n4630;
  assign n3115 = n4627 | n4628;
  assign n3120 = ~preset & (n3825 ? n3752 : \[13445] );
  assign n3125 = n4626 | (n3744 & n3767);
  assign n3130 = n4625 | (n3748 & n3753);
  assign n3135 = (\[13490]  & n3734) | (n3735 & n3743);
  assign n3140 = (n3746_1 & n3764) | (\[13505]  & n3763_1);
  assign n3145 = n6005 | n6002 | n6003;
  assign n3149 = n6006 | n4612 | n4613;
  assign n3154 = n4608 | n4610 | n4611 | n6008;
  assign n3158 = n4607 | (pdata_15_15_ & n3703);
  assign n3163 = ~preset & (n3792_1 ? pdata_13_13_ : \[13595] );
  assign n3168 = n4606 | (pdata_10_10_ & n3705);
  assign n3173 = ~preset & (n3817_1 ? pdata_3_3_ : \[13625] );
  assign n3178 = n4604 | n4605;
  assign n3183 = n4602 | n4603;
  assign n3188 = n4600 | n4601;
  assign n3193 = n4598_1 | n4599;
  assign n3198 = n4597 | (\[13700]  & n3713);
  assign n3203 = n4596 | (\[13715]  & n3704);
  assign n3208 = (n4427 & n3719) | (\[13730]  & n3704);
  assign n3213 = n4594_1 | n4595;
  assign n3218 = n4593 | (n3962 & n3714);
  assign n3223 = n4591 | n4592;
  assign n3228 = ~preset & (n3825 ? n3745 : \[13805] );
  assign n3233 = n4590 | (n3731_1 & n3767);
  assign n3238 = n4589_1 | (n3736_1 & n3748);
  assign n3243 = (n3726_1 & n3735) | (\[13850]  & n3734);
  assign n3248 = (n3724 & n3764) | (\[13865]  & n3763_1);
  assign n3253 = n4588 | (n3764 & (~n3930 ^ n3931));
  assign n3258 = n4587 | (pdata_8_8_ & n3696_1);
  assign n3263 = n6014 | n6012 | n6013;
  assign n3267 = n6018 | n4577 | n6016;
  assign n3271 = n4560 | n4562 | n4563 | n6020;
  assign n3275 = n4559 | (pdata_5_5_ & n3703);
  assign n3280 = n4558 | (pdata_0_0_ & n3705);
  assign n3285 = n4557_1 | (pdata_7_7_ & n3705);
  assign n3290 = ~preset & (n3817_1 ? pdata_2_2_ : \[14000] );
  assign n3295 = n4556 | (pdata_13_13_ & n3708);
  assign n3300 = n4555 | (pdata_8_8_ & n4504);
  assign n3305 = n4553 | n4554;
  assign n3310 = n4551 | n4552_1;
  assign n3315 = n4549 | n4550;
  assign n3320 = n4548 | (pdata_11_11_ & n3711_1);
  assign n3325 = n4547_1 | (\[14105]  & n3704);
  assign n3330 = (n4427 & n3714) | (\[14120]  & n3704);
  assign n3335 = n4546 | (n3715 & n3741_1);
  assign n3340 = n4544 | n4545;
  assign n3345 = n4543 | (n3962 & n3720);
  assign n3350 = n4542_1 | (n4106 & n3747);
  assign n3355 = n4541 | (n3724 & n3767);
  assign n3360 = n4540 | (n3748 & n3749);
  assign n3365 = (\[14240]  & n3734) | (n3735 & n3745);
  assign n3370 = (n3733 & n3764) | (\[14255]  & n3763_1);
  assign n3375 = (n3752 & n3764) | (\[14270]  & n3763_1);
  assign n3380 = n4539 | (pdata_7_7_ & n3696_1);
  assign n3385 = n4537_1 | n6022 | n6023 | n6024;
  assign n3389 = n6028 | n4527 | n6026;
  assign n3393 = n6032 | n4513 | n6030;
  assign n3397 = n4496 | n4498 | n4499_1 | n6034;
  assign n3401 = n4495 | (pdata_4_4_ & n3703);
  assign n3406 = n4494_1 | (pdata_13_13_ & n3703);
  assign n3411 = ~preset & (n3792_1 ? pdata_15_15_ : \[14390] );
  assign n3416 = n4493 | (pdata_8_8_ & n3705);
  assign n3421 = ~preset & (n3817_1 ? pdata_1_1_ : \[14420] );
  assign n3426 = n4492 | (pdata_14_14_ & n3708);
  assign n3431 = n4491 | (pdata_7_7_ & n4504);
  assign n3436 = n4489_1 | n4490;
  assign n3441 = n4487 | n4488;
  assign n3446 = n4485_1 | n4486;
  assign n3451 = n4484 | (pdata_1_1_ & n3711_1);
  assign n3456 = n4483 | (\[14525]  & n3704);
  assign n3461 = n4482 | (\[14540]  & n3704);
  assign n3466 = n4480_1 | n4481;
  assign n3471 = n4479 | (n3962 & n3712);
  assign n3476 = n4477 | n4478;
  assign n3481 = n4475_1 | n4476;
  assign n3486 = n4474 | (n3725 & (~n3930 ^ n3931));
  assign n3491 = n4473 | (n3742 & n3767);
  assign n3496 = (\[14660]  & n3734) | (n3735 & n3737);
  assign n3501 = (n3728 & n3764) | (\[14675]  & n3763_1);
  assign n3506 = (n3745 & n3764) | (\[14690]  & n3763_1);
  assign n3511 = n4472 | (pdata_6_6_ & n3696_1);
  assign n3516 = n4470_1 | n6036 | n6037 | n6038;
  assign n3520 = n6044 | n6042 | n6043;
  assign n3524 = n6048 | n4451 | n6046;
  assign n3528 = n6049 | n4435 | n4436;
  assign n3533 = n6055 | n6053 | n6054;
  assign n3537 = n4417_1 | n4419 | n4420 | n6057;
  assign n3541 = ~preset & (n3792_1 ? pdata_10_10_ : \[14810] );
  assign n3546 = n4416 | (pdata_5_5_ & n3705);
  assign n3551 = ~preset & (n3817_1 ? pdata_0_0_ : \[14840] );
  assign n3556 = ~preset & (n3817_1 ? pdata_9_9_ : \[14855] );
  assign n3561 = n4415 | (pdata_4_4_ & n3708);
  assign n3566 = n4413 | n4414;
  assign n3571 = n4411 | n4412_1;
  assign n3576 = n4409 | n4410;
  assign n3581 = ~preset & (n3813 ? pdata_7_7_ : \[14930] );
  assign n3586 = n4408 | (\[14960]  & n3704);
  assign n3591 = n4406 | n4407_1;
  assign n3596 = n4404 | n4405;
  assign n3601 = n4402_1 | n4403;
  assign n3606 = n4401 | (n4106 & n3712);
  assign n3611 = n4400 | (n3728 & n3767);
  assign n3616 = n4399 | (n3767 & (~n3930 ^ n3931));
  assign n3621 = (n3737 & n3764) | (\[15065]  & n3763_1);
  assign n3626 = n4398 | (pdata_5_5_ & n3696_1);
  assign n3631 = n4396 | n6059 | n6060 | n6061;
  assign n3635 = n6067 | n6065 | n6066;
  assign n3639 = n6071 | n4378_1 | n6069;
  assign n3643 = n6072 | n4362 | n4363_1;
  assign n3648 = n6078 | n6076 | n6077;
  assign n3652 = n4344 | n4346 | n4347 | n6080;
  assign n3656 = ~preset & (n3792_1 ? pdata_9_9_ : \[15185] );
  assign n3661 = n4343_1 | (pdata_6_6_ & n3705);
  assign n3666 = n4342 | (pdata_15_15_ & n3705);
  assign n3671 = ~preset & (n3817_1 ? pdata_10_10_ : \[15230] );
  assign n3676 = n4341 | (pdata_3_3_ & n3708);
  assign n3681 = n4339 | n4340;
  assign n3686 = n4337 | n4338_1;
  assign n3691 = n4335 | n4336;
  assign n3696 = ~preset & (n3813 ? pdata_13_13_ : \[15305] );
  assign n3701 = (n4160 & n3719) | (\[15320]  & n3713);
  assign n3706 = n4334 | (\[15335]  & n3704);
  assign n3711 = n4333_1 | (n3715 & n3747);
  assign n3716 = n4331 | n4332;
  assign n3721 = n4330 | (n4106 & (n3893_1 ^ n3894));
  assign n3726 = n4329 | (n3746_1 & n3767);
  assign n3731 = n4328_1 | (n3752 & n3767);
  assign n3736 = (n3753 & n3764) | (\[15425]  & n3763_1);
  assign n3741 = n4327 | (pdata_4_4_ & n3696_1);
  assign n3746 = n4325 | n6082 | n6083 | n6084;
  assign n3750 = n4315 | n6085 | n6086 | n6087;
  assign n3754 = n6091 | n4302 | n6089;
  assign n3758 = n6092 | n4286 | n4287;
  assign n3763 = n6093 | n4283 | n4284;
  assign n3768 = n6099 | n6097 | n6098;
  assign n3772 = ~preset & (n3792_1 ? pdata_12_12_ : \[15545] );
  assign n3777 = n4268 | (pdata_3_3_ & n3705);
  assign n3782 = n4267 | (pdata_14_14_ & n3705);
  assign n3787 = ~preset & (n3817_1 ? pdata_5_5_ : \[15590] );
  assign n3792 = ~preset & (n3817_1 ? pdata_0_0_ : \[15605] );
  assign n3797 = n4265_1 | n4266;
  assign n3802 = n4263 | n4264;
  assign n3807 = n4261_1 | n4262;
  assign n3812 = ~preset & (n3813 ? pdata_3_3_ : \[15665] );
  assign n3817 = (n4427 & n3712) | (\[15680]  & n3704);
  assign n3822 = n4260 | (\[15695]  & n3704);
  assign n3827 = n4258 | n4259;
  assign n3832 = n4257 | (n4547 & n3719);
  assign n3837 = ~preset & (n3825 ? n3737 : \[15755] );
  assign n3842 = (n3731_1 & n3735) | (\[15770]  & n3734);
  assign n3847 = n4256_1 | (pdata_3_3_ & n3696_1);
  assign n3852 = n6103 | n6100 | n6101;
  assign n3856 = n6109 | n6107 | n6108;
  assign n3860 = n6113 | n4237_1 | n6111;
  assign n3864 = n6114 | n4221 | n4222;
  assign n3869 = n6115 | n4218_1 | n4219;
  assign n3874 = n6121 | n6119 | n6120;
  assign n3878 = ~preset & (n3792_1 ? pdata_11_11_ : \[15890] );
  assign n3883 = n4203_1 | (pdata_4_4_ & n3705);
  assign n3888 = n4202 | (pdata_13_13_ & n3705);
  assign n3893 = ~preset & (n3817_1 ? pdata_6_6_ : \[15935] );
  assign n3898 = ~preset & (n3817_1 ? pdata_15_15_ : \[15950] );
  assign n3903 = n4200 | n4201;
  assign n3908 = n4198 | n4199_1;
  assign n3913 = n4196 | n4197;
  assign n3918 = n4194_1 | n4195;
  assign n3923 = n4193 | (n4427 & (n3893_1 ^ n3894));
  assign n3928 = (n4427 & n3720) | (\[16040]  & n3704);
  assign n3933 = n4192 | (n3712 & n3715);
  assign n3938 = n4191 | (n4547 & n3740);
  assign n3943 = n4190 | (n3962 & n3741_1);
  assign n3948 = ~preset & (n3825 ? n3743 : \[16100] );
  assign n3953 = n6140 | n6141;
  assign n3957 = n4175 | n6142;
  assign n3962 = n3876 & n3798 & ~preset & ~\[16920] ;
  assign n3967 = n4141 | (n3798 & n3803 & n6143);
  assign n3972 = n6149 | n6150;
  assign n3976 = n4163 | n6151;
  assign n3981 = \[16972]  & ~preset & ~\[16920] ;
  assign n3986 = ~\[18389]  & ~preset & \[16985] ;
  assign n3991 = n4161 | n6152;
  assign n3996 = ~preset & (\[17011]  | n3858 | n3859);
  assign n4001 = ~preset & ~pdn;
  assign n4006 = ~preset & ~\[17102]  & (\[17037]  | \[18025] );
  assign n4011 = \[17115]  & ~preset & ~\[17050] ;
  assign n4016 = n4159 | n6153;
  assign n4021 = n4157 | n6154;
  assign n4026 = \[17089]  & ~preset & ~pdn;
  assign n4031 = ~\[17102]  & ~preset & \[17037] ;
  assign n4036 = n4011 | (n3798 & n3826 & n6155);
  assign n4041 = n4155_1 | n6156;
  assign n4046 = ~preset & (\[17141]  | n3858 | n3859);
  assign n4051 = \[17154]  & ~preset & ~\[17102] ;
  assign n4056 = n3819 & n3798 & ~preset & ~\[17167] ;
  assign n4061 = n4081 | (n3798 & n3827_1 & n6157);
  assign n4066 = n4153 | n6158;
  assign n4071 = n4096 | (n3798 & n3808 & n6159);
  assign n4076 = \[17219]  & ~preset & ~\[17050] ;
  assign n4081 = ~\[17232]  & ~preset & \[17180] ;
  assign n4086 = ~preset & \[17245]  & (~n3798 | ~n3811);
  assign n4091 = n4151 | n6160;
  assign n4096 = ~\[17271]  & ~preset & \[17206] ;
  assign n4101 = n4504 | (n3798 & n3802_1 & n6161);
  assign n4106 = n3812_1 & n3798 & ~preset & ~\[17297] ;
  assign n4111 = ~\[17388]  & ~preset & \[17310] ;
  assign n4116 = n4149 | n6162;
  assign n4121 = ~preset & (\[17336]  | n3858 | n3859);
  assign n4126 = \[17349]  & ~preset & ~\[17271] ;
  assign n4131 = \[17362]  & ~preset & ~\[17167] ;
  assign n4136 = \[17375]  & ~preset & ~\[17297] ;
  assign n4141 = ~\[17388]  & ~preset & \[16933] ;
  assign n4146 = n6168 | n6169;
  assign n4150 = \[17843]  & ~preset & ~\[17414] ;
  assign n4155 = ~preset & ~\[17700]  & (\[17427]  | \[17518] );
  assign n4160 = n5734 & n5729 & ~preset & n3798;
  assign n4165 = n6175 | n6176;
  assign n4169 = ~preset & (\[17479]  | n3858 | n3859);
  assign n4174 = n4127 | n6177;
  assign n4179 = \[17505]  & ~preset & ~\[17414] ;
  assign n4184 = ~preset & ~\[17700]  & (\[17518]  | \[17817] );
  assign n4189 = n4126_1 | (\[17531]  & n3784);
  assign n4194 = ~preset & (n3877 ? ppeaki_7_7_ : \[17544] );
  assign n4199 = n6183 | n6184;
  assign n4203 = ~preset & ~n3786 & (\[17570]  | n3785);
  assign n4208 = ~preset & ~\[17700]  & (\[17583]  | \[17648] );
  assign n4213 = n4114 | (~n3786 & n6195);
  assign n4218 = ~preset & (n3877 ? ppeaki_6_6_ : \[17609] );
  assign n4223 = n6201 | n6202;
  assign n4227 = ~preset & ~n3786 & (\[17570]  | \[17635] );
  assign n4232 = ~preset & ~\[17700]  & (\[17427]  | \[17648] );
  assign n4237 = n6191 & n6188 & ~preset & n6187;
  assign n4242 = ~preset & (n3877 ? ppeaki_5_5_ : \[17674] );
  assign n4247 = n6208 | n6209;
  assign n4251 = \[18142]  & ~preset & ~\[17700] ;
  assign n4256 = ~preset & (n3877 ? ppeaki_4_4_ : \[17713] );
  assign n4261 = n6215 | n6216;
  assign n4265 = \[17739]  & ~preset & ~\[17700] ;
  assign n4270 = n3784 & (\[17752]  | (n3798 & n5729));
  assign n4275 = n4082 | n6217;
  assign n4280 = n4080 | n6218;
  assign n4285 = ~preset & ~\[17414]  & (\[17791]  | n3788);
  assign n4290 = n3786 & ~preset & ~pdn;
  assign n4295 = n4079 | (~preset & ~\[17700]  & \[17817] );
  assign n4300 = n6229 | n6227 | n6228;
  assign n4304 = ~preset & ~\[17414]  & (\[17843]  | (\[17791]  & ~\[17843] ));
  assign n4309 = ~preset & (\[17856]  | n3790);
  assign n4314 = ~preset & (\[17869]  | n3858 | n3859);
  assign n4319 = ~preset & (\[17882]  | n3858 | n3859);
  assign n4324 = n6254 | n6251 | n6252;
  assign n4328 = ~preset & (\[17908]  | n3858 | n3859);
  assign n4333 = n4077 | n6255;
  assign n4338 = ~preset & (\[17934]  | n3858 | n3859);
  assign n4343 = ~preset & (\[17947]  | n3858 | n3859);
  assign n4348 = ~preset & (\[17960]  | n3858 | n3859);
  assign n4353 = n4075 | n6256;
  assign n4358 = ~preset & ~n3786 & (\[17635]  | \[17986] );
  assign n4363 = ~preset & ~\[17700]  & (\[17999]  | \[18077] );
  assign n4368 = n4073 | n4074;
  assign n4373 = n3779 & (\[18025]  | (n3798 & n3806));
  assign n4378 = ~preset & (\[18038]  | n3858 | n3859);
  assign n4383 = ~preset & ~pdn & (\[17414]  | n3786);
  assign n4387 = n4072 | (~preset & ~pdn & \[18064] );
  assign n4392 = ~preset & ~\[17700]  & (\[17583]  | \[18077] );
  assign n4397 = n4070 | n4071_1;
  assign n4402 = ~\[18168]  & ~preset & \[18103] ;
  assign n4407 = ~preset & (\[18116]  | n3858 | n3859);
  assign n4412 = n4068 | n4069;
  assign n4417 = ~preset & ~\[17700]  & (\[18142]  | \[18220] );
  assign n4422 = n4066_1 | n4067;
  assign n4427 = n5730 & n5729 & ~preset & n3798;
  assign n4432 = ~preset & (\[18181]  | n3858 | n3859);
  assign n4437 = n4064 | n6258;
  assign n4442 = ~preset & ~pdn & (\[18207]  | n3790);
  assign n4447 = ~preset & ~\[17700]  & (\[17999]  | \[18220] );
  assign n4452 = n4062 | n4063;
  assign n4457 = \[18246]  & ~preset & ~\[17453] ;
  assign n4462 = n6264 | n6265;
  assign n4466 = n4050 | n4251 | n4049;
  assign n4470 = n4048 | (n3798 & n3800 & n6266);
  assign n4475 = ~\[18376]  & ~preset & \[18298] ;
  assign n4480 = ~preset & ~\[18389]  & (\[18311]  | \[18506] );
  assign n4485 = n6272 | n6273;
  assign n4489 = n4035 | n6274;
  assign n4494 = ~preset & (\[18350]  | n3858 | n3859);
  assign n4499 = ~preset & ~\[18415]  & (\[18363]  | (\[18285]  & ~\[18363] ));
  assign n4504 = ~\[18376]  & ~preset & \[17284] ;
  assign n4509 = ~\[18389]  & ~preset & \[18311] ;
  assign n4514 = n6280 | n6281;
  assign n4518 = ~\[18415]  & ~preset & \[18363] ;
  assign n4523 = ~\[18493]  & ~preset & \[18428] ;
  assign n4528 = \[18441]  & ~preset & ~\[17232] ;
  assign n4533 = n6287 | n6288;
  assign n4537 = n4013 | n4014;
  assign n4542 = \[18480]  & ~preset & ~\[18415] ;
  assign n4547 = n3821 & n3798 & ~preset & ~\[18493] ;
  assign n4552 = n3778 & (\[18506]  | (n3798 & n3801));
  assign n4557 = n6295 | n6296;
  assign n4561 = n6302 | n6303;
  assign n4565 = ~preset & ((\[18545]  & (pdn | n3874_1)) | (~pdn & n3874_1));
  assign n4570 = n6309 | n6310;
  assign n4574 = ~preset & (\[18571]  | n3858 | n3859);
  assign n4579 = ~preset & (\[18584]  | n3858 | n3859);
  assign n4584 = n3982 | (~preset & ~pdn & \[18597] );
  assign n4589 = n6316 | (\[18610]  & n3784) | n6317;
  assign n4594 = n6323 | n6324;
  assign n4598 = n6332 | n3970 | n6331;
  assign n3696_1 = ~\[17843]  & ~preset & \[17791] ;
  assign n3697 = n3857 & n3815 & n3756 & n3796;
  assign n3698 = n3857 & n3814 & n3756 & n3796;
  assign n3699 = n3857 & (n3702 | (n3756 & n3828));
  assign n3700 = n3857 & n3843 & n3756 & n3796;
  assign n3701_1 = n3962_1 & n3756 & n3857;
  assign n3702 = n3804 & (n5628 | (~n3955 & n3963));
  assign n3703 = ~\[18246]  & ~preset & \[17453] ;
  assign n3704 = ~preset & (~n3798 | ~n5729 | ~n5730);
  assign n3705 = ~\[17154]  & ~preset & \[17102] ;
  assign n3706_1 = n3800 & n3798 & ~preset & ~\[18285] ;
  assign n3707 = ~preset & (\[18285]  | ~n3798 | ~n3800);
  assign n3708 = ~\[17362]  & ~preset & \[17167] ;
  assign n3709 = n3801 & n3798 & ~preset & ~\[18506] ;
  assign n3710 = ~preset & (\[18506]  | ~n3798 | ~n3801);
  assign n3711_1 = \[17388]  & ~preset & ~\[17310] ;
  assign n3712 = ((~n3891 ^ n3945) & (~n3893_1 | (n3893_1 & n3894))) | (n3893_1 & ~n3894 & (n3891 ^ n3945));
  assign n3713 = ~preset & (~n3798 | ~n5729 | ~n5734);
  assign n3714 = ((n5483 | n5484) & (~n3880 ^ n3902)) | (~n5483 & ~n5484 & (~n3880 ^ ~n3902));
  assign n3715 = \[18168]  & ~preset & ~\[18103] ;
  assign n3716_1 = ~\[18363]  & ~preset & \[18285] ;
  assign n3717 = ~preset & (\[17284]  | ~n3798 | ~n3802_1);
  assign n3718 = n3802_1 & n3798 & ~preset & ~\[17284] ;
  assign n3719 = n3916 ? ((n3914 & n3915) | (n3892 & (n3914 ^ n3915))) : (n3892 ? (~n3914 & ~n3915) : (~n3914 | (n3914 & ~n3915)));
  assign n3720 = ((n5485 | n5486) & (~n3896 ^ n3917)) | (~n5485 & ~n5486 & (~n3896 ^ ~n3917));
  assign n3721_1 = \[18506]  & ~preset & ~\[18311] ;
  assign n3722 = ~preset & (\[16933]  | ~n3798 | ~n3803);
  assign n3723 = n3803 & n3798 & ~preset & ~\[16933] ;
  assign n3724 = (ppeaka_6_6_ & n3810 & (n3861 ^ ~n3924)) | ((~ppeaka_6_6_ | ~n3810) & (~n3861 ^ ~n3924));
  assign n3725 = ~preset & n3825;
  assign n3726_1 = (ppeaka_10_10_ & n3810 & (n3866 ^ ~n3926)) | ((~ppeaka_10_10_ | ~n3810) & (~n3866 ^ ~n3926));
  assign n3727 = ~\[17986]  & ~preset & \[17635] ;
  assign n3728 = (ppeaka_4_4_ & n3810 & (n3872 ^ ~n3929)) | ((~ppeaka_4_4_ | ~n3810) & (~n3872 ^ ~n3929));
  assign n3729 = ~preset & (\[18025]  | ~n3798 | ~n3806);
  assign n3730 = n3806 & n3798 & ~preset & ~\[18025] ;
  assign n3731_1 = (ppeaka_9_9_ & n3810 & (n3864_1 ^ ~n3932)) | ((~ppeaka_9_9_ | ~n3810) & (~n3864_1 ^ ~n3932));
  assign n3732 = \[18025]  & ~preset & ~\[17037] ;
  assign n3733 = (ppeaka_3_3_ & n3810 & (n3850 ^ ~n3933_1)) | ((~ppeaka_3_3_ | ~n3810) & (~n3850 ^ ~n3933_1));
  assign n3734 = ~preset & (\[17206]  | ~n3798 | ~n3808);
  assign n3735 = n3808 & n3798 & ~preset & ~\[17206] ;
  assign n3736_1 = ((n3870 ^ n3934) & (n3780 | ~n3944)) | (~n3780 & n3944 & (~n3870 ^ n3934));
  assign n3737 = (ppeaka_12_12_ & n3810 & (n3860_1 ^ ~n3935)) | ((~ppeaka_12_12_ | ~n3810) & (~n3860_1 ^ ~n3935));
  assign n3738 = ~preset & (\[17245]  | ~n3798 | ~n3811);
  assign n3739 = n3811 & n3798 & ~preset & ~\[17245] ;
  assign n3740 = n3937 ? ((n3903_1 & n3920) | (n3885 & (n3903_1 | n3920))) : ((~n3903_1 & ~n3920) | (~n3885 & (~n3903_1 | ~n3920)));
  assign n3741_1 = ((n5487 | n5488) & (~n3898_1 ^ n3938_1)) | (~n5487 & ~n5488 & (~n3898_1 ^ ~n3938_1));
  assign n3742 = (ppeaka_7_7_ & n3810 & (n3873 ^ ~n3925)) | ((~ppeaka_7_7_ | ~n3810) & (~n3873 ^ ~n3925));
  assign n3743 = (ppeaka_11_11_ & n3810 & (n3869_1 ^ ~n3927)) | ((~ppeaka_11_11_ | ~n3810) & (~n3869_1 ^ ~n3927));
  assign n3744 = (ppeaka_8_8_ & n3810 & (n3865 ^ ~n3939)) | ((~ppeaka_8_8_ | ~n3810) & (~n3865 ^ ~n3939));
  assign n3745 = (ppeaka_13_13_ & n3810 & (n3863 ^ ~n3936)) | ((~ppeaka_13_13_ | ~n3810) & (~n3863 ^ ~n3936));
  assign n3746_1 = (ppeaka_5_5_ & n3810 & (n3871 ^ ~n3928_1)) | ((~ppeaka_5_5_ | ~n3810) & (~n3871 ^ ~n3928_1));
  assign n3747 = ((n5493 | n5761) & (~n3884 ^ n3919)) | (~n5493 & ~n5761 & (~n3884 ^ ~n3919));
  assign n3748 = \[18077]  & ~preset & ~\[17999] ;
  assign n3749 = (~n5814 & ((~n3848 & n5811) | (~ppeaks_0_0_ & (n3848 | n5811)))) | (~n3848 & ~n5811 & n5814);
  assign n3750_1 = n3827_1 & n3798 & ~preset & ~\[17180] ;
  assign n3751 = ~preset & (\[17180]  | ~n3798 | ~n3827_1);
  assign n3752 = (ppeaka_14_14_ & n3810 & (n3867 ^ ~n3940)) | ((~ppeaka_14_14_ | ~n3810) & (~n3867 ^ ~n3940));
  assign n3753 = (ppeaka_2_2_ & n3810 & (n3849 ^ ~n3943_1)) | ((~ppeaka_2_2_ | ~n3810) & (~n3849 ^ ~n3943_1));
  assign n3754_1 = ~\[17505]  & ~preset & \[17414] ;
  assign n3755 = (ppeaki_10_10_ & n3883_1) | (ppeaki_14_14_ & n3796);
  assign n3756 = ~preset & (\[18636]  | (~n3798 & n5672));
  assign n3757 = \[18220]  & ~preset & ~\[18142] ;
  assign n3758_1 = (ppeaki_12_12_ & n3796) | (ppeaki_8_8_ & n3883_1);
  assign n3759 = (ppeaki_13_13_ & n3796) | (ppeaki_9_9_ & n3883_1);
  assign n3760 = ~\[17635]  & ~preset & \[17570] ;
  assign n3761 = ppeaki_13_13_ & n3883_1;
  assign n3762 = ppeaki_12_12_ & n3883_1;
  assign n3763_1 = ~preset & (\[17115]  | ~n3798 | ~n3826);
  assign n3764 = n3826 & n3798 & ~preset & ~\[17115] ;
  assign n3765 = (ppeaki_11_11_ & n3883_1) | (ppeaki_15_15_ & n3796);
  assign n3766 = (ppeaki_10_10_ & n3796) | (ppeaki_6_6_ & n3883_1);
  assign n3767 = ~\[17648]  & ~preset & \[17427] ;
  assign n3768_1 = (ppeaki_7_7_ & n3883_1) | (ppeaki_11_11_ & n3796);
  assign n3769 = ppeaki_15_15_ & n3883_1;
  assign n3770 = (ppeaki_8_8_ & n3796) | (ppeaki_4_4_ & n3883_1);
  assign n3771 = ppeaki_14_14_ & n3883_1;
  assign n3772_1 = (ppeaki_9_9_ & n3796) | (ppeaki_5_5_ & n3883_1);
  assign n3773 = ~preset & n3824 & (n6130 | n6131);
  assign n3774 = ~preset & n3813 & (n6130 | n6131);
  assign n3775 = ~preset & n3818 & (n6130 | n6131);
  assign n3776 = ~preset & n3807_1 & (n6130 | n6131);
  assign n3777_1 = ~preset & n3820 & (n6130 | n6131);
  assign n3778 = ~preset & ~\[18389] ;
  assign n3779 = ~preset & ~\[17102] ;
  assign n3780 = \[17180]  & ~\[17232] ;
  assign n3781 = \[17206]  & ~\[17271] ;
  assign n3782_1 = ~preset & ~\[17700] ;
  assign n3783 = \[18636]  | (~n3798 & n5672);
  assign n3784 = ~preset & ~\[18636]  & (n3798 | ~n5672);
  assign n3785 = \[18467]  | (n3795 & ~n3804);
  assign n3786 = n6193 | (n6190 & n6191 & n6192);
  assign n3787_1 = n3798 & ~n3797_1 & ~\[18610]  & n3796;
  assign n3788 = ~pdn & (\[17024]  ? \[18545]  : preset_0_0_);
  assign n3789 = (~\[17518]  & \[17817] ) | (~\[17037]  & \[18025] );
  assign n3790 = ~n5631 & (~n5677 | ~n5678) & n5679;
  assign n3791 = n4160 | n4427 | n6133 | n6134;
  assign n3792_1 = n5729 & n3814 & ~\[18168]  & n3798;
  assign n3793 = \[17999]  & ~\[18220] ;
  assign n3794 = \[18363]  & ~\[18415] ;
  assign n3795 = ~pdn & ((\[17024]  & ~\[18545] ) | (~preset_0_0_ & (~\[17024]  | ~\[18545] )));
  assign n3796 = ~n3881 & n3875 & ~n3829 & ~n3862;
  assign n3797_1 = n5659 | n5660 | n5661 | n5662;
  assign n3798 = n5671 | (~n3797_1 & (n5664 | n5668));
  assign n3799 = pdn & ~\[17089] ;
  assign n3800 = ~n3881 & ~n3875 & n3829 & ~n3862;
  assign n3801 = ~n3881 & n3875 & n3829 & n3862;
  assign n3802_1 = n3881 & n3875 & n3829 & ~n3862;
  assign n3803 = n3881 & ~n3875 & n3829 & n3862;
  assign n3804 = \[18064]  ? \[18129]  : pirq_0_0_;
  assign n3805 = \[17635]  & ~\[17986] ;
  assign n3806 = ~n3875 & ~n3829 & ~n3862 & n3881;
  assign n3807_1 = ~\[17037]  & \[18025] ;
  assign n3808 = n3881 & n3875 & ~n3829 & ~n3862;
  assign n3809 = n3808 & ~\[17206]  & n3798;
  assign n3810 = n3803 & ~\[16933]  & n3798;
  assign n3811 = n3881 & n3875 & n3829 & n3862;
  assign n3812_1 = n3881 & ~n3875 & ~n3829 & n3862;
  assign n3813 = n3801 & ~\[18506]  & n3798;
  assign n3814 = (n5680 & n5681) | (n3852_1 & n5682);
  assign n3815 = (n5683 & n5684) | (n3852_1 & n5685);
  assign n3816 = ~\[17570]  & (\[18467]  | (n3795 & ~n3804));
  assign n3817_1 = n3800 & ~\[18285]  & n3798;
  assign n3818 = ~\[17583]  & \[17648] ;
  assign n3819 = n3881 & ~n3875 & n3829 & ~n3862;
  assign n3820 = n3802_1 & ~\[17284]  & n3798;
  assign n3821 = ~n3881 & ~n3875 & ~n3829 & n3862;
  assign n3822_1 = n3826 & ~\[17115]  & n3798;
  assign n3823 = n3827_1 & ~\[17180]  & n3798;
  assign n3824 = ~\[17518]  & \[17817] ;
  assign n3825 = n3804 & n3795 & ~\[17817]  & ~\[18467] ;
  assign n3826 = ~n3881 & n3875 & n3829 & ~n3862;
  assign n3827_1 = n3881 & n3875 & ~n3829 & n3862;
  assign n3828 = ~n3881 & ~n3875 & n3829 & n3862;
  assign n3829 = \[17531]  ? \[18012]  : ppeaki_2_2_;
  assign n3830 = (n3845 & n5633) | (n3844 & n5634);
  assign n3831 = (n3845 & n3847_1) | (n5635 & n5636);
  assign n3832_1 = (n3852_1 & n5637) | (n3851 & n5638);
  assign n3833 = (n3853 & n5640) | (n3847_1 & n5639);
  assign n3834 = (n3846 & n5641) | (n3845 & n3854);
  assign n3835 = (n3855 & n5642) | (n3851 & n5643);
  assign n3836 = (n3853 & n5645) | (n3847_1 & n5644);
  assign n3837_1 = (n3847_1 & n3855) | (n5646 & n5647);
  assign n3838 = (n3854 & n5648) | (n3853 & n5649);
  assign n3839 = (n3852_1 & n5650) | (n3851 & n5651);
  assign n3840 = (n3854 & n5652) | (n3853 & n5653);
  assign n3841 = (n3851 & n5655) | (n3845 & n5654);
  assign n3842_1 = (n3854 & n3855) | (n3846 & n5656);
  assign n3843 = (n3855 & n5657) | (n3844 & n5658);
  assign n3844 = ~\[17609]  & \[17674] ;
  assign n3845 = ppeaki_4_4_ & ppeaki_5_5_;
  assign n3846 = \[17544]  & \[17752] ;
  assign n3847_1 = ~\[17752]  & ppeaki_6_6_ & ppeaki_7_7_;
  assign n3848 = n3809 | n3822_1 | n3823 | n5791;
  assign n3849 = n5806 | (ppeaks_2_2_ & n3848);
  assign n3850 = n5803 | (ppeaks_3_3_ & n3848);
  assign n3851 = \[17752]  & ~\[17544]  & \[17609] ;
  assign n3852_1 = ~\[17752]  & ~ppeaki_5_5_ & ~ppeaki_7_7_;
  assign n3853 = \[17752]  & \[17544]  & ~\[17674] ;
  assign n3854 = ~\[17752]  & ~ppeaki_6_6_ & ppeaki_7_7_;
  assign n3855 = ~ppeaki_4_4_ & ppeaki_5_5_;
  assign n3856_1 = (pdn & ~\[17089] ) | (~\[17596]  & n3790);
  assign n3857 = n3856_1 | \[18636]  | (~n3798 & n5672);
  assign n3858 = n3818 | (~\[17284]  & n3798 & n3802_1);
  assign n3859 = n3789 | n3809 | n3822_1 | n3823;
  assign n3860_1 = n5851 | (ppeaks_12_12_ & n3848);
  assign n3861 = n5794 | (ppeaks_6_6_ & n3848);
  assign n3862 = \[17531]  ? \[18090]  : ppeaki_3_3_;
  assign n3863 = n5848 | (ppeaks_13_13_ & n3848);
  assign n3864_1 = n5829 | (ppeaks_9_9_ & n3848);
  assign n3865 = n5832 | (ppeaks_8_8_ & n3848);
  assign n3866 = n5826 | (ppeaks_10_10_ & n3848);
  assign n3867 = n5845 | (ppeaks_14_14_ & n3848);
  assign n3868 = n5842 | (ppeaks_15_15_ & n3848);
  assign n3869_1 = n5854 | (ppeaks_11_11_ & n3848);
  assign n3870 = n5817 | (ppeaks_1_1_ & n3848);
  assign n3871 = n5797 | (ppeaks_5_5_ & n3848);
  assign n3872 = n5800 | (ppeaks_4_4_ & n3848);
  assign n3873 = n5835 | (ppeaks_7_7_ & n3848);
  assign n3874_1 = \[17024]  ? \[18545]  : preset_0_0_;
  assign n3875 = \[17531]  ? \[18155]  : ppeaki_0_0_;
  assign n3876 = ~n3881 & n3875 & ~n3829 & n3862;
  assign n3877 = n5728 & n3798 & ~\[17752]  & ~n3797_1;
  assign n3878_1 = n5736 | n5735 | (~\[18103]  & \[18168] );
  assign n3879 = (\[17037]  & ~\[17102] ) | (\[17284]  & ~\[18376] );
  assign n3880 = n5745 | (ppeaks_12_12_ & (n3878_1 | n5737));
  assign n3881 = \[17531]  ? \[18233]  : ppeaki_1_1_;
  assign n3882 = n5786 | (ppeaks_15_15_ & (n3878_1 | n5737));
  assign n3883_1 = n3829 | (~n3829 & n3862) | (~n3829 & ~n3862 & n3881);
  assign n3884 = n5759 | (ppeaks_3_3_ & (n3878_1 | n5737));
  assign n3885 = n5780 | (ppeaks_13_13_ & (n3878_1 | n5737));
  assign n3886 = n5772 | (ppeaks_8_8_ & (n3878_1 | n5737));
  assign n3887 = n5763 | (ppeaks_4_4_ & (n3878_1 | n5737));
  assign n3888_1 = n5757 | (ppeaks_2_2_ & (n3878_1 | n5737));
  assign n3889 = n5765 | (ppeaks_5_5_ & (n3878_1 | n5737));
  assign n3890 = n5770 | (ppeaks_7_7_ & (n3878_1 | n5737));
  assign n3891 = n5743 | (ppeaks_1_1_ & (n3878_1 | n5737));
  assign n3892 = n5782 | (ppeaks_14_14_ & (n3878_1 | n5737));
  assign n3893_1 = n3810 | n3820 | n3878_1 | n5739;
  assign n3894 = n5741 | (ppeaks_0_0_ & (n3878_1 | n5737));
  assign n3895 = n5778 | (ppeaks_11_11_ & (n3878_1 | n5737));
  assign n3896 = n5774 | (ppeaks_9_9_ & (n3878_1 | n5737));
  assign n3897 = n5776 | (ppeaks_10_10_ & (n3878_1 | n5737));
  assign n3898_1 = n5767 | (ppeaks_6_6_ & (n3878_1 | n5737));
  assign n3899 = n5716 | n5717 | n5718 | n5719;
  assign n3900 = (~n3878_1 & ~n3945 & ~n5737 & ~n5739) | (n3945 & (n3878_1 | n5737 | n5739));
  assign n3901 = (n3893_1 & ((n3894 & n3945) | (n3891 & (n3894 | n3945)))) | (n3891 & ~n3893_1 & ~n3945);
  assign n3902 = n5755 | (~ppeaka_12_12_ & ~n5532 & ~n5533);
  assign n3903_1 = (n3880 & n3902) | ((n3880 | n3902) & (n5483 | n5484));
  assign n3904 = n5535 | n5534 | (~ppeaka_11_11_ & ~n3952);
  assign n3905 = (n3910 & n3911) | (n3897 & (n3910 | n3911));
  assign n3906 = n3895 | n5534 | n5535 | n5536;
  assign n3907 = n5749 | (n3948_1 & ~n5541 & ~n5542);
  assign n3908_1 = (n3912 & n3913_1) | (n3887 & (n3912 | n3913_1));
  assign n3909 = n5749 | n3889 | n5539;
  assign n3910 = ~n3952 ^ (~n5537 & (n3941 | ~n5751));
  assign n3911 = (n3896 & n3917) | ((n3896 | n3917) & (n5485 | n5486));
  assign n3912 = ~n3947 ^ ((n3792_1 | n3900) & ~n5541);
  assign n3913_1 = (n3884 & n3919) | ((n3884 | n3919) & (n5493 | n5761));
  assign n3914 = n5468 | n5784;
  assign n3915 = (n3903_1 & n3920) | (n3885 & (n3903_1 | n3920));
  assign n3916 = (~n3882 & ~n5462 & ~n5463 & ~n5790) | (n3882 & (n5462 | n5463 | n5790));
  assign n3917 = n5519 | n5518 | (~n3792_1 & ~n3949);
  assign n3918_1 = n5544 | n5543 | (~ppeaka_2_2_ & ~n3945);
  assign n3919 = (n3901 & n3918_1) | (n3888_1 & (n3901 | n3918_1));
  assign n3920 = n3950 ^ (n5532 | n5533);
  assign n3921 = ~n3949 ^ ~n3953_1;
  assign n3922 = (n3898_1 & n3938_1) | ((n3898_1 | n3938_1) & (n5487 | n5488));
  assign n3923_1 = (n3890 & n3922) | ((n3890 | n3922) & (~n3949 ^ ~n3953_1));
  assign n3924 = (n3928_1 & n5822) | (n3871 & (n3928_1 | n5822));
  assign n3925 = (n3924 & n5823) | (n3861 & (n3924 | n5823));
  assign n3926 = (n3932 & n5838) | (n3864_1 & (n3932 | n5838));
  assign n3927 = (n3926 & n5839) | (n3866 & (n3926 | n5839));
  assign n3928_1 = (n3929 & n5821) | (n3872 & (n3929 | n5821));
  assign n3929 = (n3933_1 & n5820) | (n3850 & (n3933_1 | n5820));
  assign n3930 = n3868 ? ((~n3940 & ~n5858) | (~n3867 & (~n3940 | ~n5858))) : ((n3940 & n5858) | (n3867 & (n3940 | n5858)));
  assign n3931 = ~ppeaka_15_15_ | \[16933]  | ~n3798 | ~n3803;
  assign n3932 = (n3939 & n5837) | (n3865 & (n3939 | n5837));
  assign n3933_1 = (n3943_1 & n5819) | (n3849 & (n3943_1 | n5819));
  assign n3934 = (~ppeaks_0_0_ & ~n5814) | (~n3848 & (~n5811 | ~n5814));
  assign n3935 = (n3927 & n5855) | (n3869_1 & (n3927 | n5855));
  assign n3936 = (n3935 & n5856) | (n3860_1 & (n3935 | n5856));
  assign n3937 = ~n3892 ^ (n5468 | n5784);
  assign n3938_1 = ~n3949 & (~ppeaka_6_6_ | ~n3792_1 | n5768);
  assign n3939 = (n3925 & n5836) | (n3873 & (n3925 | n5836));
  assign n3940 = (n3936 & n5857) | (n3863 & (n3936 | n5857));
  assign n3941 = (~ppeaka_8_8_ & (~n3949 | (ppeaka_7_7_ & n3792_1))) | (~n3792_1 & ~n3949) | (n3792_1 & n3949 & ~ppeaka_7_7_ & ppeaka_8_8_);
  assign n3942 = n3886 | n3941;
  assign n3943_1 = (n3944 & n5818 & ~n3780 & n3870) | ((n3780 | ~n3944) & (n3870 | (~n3870 & n5818)));
  assign n3944 = ~ppeaka_1_1_ | \[16933]  | ~n3798 | ~n3803;
  assign n3945 = ~ppeaka_1_1_ | ~n3798 | ~n5729 | ~n5730;
  assign n3946 = ~ppeaka_2_2_ | ~n3798 | ~n5729 | ~n5730;
  assign n3947 = ~ppeaka_4_4_ | ~n3798 | ~n5729 | ~n5730;
  assign n3948_1 = ~ppeaka_5_5_ | ~n3798 | ~n5729 | ~n5730;
  assign n3949 = n5538 | (~n5539 & ~n5749 & n5750);
  assign n3950 = ~ppeaka_13_13_ | ~n3798 | ~n5729 | ~n5730;
  assign n3951 = n5537 | (~ppeaka_8_8_ & ~ppeaka_9_9_ & ~n3941);
  assign n3952 = ~ppeaka_10_10_ | ~n3798 | ~n5729 | ~n5730;
  assign n3953_1 = ~ppeaka_7_7_ | ~n3798 | ~n5729 | ~n5730;
  assign n3954 = ~ppeaka_11_11_ | ~n3798 | ~n5729 | ~n5730;
  assign n3955 = n3874_1 | (~n5631 & (~n5677 | ~n5678));
  assign n3956 = n3829 & n3881 & (~n3862 ^ n3875);
  assign n3957_1 = n3875 & (n3829 ? (~n3862 & ~n3881) : (n3862 & n3881));
  assign n3958 = n3881 & (n3829 ? (~n3862 & n3875) : (n3862 & ~n3875));
  assign n3959 = n3829 & (n3862 ? (n3875 ^ ~n3881) : (~n3875 & n3881));
  assign n3960 = n3959 | (n3796 & n3843);
  assign n3961 = ~n3829 & ~n3862 & n3881;
  assign n3962_1 = (~n3829 & n3862 & ~n3875) | (n3875 & (n3829 ? (~n3862 & n3881) : (n3862 & ~n3881)));
  assign n3963 = ~\[17089]  & ~preset & pdn;
  assign n3964 = (n3829 & ~n3875 & (~n3862 ^ n3881)) | (~n3829 & ~n3862 & n3875 & ~n3881);
  assign n3965 = ~preset & n3816 & (n6130 | n6131);
  assign n3966 = (~n3829 & n3881 & (~n3862 | (n3862 & n3875))) | (n3829 & ~n3862 & n3875 & ~n3881);
  assign n3967_1 = (n3829 & ~n3862 & n3881) | (~n3829 & n3862 & ~n3881) | (n3862 & (n3829 ? (n3875 ^ ~n3881) : (~n3875 & n3881)));
  assign n3968 = n5629 | (~preset & (~n3857 | n5630));
  assign n3969 = n3798 & ~preset & \[16920] ;
  assign n3970 = n3798 & (n3981_1 | n6316 | n6317);
  assign n3971 = \[8255]  & n4081 & (n6130 | n6131);
  assign n3972_1 = \[6065]  & n4518 & (n6130 | n6131);
  assign n3973 = \[9410]  & n4509 & (n6130 | n6131);
  assign n3974 = \[10970]  & n4096 & (n6130 | n6131);
  assign n3975 = ppeaks_7_7_ & n3791 & (n6130 | n6131);
  assign n3976_1 = ~n6131 & ~n6130 & ~preset & paddress_7_7_;
  assign n3977 = \[12905]  & n4011 & (n6130 | n6131);
  assign n3978 = n3965 & \[11075]  & n3804;
  assign n3979 = ppeaka_7_7_ & (n4187 | n4188);
  assign n3980 = ppeakp_7_7_ & (n4189_1 | (~n3804 & n3965));
  assign n3981_1 = \[18610]  & n3784;
  assign n3982 = n6311 & n6191 & ~preset & n6190;
  assign n3983 = \[7625]  & n4081 & (n6130 | n6131);
  assign n3984 = \[6740]  & n4518 & (n6130 | n6131);
  assign n3985 = \[7475]  & n4509 & (n6130 | n6131);
  assign n3986_1 = \[11690]  & n4096 & (n6130 | n6131);
  assign n3987 = ppeaks_6_6_ & n3791 & (n6130 | n6131);
  assign n3988 = ~n6131 & ~n6130 & ~preset & paddress_6_6_;
  assign n3989 = \[13865]  & n4011 & (n6130 | n6131);
  assign n3990 = n3965 & \[9950]  & n3804;
  assign n3991_1 = ppeaka_6_6_ & (n4187 | n4188);
  assign n3992 = ppeakp_6_6_ & (n4189_1 | (~n3804 & n3965));
  assign n3993 = \[6995]  & n4081 & (n6130 | n6131);
  assign n3994 = \[4670]  & n4518 & (n6130 | n6131);
  assign n3995 = \[8105]  & n4509 & (n6130 | n6131);
  assign n3996_1 = \[11465]  & n4096 & (n6130 | n6131);
  assign n3997 = ppeaks_5_5_ & n3791 & (n6130 | n6131);
  assign n3998 = ~n6131 & ~n6130 & ~preset & paddress_5_5_;
  assign n3999 = \[13505]  & n4011 & (n6130 | n6131);
  assign n4000 = n3965 & \[10220]  & n3804;
  assign n4001_1 = ppeaka_5_5_ & (n4187 | n4188);
  assign n4002 = ppeakp_5_5_ & (n4189_1 | (~n3804 & n3965));
  assign n4003 = \[12245]  & n4081 & (n6130 | n6131);
  assign n4004 = \[5375]  & n4518 & (n6130 | n6131);
  assign n4005 = \[6170]  & n4509 & (n6130 | n6131);
  assign n4006_1 = \[5615]  & n4096 & (n6130 | n6131);
  assign n4007 = ppeaks_4_4_ & n3791 & (n6130 | n6131);
  assign n4008 = ~n6131 & ~n6130 & ~preset & paddress_4_4_;
  assign n4009 = \[14675]  & n4011 & (n6130 | n6131);
  assign n4010 = n3965 & \[10505]  & n3804;
  assign n4011_1 = ppeaka_4_4_ & (n4187 | n4188);
  assign n4012 = ppeakp_4_4_ & (n4189_1 | (~n3804 & n3965));
  assign n4013 = n6289 & n3804 & ~\[18467]  & n3795;
  assign n4014 = n4001 & (\[18467]  | (n3795 & ~n3804));
  assign n4015 = \[12455]  & n4081 & (n6130 | n6131);
  assign n4016_1 = \[9995]  & n4518 & (n6130 | n6131);
  assign n4017 = \[6845]  & n4509 & (n6130 | n6131);
  assign n4018 = \[4910]  & n4096 & (n6130 | n6131);
  assign n4019 = ppeaks_3_3_ & n3791 & (n6130 | n6131);
  assign n4020 = ~n6131 & ~n6130 & ~preset & paddress_3_3_;
  assign n4021_1 = \[14255]  & n4011 & (n6130 | n6131);
  assign n4022 = n3965 & \[10790]  & n3804;
  assign n4023 = ppeaka_3_3_ & (n4187 | n4188);
  assign n4024 = ppeakp_3_3_ & (n4189_1 | (~n3804 & n3965));
  assign n4025 = \[12680]  & n4081 & (n6130 | n6131);
  assign n4026_1 = \[9725]  & n4518 & (n6130 | n6131);
  assign n4027 = \[4760]  & n4509 & (n6130 | n6131);
  assign n4028 = \[6980]  & n4096 & (n6130 | n6131);
  assign n4029 = ppeaks_2_2_ & n3791 & (n6130 | n6131);
  assign n4030 = ~n6131 & ~n6130 & ~preset & paddress_2_2_;
  assign n4031_1 = \[15425]  & n4011 & (n6130 | n6131);
  assign n4032 = n3965 & \[11060]  & n3804;
  assign n4033 = ppeaka_2_2_ & (n4187 | n4188);
  assign n4034 = ppeakp_2_2_ & (n4189_1 | (~n3804 & n3965));
  assign n4035 = ~n3859 & ~n3858 & ~preset & \[18337] ;
  assign n4036_1 = n3858 & ~preset & ppeaka_0_0_;
  assign n4037 = \[12920]  & n4081 & (n6130 | n6131);
  assign n4038 = \[9290]  & n4518 & (n6130 | n6131);
  assign n4039 = \[10310]  & n4509 & (n6130 | n6131);
  assign n4040 = \[6305]  & n4096 & (n6130 | n6131);
  assign n4041_1 = ppeaks_1_1_ & n3791 & (n6130 | n6131);
  assign n4042 = ~n6131 & ~n6130 & ~preset & paddress_1_1_;
  assign n4043 = \[12005]  & n4011 & (n6130 | n6131);
  assign n4044 = n3965 & \[11315]  & n3804;
  assign n4045 = ppeaka_1_1_ & (n4187 | n4188);
  assign n4046_1 = ppeakp_1_1_ & (n4189_1 | (~n3804 & n3965));
  assign n4047 = ~preset & n3793 & (n6130 | n6131);
  assign n4048 = ~\[18415]  & ~preset & \[18285] ;
  assign n4049 = \[17739]  & ~preset & piack_0_0_;
  assign n4050 = ~\[17700]  & ~preset & piack_0_0_;
  assign n4051_1 = \[13175]  & n4081 & (n6130 | n6131);
  assign n4052 = \[8630]  & n4518 & (n6130 | n6131);
  assign n4053 = \[10025]  & n4509 & (n6130 | n6131);
  assign n4054 = \[8240]  & n4096 & (n6130 | n6131);
  assign n4055 = ppeaks_0_0_ & n3791 & (n6130 | n6131);
  assign n4056_1 = ~n6131 & ~n6130 & ~preset & paddress_0_0_;
  assign n4057 = \[12890]  & n4011 & (n6130 | n6131);
  assign n4058 = n3965 & \[11555]  & n3804;
  assign n4059 = ppeaka_0_0_ & (n4187 | n4188);
  assign n4060 = ppeakp_0_0_ & (n4189_1 | (~n3804 & n3965));
  assign n4061_1 = n4150 & (n6130 | n6131);
  assign n4062 = ~preset & \[18233]  & (\[17531]  | ~n3798);
  assign n4063 = n3798 & ~\[17531]  & ~preset & ppeaki_1_1_;
  assign n4064 = ~n3859 & ~n3858 & ~preset & \[18194] ;
  assign n4065 = n3858 & ~preset & ppeaka_11_11_;
  assign n4066_1 = ~preset & \[18155]  & (\[17531]  | ~n3798);
  assign n4067 = n3798 & ~\[17531]  & ~preset & ppeaki_0_0_;
  assign n4068 = n6257 & (\[18467]  | ~n3795 | (n3795 & ~n3804));
  assign n4069 = n3804 & n3795 & ~preset & ~\[18467] ;
  assign n4070 = ~preset & \[18090]  & (\[17531]  | ~n3798);
  assign n4071_1 = n3798 & ~\[17531]  & ~preset & ppeaki_3_3_;
  assign n4072 = n3804 & n3795 & n4001 & ~\[18467] ;
  assign n4073 = ~preset & \[18012]  & (\[17531]  | ~n3798);
  assign n4074 = n3798 & ~\[17531]  & ~preset & ppeaki_2_2_;
  assign n4075 = ~n3859 & ~n3858 & ~preset & \[17973] ;
  assign n4076_1 = n3858 & ~preset & ppeaka_12_12_;
  assign n4077 = ~n3859 & ~n3858 & ~preset & \[17921] ;
  assign n4078 = n3858 & ~preset & ppeaka_10_10_;
  assign n4079 = n3804 & n3795 & ~\[18467]  & n3782_1;
  assign n4080 = ~n3859 & ~n3858 & ~preset & \[17778] ;
  assign n4081_1 = n3858 & ~preset & ppeaka_14_14_;
  assign n4082 = ~n3859 & ~n3858 & ~preset & \[17765] ;
  assign n4083 = n3858 & ~preset & ppeaka_9_9_;
  assign n4084 = \[10985]  & n4081 & (n6130 | n6131);
  assign n4085 = \[6080]  & n4518 & (n6130 | n6131);
  assign n4086_1 = \[5480]  & n4509 & (n6130 | n6131);
  assign n4087 = \[12650]  & n4096 & (n6130 | n6131);
  assign n4088 = ppeaks_14_14_ & n3791 & (n6130 | n6131);
  assign n4089 = ~n6131 & ~n6130 & ~preset & paddress_14_14_;
  assign n4090 = \[14270]  & n4011 & (n6130 | n6131);
  assign n4091_1 = n3965 & \[12260]  & n3804;
  assign n4092 = ppeaka_14_14_ & (n4187 | n4188);
  assign n4093 = ppeakp_14_14_ & (n4189_1 | (~n3804 & n3965));
  assign n4094 = \[6320]  & n4081 & (n6130 | n6131);
  assign n4095 = \[6755]  & n4518 & (n6130 | n6131);
  assign n4096_1 = \[8765]  & n4509 & (n6130 | n6131);
  assign n4097 = \[12425]  & n4096 & (n6130 | n6131);
  assign n4098 = ppeaks_15_15_ & n3791 & (n6130 | n6131);
  assign n4099 = ~n6131 & ~n6130 & ~preset & paddress_15_15_;
  assign n4100 = \[13880]  & n4011 & (n6130 | n6131);
  assign n4101_1 = n3965 & \[12470]  & n3804;
  assign n4102 = ppeaka_15_15_ & (n4187 | n4188);
  assign n4103 = ppeakp_15_15_ & (n4189_1 | (~n3804 & n3965));
  assign n4104 = \[10415]  & n4081 & (n6130 | n6131);
  assign n4105 = \[10010]  & n4518 & (n6130 | n6131);
  assign n4106_1 = \[6860]  & n4509 & (n6130 | n6131);
  assign n4107 = \[14660]  & n4096 & (n6130 | n6131);
  assign n4108 = ppeaks_12_12_ & n3791 & (n6130 | n6131);
  assign n4109 = ~n6131 & ~n6130 & ~preset & paddress_12_12_;
  assign n4110 = \[15065]  & n4011 & (n6130 | n6131);
  assign n4111_1 = n3965 & \[12050]  & n3804;
  assign n4112 = ppeaka_12_12_ & (n4187 | n4188);
  assign n4113 = ppeakp_12_12_ & (n4189_1 | (~n3804 & n3965));
  assign n4114 = n6194 & (~n6187 | ~n6188 | ~n6191);
  assign n4115 = \[17986]  & (n5631 | (n5677 & n5678));
  assign n4116_1 = \[10700]  & n4081 & (n6130 | n6131);
  assign n4117 = \[9740]  & n4518 & (n6130 | n6131);
  assign n4118 = \[4775]  & n4509 & (n6130 | n6131);
  assign n4119 = \[14240]  & n4096 & (n6130 | n6131);
  assign n4120 = ppeaks_13_13_ & n3791 & (n6130 | n6131);
  assign n4121_1 = ~n6131 & ~n6130 & ~preset & paddress_13_13_;
  assign n4122 = \[14690]  & n4011 & (n6130 | n6131);
  assign n4123 = n3965 & \[12170]  & n3804;
  assign n4124 = ppeaka_13_13_ & (n4187 | n4188);
  assign n4125 = ppeakp_13_13_ & (n4189_1 | (~n3804 & n3965));
  assign n4126_1 = n3798 & ~preset & ~\[18636] ;
  assign n4127 = ~n3859 & ~n3858 & ~preset & \[17492] ;
  assign n4128 = n3858 & ~preset & ppeaka_13_13_;
  assign n4129 = \[9860]  & n4081 & (n6130 | n6131);
  assign n4130 = \[9305]  & n4518 & (n6130 | n6131);
  assign n4131_1 = \[9770]  & n4509 & (n6130 | n6131);
  assign n4132 = \[13850]  & n4096 & (n6130 | n6131);
  assign n4133 = ppeaks_10_10_ & n3791 & (n6130 | n6131);
  assign n4134 = ~n6131 & ~n6130 & ~preset & paddress_10_10_;
  assign n4135 = \[12665]  & n4011 & (n6130 | n6131);
  assign n4136_1 = n3965 & \[11795]  & n3804;
  assign n4137 = ppeaka_10_10_ & (n4187 | n4188);
  assign n4138 = ppeakp_10_10_ & (n4189_1 | (~n3804 & n3965));
  assign n4139 = \[10130]  & n4081 & (n6130 | n6131);
  assign n4140 = \[8645]  & n4518 & (n6130 | n6131);
  assign n4141_1 = \[10595]  & n4509 & (n6130 | n6131);
  assign n4142 = \[13490]  & n4096 & (n6130 | n6131);
  assign n4143 = ppeaks_11_11_ & n3791 & (n6130 | n6131);
  assign n4144 = ~n6131 & ~n6130 & ~preset & paddress_11_11_;
  assign n4145 = \[12125]  & n4011 & (n6130 | n6131);
  assign n4146_1 = n3965 & \[11915]  & n3804;
  assign n4147 = ppeaka_11_11_ & (n4187 | n4188);
  assign n4148 = ppeakp_11_11_ & (n4189_1 | (~n3804 & n3965));
  assign n4149 = ~n3859 & ~n3858 & ~preset & \[17323] ;
  assign n4150_1 = n3858 & ~preset & ppeaka_2_2_;
  assign n4151 = ~n3859 & ~n3858 & ~preset & \[17258] ;
  assign n4152 = n3858 & ~preset & ppeaka_1_1_;
  assign n4153 = ~n3859 & ~n3858 & ~preset & \[17193] ;
  assign n4154 = n3858 & ~preset & ppeaka_4_4_;
  assign n4155_1 = ~n3859 & ~n3858 & ~preset & \[17128] ;
  assign n4156 = n3858 & ~preset & ppeaka_3_3_;
  assign n4157 = ~n3859 & ~n3858 & ~preset & \[17076] ;
  assign n4158 = n3858 & ~preset & ppeaka_15_15_;
  assign n4159 = ~n3859 & ~n3858 & ~preset & \[17063] ;
  assign n4160_1 = n3858 & ~preset & ppeaka_6_6_;
  assign n4161 = ~n3859 & ~n3858 & ~preset & \[16998] ;
  assign n4162 = n3858 & ~preset & ppeaka_5_5_;
  assign n4163 = ~n3859 & ~n3858 & ~preset & \[16959] ;
  assign n4164 = n3858 & ~preset & ppeaka_8_8_;
  assign n4165_1 = \[9590]  & n4081 & (n6130 | n6131);
  assign n4166 = \[7370]  & n4518 & (n6130 | n6131);
  assign n4167 = \[10040]  & n4509 & (n6130 | n6131);
  assign n4168 = \[15770]  & n4096 & (n6130 | n6131);
  assign n4169_1 = ppeaks_9_9_ & n3791 & (n6130 | n6131);
  assign n4170 = ~n6131 & ~n6130 & ~preset & paddress_9_9_;
  assign n4171 = \[12440]  & n4011 & (n6130 | n6131);
  assign n4172 = n3965 & \[11570]  & n3804;
  assign n4173 = ppeaka_9_9_ & (n4187 | n4188);
  assign n4174_1 = ppeakp_9_9_ & (n4189_1 | (~n3804 & n3965));
  assign n4175 = ~n3859 & ~n3858 & ~preset & \[16907] ;
  assign n4176 = n3858 & ~preset & ppeaka_7_7_;
  assign n4177 = \[8915]  & n4081 & (n6130 | n6131);
  assign n4178 = \[8000]  & n4518 & (n6130 | n6131);
  assign n4179_1 = \[8750]  & n4509 & (n6130 | n6131);
  assign n4180 = \[11225]  & n4096 & (n6130 | n6131);
  assign n4181 = ppeaks_8_8_ & n3791 & (n6130 | n6131);
  assign n4182 = ~n6131 & ~n6130 & ~preset & paddress_8_8_;
  assign n4183 = \[13160]  & n4011 & (n6130 | n6131);
  assign n4184_1 = n3965 & \[11330]  & n3804;
  assign n4185 = ppeaka_8_8_ & (n4187 | n4188);
  assign n4186 = ppeakp_8_8_ & (n4189_1 | (~n3804 & n3965));
  assign n4187 = ~preset & n3817_1 & (n6130 | n6131);
  assign n4188 = n4056 & (n6130 | n6131);
  assign n4189_1 = n4031 & (n6130 | n6131);
  assign n4190 = ~preset & \[16085]  & (~n3798 | ~n5732);
  assign n4191 = ~preset & \[16070]  & (~n3798 | ~n5731);
  assign n4192 = ~preset & \[16055]  & (\[18103]  | ~\[18168] );
  assign n4193 = \[16025]  & n3704;
  assign n4194_1 = ~preset & \[16010]  & (~n3798 | ~n5733);
  assign n4195 = n5733 & n3798 & ~preset & pdata_9_9_;
  assign n4196 = ~preset & \[15995]  & (~n3798 | ~n5733);
  assign n4197 = n5733 & n3798 & ~preset & pdata_0_0_;
  assign n4198 = ~preset & \[15980]  & (~n3798 | ~n5732);
  assign n4199_1 = n5732 & n3798 & ~preset & pdata_7_7_;
  assign n4200 = ~preset & \[15965]  & (~n3798 | ~n5731);
  assign n4201 = n5731 & n3798 & ~preset & pdata_14_14_;
  assign n4202 = ~preset & \[15920]  & (~\[17102]  | \[17154] );
  assign n4203_1 = ~preset & \[15905]  & (~\[17102]  | \[17154] );
  assign n4204 = n3857 & n3827_1 & \[9860]  & n3756;
  assign n4205 = n3963 & n3874_1 & \[10205]  & n3857;
  assign n4206 = n3857 & n3826 & \[12665]  & n3756;
  assign n4207 = n3857 & n3808 & \[13850]  & n3756;
  assign n4208_1 = n3857 & n3806 & \[10400]  & n3756;
  assign n4209 = n3857 & n3812_1 & \[6155]  & n3756;
  assign n4210 = n3857 & n3801 & \[8135]  & n3756;
  assign n4211 = n3876 & n3857 & \[14585]  & n3756;
  assign n4212 = n3857 & n3821 & \[5450]  & n3756;
  assign n4213_1 = n3857 & n3802_1 & \[8060]  & n3756;
  assign n4214 = n3857 & n3803 & \[8810]  & n3756;
  assign n4215 = n3857 & \[12860]  & n3702;
  assign n4216 = n3857 & n3800 & \[4700]  & n3756;
  assign n4217 = ppeaks_10_10_ & (n5708 | n5709);
  assign n4218_1 = n3801 & \[15665]  & n3756;
  assign n4219 = \[15860]  & (n3968 | n5701 | n5702);
  assign n4220 = \[13130]  & n3804 & (n5627 | n5628);
  assign n4221 = n3801 & \[9980]  & n3756;
  assign n4222 = \[15845]  & (n3968 | n5701 | n5702);
  assign n4223_1 = \[9500]  & n3804 & (n5627 | n5628);
  assign n4224 = n3843 & n3796 & ppeaka_6_6_ & n3756;
  assign n4225 = n3957_1 & \[8330]  & n3756;
  assign n4226 = n3811 & \[5660]  & n3756;
  assign n4227_1 = n3962_1 & ppeakb_5_5_ & n3756;
  assign n4228 = n3819 & \[6560]  & n3756;
  assign n4229 = n3808 & \[11465]  & n3756;
  assign n4230 = n3800 & \[15590]  & n3756;
  assign n4231 = n3814 & n3796 & \[14105]  & n3756;
  assign n4232_1 = n3803 & \[7670]  & n3756;
  assign n4233 = n3815 & n3796 & ~ppeaka_5_5_ & n3756;
  assign n4234 = n3815 & n3796 & ~ppeakb_5_5_ & n3756;
  assign n4235 = ppeakp_5_5_ & (n3702 | (n3756 & n3828));
  assign n4236 = n3806 & \[14825]  & n3756;
  assign n4237_1 = ppeaka_5_5_ & ((n3756 & n3801) | n3968);
  assign n4238 = n3857 & n3811 & \[8315]  & n3756;
  assign n4239 = n3857 & n3819 & \[14435]  & n3756;
  assign n4240 = n3957_1 & n3857 & \[15140]  & n3756;
  assign n4241 = n3857 & n3808 & \[12650]  & n3756;
  assign n4242_1 = n3857 & n3806 & \[15575]  & n3756;
  assign n4243 = n3857 & n3803 & \[6335]  & n3756;
  assign n4244 = n3857 & n3800 & \[9080]  & n3756;
  assign n4245 = ppeaka_14_14_ & ((n3756 & n3801) | n3968);
  assign n4246 = n3966 & n3857 & ppeaka_7_7_ & n3756;
  assign n4247_1 = n3857 & n3812_1 & \[13340]  & n3756;
  assign n4248 = n3857 & n3801 & \[14930]  & n3756;
  assign n4249 = n3876 & n3857 & \[15980]  & n3756;
  assign n4250 = n3857 & n3821 & \[5915]  & n3756;
  assign n4251_1 = n3857 & n3802_1 & \[14450]  & n3756;
  assign n4252 = n3857 & n3803 & \[5315]  & n3756;
  assign n4253 = n3857 & \[7055]  & n3702;
  assign n4254 = n3857 & n3800 & \[9095]  & n3756;
  assign n4255 = ppeakb_7_7_ & ((n3756 & n3960) | n3968);
  assign n4256_1 = ~preset & \[15785]  & (~\[17791]  | \[17843] );
  assign n4257 = ~preset & \[15725]  & (~n3798 | ~n5731);
  assign n4258 = ~preset & \[15710]  & (\[18103]  | ~\[18168] );
  assign n4259 = n3715 & (n3888_1 ? (n3901 ^ ~n3918_1) : (~n3901 ^ ~n3918_1));
  assign n4260 = n4427 & (n3886 ? (n3923_1 ^ ~n3941) : (~n3923_1 ^ ~n3941));
  assign n4261_1 = ~preset & \[15650]  & (~n3798 | ~n5733);
  assign n4262 = n5733 & n3798 & ~preset & pdata_1_1_;
  assign n4263 = ~preset & \[15635]  & (~n3798 | ~n5732);
  assign n4264 = n5732 & n3798 & ~preset & pdata_6_6_;
  assign n4265_1 = ~preset & \[15620]  & (~n3798 | ~n5731);
  assign n4266 = n5731 & n3798 & ~preset & pdata_15_15_;
  assign n4267 = ~preset & \[15575]  & (~\[17102]  | \[17154] );
  assign n4268 = ~preset & \[15560]  & (~\[17102]  | \[17154] );
  assign n4269 = n3857 & n3827_1 & \[13175]  & n3756;
  assign n4270_1 = n3963 & n3874_1 & \[9935]  & n3857;
  assign n4271 = n3857 & n3826 & \[12890]  & n3756;
  assign n4272 = n3857 & n3808 & \[8240]  & n3756;
  assign n4273 = n3857 & n3806 & \[10670]  & n3756;
  assign n4274 = n3857 & n3812_1 & \[15380]  & n3756;
  assign n4275_1 = n3857 & n3801 & \[7490]  & n3756;
  assign n4276 = n3876 & n3857 & \[13400]  & n3756;
  assign n4277 = n3857 & n3821 & \[6125]  & n3756;
  assign n4278 = n3857 & n3802_1 & \[7415]  & n3756;
  assign n4279 = n3857 & n3803 & \[9455]  & n3756;
  assign n4280_1 = n3857 & \[12605]  & n3702;
  assign n4281 = n3857 & n3800 & \[5390]  & n3756;
  assign n4282 = ppeaks_0_0_ & (n5708 | n5709);
  assign n4283 = n3801 & \[9710]  & n3756;
  assign n4284 = \[15515]  & (n3968 | n5701 | n5702);
  assign n4285_1 = \[13475]  & n3804 & (n5627 | n5628);
  assign n4286 = n3801 & \[15305]  & n3756;
  assign n4287 = \[15500]  & (n3968 | n5701 | n5702);
  assign n4288 = \[9800]  & n3804 & (n5627 | n5628);
  assign n4289 = n3843 & n3796 & ppeaka_5_5_ & n3756;
  assign n4290_1 = n3957_1 & \[14765]  & n3756;
  assign n4291 = n3811 & \[8975]  & n3756;
  assign n4292 = n3962_1 & ppeakb_4_4_ & n3756;
  assign n4293 = n3819 & \[14870]  & n3756;
  assign n4294 = n3808 & \[5615]  & n3756;
  assign n4295_1 = n3800 & \[13280]  & n3756;
  assign n4296 = n3814 & n3796 & \[14525]  & n3756;
  assign n4297 = n3803 & \[8300]  & n3756;
  assign n4298 = n3815 & n3796 & ~ppeaka_4_4_ & n3756;
  assign n4299 = n3815 & n3796 & ~ppeakb_4_4_ & n3756;
  assign n4300_1 = ppeakp_4_4_ & (n3702 | (n3756 & n3828));
  assign n4301 = n3806 & \[15905]  & n3756;
  assign n4302 = ppeaka_4_4_ & ((n3756 & n3801) | n3968);
  assign n4303 = n3957_1 & \[13550]  & n3756;
  assign n4304_1 = n3811 & \[6365]  & n3756;
  assign n4305 = n3962_1 & ppeakb_15_15_ & n3756;
  assign n4306 = n3819 & \[7205]  & n3756;
  assign n4307 = n3808 & \[12425]  & n3756;
  assign n4308 = n3800 & \[15950]  & n3756;
  assign n4309_1 = n3814 & n3796 & \[13730]  & n3756;
  assign n4310 = n3803 & \[7010]  & n3756;
  assign n4311 = n3815 & n3796 & ~ppeaka_15_15_ & n3756;
  assign n4312 = n3815 & n3796 & ~ppeakb_15_15_ & n3756;
  assign n4313 = ppeakp_15_15_ & (n3702 | (n3756 & n3828));
  assign n4314_1 = n3806 & \[15215]  & n3756;
  assign n4315 = ppeaka_15_15_ & ((n3756 & n3801) | n3968);
  assign n4316 = n3966 & ppeaka_6_6_ & n3756;
  assign n4317 = n3821 & \[7865]  & n3756;
  assign n4318 = n3802_1 & \[6575]  & n3756;
  assign n4319_1 = n3876 & \[15635]  & n3756;
  assign n4320 = n3800 & \[7160]  & n3756;
  assign n4321 = n3814 & n3796 & \[4385]  & n3756;
  assign n4322 = n3803 & \[4610]  & n3756;
  assign n4323 = n3815 & n3796 & \[7745]  & n3756;
  assign n4324_1 = n3801 & \[10265]  & n3756;
  assign n4325 = ppeakb_6_6_ & ((n3756 & n3960) | n3968);
  assign n4326 = \[7685]  & n3804 & (n5627 | n5628);
  assign n4327 = ~preset & \[15440]  & (~\[17791]  | \[17843] );
  assign n4328_1 = ~preset & \[15410]  & (~\[17427]  | \[17648] );
  assign n4329 = ~preset & \[15395]  & (~\[17427]  | \[17648] );
  assign n4330 = ~preset & \[15380]  & (~n3798 | ~n5733);
  assign n4331 = ~preset & \[15365]  & (~n3798 | ~n5732);
  assign n4332 = n3962 & (n3886 ? (n3923_1 ^ ~n3941) : (~n3923_1 ^ ~n3941));
  assign n4333_1 = ~preset & \[15350]  & (\[18103]  | ~\[18168] );
  assign n4334 = n4427 & (n3895 ? (n3904 ^ ~n3905) : (~n3904 ^ ~n3905));
  assign n4335 = ~preset & \[15290]  & (~n3798 | ~n5733);
  assign n4336 = n5733 & n3798 & ~preset & pdata_2_2_;
  assign n4337 = ~preset & \[15275]  & (~n3798 | ~n5732);
  assign n4338_1 = n5732 & n3798 & ~preset & pdata_9_9_;
  assign n4339 = ~preset & \[15260]  & (~n3798 | ~n5731);
  assign n4340 = n5731 & n3798 & ~preset & pdata_12_12_;
  assign n4341 = ~preset & \[15245]  & (~\[17167]  | \[17362] );
  assign n4342 = ~preset & \[15215]  & (~\[17102]  | \[17154] );
  assign n4343_1 = ~preset & \[15200]  & (~\[17102]  | \[17154] );
  assign n4344 = ppeaka_15_15_ & (n5577 | n5720);
  assign n4345 = n3963 & \[11285]  & n3874_1;
  assign n4346 = ppeakp_15_15_ & (n5722 | n5723 | n5725);
  assign n4347 = n3801 & ppeakb_15_15_ & n3756;
  assign n4348_1 = n3857 & n3827_1 & \[8915]  & n3756;
  assign n4349 = n3963 & n3874_1 & \[10775]  & n3857;
  assign n4350 = n3857 & n3826 & \[13160]  & n3756;
  assign n4351 = n3857 & n3808 & \[11225]  & n3756;
  assign n4352 = n3857 & n3806 & \[7595]  & n3756;
  assign n4353_1 = n3857 & n3812_1 & \[12590]  & n3756;
  assign n4354 = n3857 & n3801 & \[9440]  & n3756;
  assign n4355 = n3876 & n3857 & \[15365]  & n3756;
  assign n4356 = n3857 & n3821 & \[6815]  & n3756;
  assign n4357 = n3857 & n3802_1 & \[10865]  & n3756;
  assign n4358_1 = n3857 & n3803 & \[7520]  & n3756;
  assign n4359 = n3857 & \[13460]  & n3702;
  assign n4360 = n3857 & n3800 & \[6095]  & n3756;
  assign n4361 = ppeaks_8_8_ & (n5708 | n5709);
  assign n4362 = n3801 & \[5975]  & n3756;
  assign n4363_1 = \[15140]  & (n3968 | n5701 | n5702);
  assign n4364 = \[10070]  & n3804 & (n5627 | n5628);
  assign n4365 = n3843 & n3796 & ppeaka_4_4_ & n3756;
  assign n4366 = n3957_1 & \[15860]  & n3756;
  assign n4367 = n3811 & \[9920]  & n3756;
  assign n4368_1 = n3962_1 & ppeakb_3_3_ & n3756;
  assign n4369 = n3819 & \[15245]  & n3756;
  assign n4370 = n3808 & \[4910]  & n3756;
  assign n4371 = n3800 & \[13625]  & n3756;
  assign n4372 = n3814 & n3796 & \[13355]  & n3756;
  assign n4373_1 = n3803 & \[8960]  & n3756;
  assign n4374 = n3815 & n3796 & ~ppeaka_3_3_ & n3756;
  assign n4375 = n3815 & n3796 & ~ppeakb_3_3_ & n3756;
  assign n4376 = ppeakp_3_3_ & (n3702 | (n3756 & n3828));
  assign n4377 = n3806 & \[15560]  & n3756;
  assign n4378_1 = ppeaka_3_3_ & ((n3756 & n3801) | n3968);
  assign n4379 = n3857 & n3811 & \[11510]  & n3756;
  assign n4380 = n3857 & n3819 & \[7190]  & n3756;
  assign n4381 = n3957_1 & n3857 & \[15845]  & n3756;
  assign n4382 = n3857 & n3808 & \[14660]  & n3756;
  assign n4383_1 = n3857 & n3806 & \[4415]  & n3756;
  assign n4384 = n3857 & n3803 & \[4940]  & n3756;
  assign n4385 = n3857 & n3800 & \[7775]  & n3756;
  assign n4386 = ppeaka_12_12_ & ((n3756 & n3801) | n3968);
  assign n4387_1 = n3966 & ppeaka_9_9_ & n3756;
  assign n4388 = n3821 & \[4520]  & n3756;
  assign n4389 = n3802_1 & \[7850]  & n3756;
  assign n4390 = n3876 & \[15275]  & n3756;
  assign n4391 = n3800 & \[14855]  & n3756;
  assign n4392_1 = n3814 & n3796 & \[15185]  & n3756;
  assign n4393 = n3803 & \[6680]  & n3756;
  assign n4394 = n3815 & n3796 & \[8390]  & n3756;
  assign n4395 = n3801 & \[5990]  & n3756;
  assign n4396 = ppeakb_9_9_ & ((n3756 & n3960) | n3968);
  assign n4397_1 = \[5720]  & n3804 & (n5627 | n5628);
  assign n4398 = ~preset & \[15080]  & (~\[17791]  | \[17843] );
  assign n4399 = ~preset & \[15050]  & (~\[17427]  | \[17648] );
  assign n4400 = ~preset & \[15035]  & (~\[17427]  | \[17648] );
  assign n4401 = ~preset & \[15020]  & (~n3798 | ~n5733);
  assign n4402_1 = ~preset & \[15005]  & (~n3798 | ~n5732);
  assign n4403 = n3962 & (n3890 ? (n3921 ^ ~n3922) : (~n3921 ^ ~n3922));
  assign n4404 = ~preset & \[14990]  & (~n3798 | ~n5731);
  assign n4405 = n4547 & (n3885 ? (n3903_1 ^ ~n3920) : (~n3903_1 ^ ~n3920));
  assign n4406 = ~preset & \[14975]  & (\[18103]  | ~\[18168] );
  assign n4407_1 = n3715 & (n3887 ? (n3912 ^ ~n3913_1) : (~n3912 ^ ~n3913_1));
  assign n4408 = n4427 & (n3897 ? (n3910 ^ ~n3911) : (~n3910 ^ ~n3911));
  assign n4409 = ~preset & \[14915]  & (~n3798 | ~n5733);
  assign n4410 = n5733 & n3798 & ~preset & pdata_3_3_;
  assign n4411 = ~preset & \[14900]  & (~n3798 | ~n5732);
  assign n4412_1 = n5732 & n3798 & ~preset & pdata_8_8_;
  assign n4413 = ~preset & \[14885]  & (~n3798 | ~n5731);
  assign n4414 = n5731 & n3798 & ~preset & pdata_13_13_;
  assign n4415 = ~preset & \[14870]  & (~\[17167]  | \[17362] );
  assign n4416 = ~preset & \[14825]  & (~\[17102]  | \[17154] );
  assign n4417_1 = ppeaka_14_14_ & (n5577 | n5720);
  assign n4418 = n3963 & \[11525]  & n3874_1;
  assign n4419 = ppeakp_14_14_ & (n5722 | n5723 | n5725);
  assign n4420 = n3801 & ppeakb_14_14_ & n3756;
  assign n4421 = n3857 & n3827_1 & \[9590]  & n3756;
  assign n4422_1 = n3963 & n3874_1 & \[11045]  & n3857;
  assign n4423 = n3857 & n3826 & \[12440]  & n3756;
  assign n4424 = n3857 & n3808 & \[15770]  & n3756;
  assign n4425 = n3857 & n3806 & \[10685]  & n3756;
  assign n4426 = n3857 & n3812_1 & \[5465]  & n3756;
  assign n4427_1 = n3857 & n3801 & \[8780]  & n3756;
  assign n4428 = n3876 & n3857 & \[14165]  & n3756;
  assign n4429 = n3857 & n3821 & \[4745]  & n3756;
  assign n4430 = n3857 & n3802_1 & \[11135]  & n3756;
  assign n4431 = n3857 & n3803 & \[9470]  & n3756;
  assign n4432_1 = n3857 & \[13820]  & n3702;
  assign n4433 = n3857 & n3800 & \[5405]  & n3756;
  assign n4434 = ppeaks_9_9_ & (n5708 | n5709);
  assign n4435 = n3801 & \[5270]  & n3756;
  assign n4436 = \[14765]  & (n3968 | n5701 | n5702);
  assign n4437_1 = \[12875]  & n3804 & (n5627 | n5628);
  assign n4438 = n3843 & n3796 & ppeaka_3_3_ & n3756;
  assign n4439 = n3957_1 & \[15515]  & n3756;
  assign n4440 = n3811 & \[11720]  & n3756;
  assign n4441 = n3962_1 & ppeakb_2_2_ & n3756;
  assign n4442_1 = n3819 & \[7805]  & n3756;
  assign n4443 = n3808 & \[6980]  & n3756;
  assign n4444 = n3800 & \[14000]  & n3756;
  assign n4445 = n3814 & n3796 & \[13715]  & n3756;
  assign n4446 = n3803 & \[9635]  & n3756;
  assign n4447_1 = n3815 & n3796 & ~ppeaka_2_2_ & n3756;
  assign n4448 = n3815 & n3796 & ~ppeakb_2_2_ & n3756;
  assign n4449 = ppeakp_2_2_ & (n3702 | (n3756 & n3828));
  assign n4450 = n3806 & \[5105]  & n3756;
  assign n4451 = ppeaka_2_2_ & ((n3756 & n3801) | n3968);
  assign n4452_1 = n3857 & n3811 & \[10190]  & n3756;
  assign n4453 = n3962_1 & n3857 & ppeakb_13_13_ & n3756;
  assign n4454 = n3857 & n3819 & \[14015]  & n3756;
  assign n4455 = n3957_1 & n3857 & \[15500]  & n3756;
  assign n4456 = n3857 & n3808 & \[14240]  & n3756;
  assign n4457_1 = n3857 & n3806 & \[15920]  & n3756;
  assign n4458 = n3857 & n3803 & \[5645]  & n3756;
  assign n4459 = n3857 & n3800 & \[8420]  & n3756;
  assign n4460 = ppeaka_13_13_ & ((n3756 & n3801) | n3968);
  assign n4461 = n3966 & ppeaka_8_8_ & n3756;
  assign n4462_1 = n3821 & \[6605]  & n3756;
  assign n4463 = n3802_1 & \[14030]  & n3756;
  assign n4464 = n3876 & \[14900]  & n3756;
  assign n4465 = n3800 & \[8435]  & n3756;
  assign n4466_1 = n3814 & n3796 & \[5810]  & n3756;
  assign n4467 = n3803 & \[6005]  & n3756;
  assign n4468 = n3815 & n3796 & \[9050]  & n3756;
  assign n4469 = n3801 & \[6665]  & n3756;
  assign n4470_1 = ppeakb_8_8_ & ((n3756 & n3960) | n3968);
  assign n4471 = \[6410]  & n3804 & (n5627 | n5628);
  assign n4472 = ~preset & \[14705]  & (~\[17791]  | \[17843] );
  assign n4473 = ~preset & \[14630]  & (~\[17427]  | \[17648] );
  assign n4474 = ~n3825 & ~preset & \[14615] ;
  assign n4475_1 = ~preset & \[14600]  & (~n3798 | ~n5733);
  assign n4476 = n4106 & (n3888_1 ? (n3901 ^ ~n3918_1) : (~n3901 ^ ~n3918_1));
  assign n4477 = ~preset & \[14585]  & (~n3798 | ~n5732);
  assign n4478 = n3962 & (n3897 ? (n3910 ^ ~n3911) : (~n3910 ^ ~n3911));
  assign n4479 = ~preset & \[14570]  & (~n3798 | ~n5732);
  assign n4480_1 = ~preset & \[14555]  & (\[18103]  | ~\[18168] );
  assign n4481 = n3715 & (n3889 ? (n3907 ^ ~n3908_1) : (~n3907 ^ ~n3908_1));
  assign n4482 = n4427 & (n3885 ? (n3903_1 ^ ~n3920) : (~n3903_1 ^ ~n3920));
  assign n4483 = n4427 & (n3887 ? (n3912 ^ ~n3913_1) : (~n3912 ^ ~n3913_1));
  assign n4484 = ~preset & \[14510]  & (\[17310]  | ~\[17388] );
  assign n4485_1 = ~preset & \[14495]  & (~n3798 | ~n5733);
  assign n4486 = n5733 & n3798 & ~preset & pdata_4_4_;
  assign n4487 = ~preset & \[14480]  & (~n3798 | ~n5732);
  assign n4488 = n5732 & n3798 & ~preset & pdata_11_11_;
  assign n4489_1 = ~preset & \[14465]  & (~n3798 | ~n5732);
  assign n4490 = n5732 & n3798 & ~preset & pdata_2_2_;
  assign n4491 = ~preset & \[14450]  & (~\[17284]  | \[18376] );
  assign n4492 = ~preset & \[14435]  & (~\[17167]  | \[17362] );
  assign n4493 = ~preset & \[14405]  & (~\[17102]  | \[17154] );
  assign n4494_1 = ~preset & \[14375]  & (~\[17453]  | \[18246] );
  assign n4495 = ~preset & \[14360]  & (~\[17453]  | \[18246] );
  assign n4496 = ppeaka_4_4_ & (n5577 | n5720);
  assign n4497 = n3963 & \[15440]  & n3874_1;
  assign n4498 = ppeakp_4_4_ & (n5722 | n5723 | n5725);
  assign n4499_1 = n3801 & ppeakb_4_4_ & n3756;
  assign n4500 = n3843 & n3796 & ppeaka_2_2_ & n3756;
  assign n4501 = n3957_1 & \[5030]  & n3756;
  assign n4502 = n3811 & \[11495]  & n3756;
  assign n4503 = n3962_1 & ppeakb_1_1_ & n3756;
  assign n4504_1 = n3819 & \[7175]  & n3756;
  assign n4505 = n3808 & \[6305]  & n3756;
  assign n4506 = n3800 & \[14420]  & n3756;
  assign n4507 = n3814 & n3796 & \[15680]  & n3756;
  assign n4508 = n3803 & \[4925]  & n3756;
  assign n4509_1 = n3815 & n3796 & ~ppeaka_1_1_ & n3756;
  assign n4510 = n3815 & n3796 & ~ppeakb_1_1_ & n3756;
  assign n4511 = ppeakp_1_1_ & (n3702 | (n3756 & n3828));
  assign n4512 = n3806 & \[4400]  & n3756;
  assign n4513 = ppeaka_1_1_ & ((n3756 & n3801) | n3968);
  assign n4514_1 = n3843 & n3796 & ppeaka_11_11_ & n3756;
  assign n4515 = n3957_1 & \[5015]  & n3756;
  assign n4516 = n3811 & \[11015]  & n3756;
  assign n4517 = n3962_1 & ppeakb_10_10_ & n3756;
  assign n4518_1 = n3819 & \[8465]  & n3756;
  assign n4519 = n3808 & \[13850]  & n3756;
  assign n4520 = n3800 & \[6515]  & n3756;
  assign n4521 = n3814 & n3796 & \[14960]  & n3756;
  assign n4522 = n3803 & \[11705]  & n3756;
  assign n4523_1 = n3815 & n3796 & ~ppeaka_10_10_ & n3756;
  assign n4524 = n3815 & n3796 & ~ppeakb_10_10_ & n3756;
  assign n4525 = ppeakp_10_10_ & (n3702 | (n3756 & n3828));
  assign n4526 = n3806 & \[13610]  & n3756;
  assign n4527 = ppeaka_10_10_ & ((n3756 & n3801) | n3968);
  assign n4528_1 = n3966 & ppeaka_3_3_ & n3756;
  assign n4529 = n3821 & \[8510]  & n3756;
  assign n4530 = n3802_1 & \[4490]  & n3756;
  assign n4531 = n3876 & \[14045]  & n3756;
  assign n4532 = n3800 & \[6530]  & n3756;
  assign n4533_1 = n3814 & n3796 & \[7760]  & n3756;
  assign n4534 = n3803 & \[7940]  & n3756;
  assign n4535 = n3815 & n3796 & \[13220]  & n3756;
  assign n4536 = n3801 & \[9215]  & n3756;
  assign n4537_1 = ppeakb_3_3_ & ((n3756 & n3960) | n3968);
  assign n4538 = \[15860]  & n3804 & (n5627 | n5628);
  assign n4539 = ~preset & \[14285]  & (~\[17791]  | \[17843] );
  assign n4540 = ~preset & \[14225]  & (\[17999]  | ~\[18077] );
  assign n4541 = ~preset & \[14210]  & (~\[17427]  | \[17648] );
  assign n4542_1 = ~preset & \[14180]  & (~n3798 | ~n5733);
  assign n4543 = ~preset & \[14165]  & (~n3798 | ~n5732);
  assign n4544 = ~preset & \[14150]  & (~n3798 | ~n5732);
  assign n4545 = n3962 & (n3888_1 ? (n3901 ^ ~n3918_1) : (~n3901 ^ ~n3918_1));
  assign n4546 = ~preset & \[14135]  & (\[18103]  | ~\[18168] );
  assign n4547_1 = n4427 & (n3889 ? (n3907 ^ ~n3908_1) : (~n3907 ^ ~n3908_1));
  assign n4548 = ~preset & \[14090]  & (\[17310]  | ~\[17388] );
  assign n4549 = ~preset & \[14075]  & (~n3798 | ~n5733);
  assign n4550 = n5733 & n3798 & ~preset & pdata_5_5_;
  assign n4551 = ~preset & \[14060]  & (~n3798 | ~n5732);
  assign n4552_1 = n5732 & n3798 & ~preset & pdata_10_10_;
  assign n4553 = ~preset & \[14045]  & (~n3798 | ~n5732);
  assign n4554 = n5732 & n3798 & ~preset & pdata_3_3_;
  assign n4555 = ~preset & \[14030]  & (~\[17284]  | \[18376] );
  assign n4556 = ~preset & \[14015]  & (~\[17167]  | \[17362] );
  assign n4557_1 = ~preset & \[13985]  & (~\[17102]  | \[17154] );
  assign n4558 = ~preset & \[13970]  & (~\[17102]  | \[17154] );
  assign n4559 = ~preset & \[13955]  & (~\[17453]  | \[18246] );
  assign n4560 = ppeaka_5_5_ & (n5577 | n5720);
  assign n4561_1 = n3963 & \[15080]  & n3874_1;
  assign n4562 = ppeakp_5_5_ & (n5722 | n5723 | n5725);
  assign n4563 = n3801 & ppeakb_5_5_ & n3756;
  assign n4564 = n3843 & n3796 & ppeaka_1_1_ & n3756;
  assign n4565_1 = n3957_1 & \[4310]  & n3756;
  assign n4566 = n3811 & \[11255]  & n3756;
  assign n4567 = n3962_1 & ppeakb_0_0_ & n3756;
  assign n4568 = n3819 & \[9110]  & n3756;
  assign n4569 = n3808 & \[8240]  & n3756;
  assign n4570_1 = n3800 & \[14840]  & n3756;
  assign n4571 = n3814 & n3796 & \[16025]  & n3756;
  assign n4572 = n3803 & \[11480]  & n3756;
  assign n4573 = n3815 & n3796 & ~ppeaka_0_0_ & n3756;
  assign n4574_1 = n3815 & n3796 & ~ppeakb_0_0_ & n3756;
  assign n4575 = ppeakp_0_0_ & (n3702 | (n3756 & n3828));
  assign n4576 = n3806 & \[13970]  & n3756;
  assign n4577 = ppeaka_0_0_ & ((n3756 & n3801) | n3968);
  assign n4578 = n3857 & n3811 & \[11735]  & n3756;
  assign n4579_1 = n3962_1 & n3857 & ppeakb_11_11_ & n3756;
  assign n4580 = n3857 & n3819 & \[7820]  & n3756;
  assign n4581 = n3957_1 & n3857 & \[4295]  & n3756;
  assign n4582 = n3857 & n3808 & \[13490]  & n3756;
  assign n4583 = n3857 & n3806 & \[5120]  & n3756;
  assign n4584_1 = n3857 & n3803 & \[9650]  & n3756;
  assign n4585 = n3857 & n3800 & \[7145]  & n3756;
  assign n4586 = ppeaka_11_11_ & ((n3756 & n3801) | n3968);
  assign n4587 = ~preset & \[13895]  & (~\[17791]  | \[17843] );
  assign n4588 = \[13880]  & n3763_1;
  assign n4589_1 = ~preset & \[13835]  & (\[17999]  | ~\[18077] );
  assign n4590 = ~preset & \[13820]  & (~\[17427]  | \[17648] );
  assign n4591 = ~preset & \[13790]  & (~n3798 | ~n5733);
  assign n4592 = n4106 & (n3887 ? (n3912 ^ ~n3913_1) : (~n3912 ^ ~n3913_1));
  assign n4593 = ~preset & \[13775]  & (~n3798 | ~n5732);
  assign n4594_1 = ~preset & \[13745]  & (\[18103]  | ~\[18168] );
  assign n4595 = n3715 & (n3890 ? (n3921 ^ ~n3922) : (~n3921 ^ ~n3922));
  assign n4596 = n4427 & (n3888_1 ? (n3901 ^ ~n3918_1) : (~n3901 ^ ~n3918_1));
  assign n4597 = n4160 & (n3889 ? (n3907 ^ ~n3908_1) : (~n3907 ^ ~n3908_1));
  assign n4598_1 = ~preset & \[13685]  & (~n3798 | ~n5733);
  assign n4599 = n5733 & n3798 & ~preset & pdata_6_6_;
  assign n4600 = ~preset & \[13670]  & (~n3798 | ~n5732);
  assign n4601 = n5732 & n3798 & ~preset & pdata_13_13_;
  assign n4602 = ~preset & \[13655]  & (~n3798 | ~n5732);
  assign n4603 = n5732 & n3798 & ~preset & pdata_0_0_;
  assign n4604 = ~preset & \[13640]  & (~n3798 | ~n5731);
  assign n4605 = n5731 & n3798 & ~preset & pdata_2_2_;
  assign n4606 = ~preset & \[13610]  & (~\[17102]  | \[17154] );
  assign n4607 = ~preset & \[13580]  & (~\[17453]  | \[18246] );
  assign n4608 = ppeaka_6_6_ & (n5577 | n5720);
  assign n4609 = n3963 & \[14705]  & n3874_1;
  assign n4610 = ppeakp_6_6_ & (n5722 | n5723 | n5725);
  assign n4611 = n3801 & ppeakb_6_6_ & n3756;
  assign n4612 = n3801 & \[6650]  & n3756;
  assign n4613 = \[13550]  & (n3968 | n5701 | n5702);
  assign n4614 = \[10355]  & n3804 & (n5627 | n5628);
  assign n4615 = n3966 & n3857 & ppeaka_5_5_ & n3756;
  assign n4616 = n3857 & n3812_1 & \[14075]  & n3756;
  assign n4617 = n3857 & n3801 & \[7910]  & n3756;
  assign n4618 = n3876 & n3857 & \[5240]  & n3756;
  assign n4619 = n3857 & n3821 & \[7235]  & n3756;
  assign n4620 = n3857 & n3802_1 & \[5885]  & n3756;
  assign n4621 = n3857 & n3803 & \[9245]  & n3756;
  assign n4622 = n3857 & \[8330]  & n3702;
  assign n4623 = n3857 & n3800 & \[7790]  & n3756;
  assign n4624 = ppeakb_5_5_ & ((n3756 & n3960) | n3968);
  assign n4625 = ~preset & \[13475]  & (\[17999]  | ~\[18077] );
  assign n4626 = ~preset & \[13460]  & (~\[17427]  | \[17648] );
  assign n4627 = ~preset & \[13430]  & (~n3798 | ~n5733);
  assign n4628 = n4106 & (n3889 ? (n3907 ^ ~n3908_1) : (~n3907 ^ ~n3908_1));
  assign n4629 = ~preset & \[13415]  & (~n3798 | ~n5732);
  assign n4630 = n3962 & (n3895 ? (n3904 ^ ~n3905) : (~n3904 ^ ~n3905));
  assign n4631 = ~preset & \[13400]  & (~n3798 | ~n5732);
  assign n4632 = ~preset & \[13385]  & (\[18103]  | ~\[18168] );
  assign n4633 = n3715 & (n3886 ? (n3923_1 ^ ~n3941) : (~n3923_1 ^ ~n3941));
  assign n4634 = ~preset & \[13340]  & (~n3798 | ~n5733);
  assign n4635 = n5733 & n3798 & ~preset & pdata_7_7_;
  assign n4636 = ~preset & \[13325]  & (~n3798 | ~n5732);
  assign n4637 = n5732 & n3798 & ~preset & pdata_12_12_;
  assign n4638 = ~preset & \[13310]  & (~n3798 | ~n5732);
  assign n4639 = n5732 & n3798 & ~preset & pdata_1_1_;
  assign n4640 = ~preset & \[13295]  & (~n3798 | ~n5731);
  assign n4641 = n5731 & n3798 & ~preset & pdata_1_1_;
  assign n4642 = ~preset & \[13265]  & (~\[17102]  | \[17154] );
  assign n4643 = ~preset & \[13235]  & (~\[17453]  | \[18246] );
  assign n4644 = ~preset & \[13220]  & (~\[17453]  | \[18246] );
  assign n4645 = n3857 & n3811 & \[11270]  & n3756;
  assign n4646 = n3857 & n3819 & \[9125]  & n3756;
  assign n4647 = n3957_1 & n3857 & \[5720]  & n3756;
  assign n4648 = n3857 & n3808 & \[15770]  & n3756;
  assign n4649 = n3857 & n3806 & \[13265]  & n3756;
  assign n4650 = n3857 & n3803 & \[9905]  & n3756;
  assign n4651 = n3857 & n3800 & \[5825]  & n3756;
  assign n4652 = ppeaka_9_9_ & ((n3756 & n3801) | n3968);
  assign n4653 = n3966 & n3857 & ppeaka_4_4_ & n3756;
  assign n4654 = n3857 & n3812_1 & \[14495]  & n3756;
  assign n4655 = n3857 & n3801 & \[7280]  & n3756;
  assign n4656 = n3876 & n3857 & \[12545]  & n3756;
  assign n4657 = n3857 & n3821 & \[9170]  & n3756;
  assign n4658 = n3857 & n3802_1 & \[5195]  & n3756;
  assign n4659 = n3857 & n3803 & \[8585]  & n3756;
  assign n4660 = n3857 & \[14765]  & n3702;
  assign n4661 = n3857 & n3800 & \[5840]  & n3756;
  assign n4662 = ppeakb_4_4_ & ((n3756 & n3960) | n3968);
  assign n4663 = ~preset & \[13130]  & (\[17999]  | ~\[18077] );
  assign n4664 = ~preset & \[13115]  & (~\[17427]  | \[17648] );
  assign n4665 = ~preset & \[13100]  & (~\[17427]  | \[17648] );
  assign n4666 = ~preset & \[13085]  & (~n3798 | ~n5733);
  assign n4667 = ~preset & \[13070]  & (~n3798 | ~n5732);
  assign n4668 = ~preset & \[13055]  & (~n3798 | ~n5732);
  assign n4669 = n3962 & (n3889 ? (n3907 ^ ~n3908_1) : (~n3907 ^ ~n3908_1));
  assign n4670 = ~preset & \[13040]  & (\[18103]  | ~\[18168] );
  assign n4671 = ~preset & \[13025]  & (\[18103]  | ~\[18168] );
  assign n4672 = ~preset & \[13010]  & (~n3798 | ~n5733);
  assign n4673 = n5733 & n3798 & ~preset & pdata_8_8_;
  assign n4674 = ~preset & ppeaki_1_1_ & (~n3857 | n5630);
  assign n4675 = \[10805]  & (n5628 | (~n3955 & n3963));
  assign n4676 = ~preset & ppeaki_10_10_ & (~n3857 | n5630);
  assign n4677 = \[12935]  & (n5628 | (~n3955 & n3963));
  assign n4678 = ~preset & \[12935]  & (~\[17570]  | \[17635] );
  assign n4679 = ~preset & \[12875]  & (\[17999]  | ~\[18077] );
  assign n4680 = ~preset & \[12860]  & (~\[17427]  | \[17648] );
  assign n4681 = ~preset & \[12845]  & (~\[17427]  | \[17648] );
  assign n4682 = ~preset & \[12830]  & (~n3798 | ~n5733);
  assign n4683 = n4106 & (n3890 ? (n3921 ^ ~n3922) : (~n3921 ^ ~n3922));
  assign n4684 = ~preset & \[12815]  & (~n3798 | ~n5732);
  assign n4685 = n3962 & (n3885 ? (n3903_1 ^ ~n3920) : (~n3903_1 ^ ~n3920));
  assign n4686 = ~preset & \[12800]  & (\[18103]  | ~\[18168] );
  assign n4687 = n3715 & (n3897 ? (n3910 ^ ~n3911) : (~n3910 ^ ~n3911));
  assign n4688 = ~preset & \[12770]  & (~n3798 | ~n5732);
  assign n4689 = n5732 & n3798 & ~preset & pdata_14_14_;
  assign n4690 = ~preset & ppeaki_0_0_ & (~n3857 | n5630);
  assign n4691 = \[12695]  & (n5628 | (~n3955 & n3963));
  assign n4692 = ~preset & ppeaki_11_11_ & (~n3857 | n5630);
  assign n4693 = \[11600]  & (n5628 | (~n3955 & n3963));
  assign n4694 = ~preset & \[12695]  & (~\[17570]  | \[17635] );
  assign n4695 = ~preset & \[12635]  & (\[17999]  | ~\[18077] );
  assign n4696 = ~preset & \[12620]  & (~\[17427]  | \[17648] );
  assign n4697 = ~preset & \[12605]  & (~\[17427]  | \[17648] );
  assign n4698 = ~preset & \[12590]  & (~n3798 | ~n5733);
  assign n4699 = n4106 & (n3886 ? (n3923_1 ^ ~n3941) : (~n3923_1 ^ ~n3941));
  assign n4700 = ~preset & \[12575]  & (~n3798 | ~n5732);
  assign n4701 = ~preset & \[12545]  & (~n3798 | ~n5732);
  assign n4702 = n5732 & n3798 & ~preset & pdata_4_4_;
  assign n4703 = ~preset & ppeaki_3_3_ & (~n3857 | n5630);
  assign n4704 = \[11345]  & (n5628 | (~n3955 & n3963));
  assign n4705 = ~preset & ppeaki_12_12_ & (~n3857 | n5630);
  assign n4706 = ~preset & \[12485]  & (~\[17570]  | \[17635] );
  assign n4707 = ~preset & \[12470]  & (\[18142]  | ~\[18220] );
  assign n4708 = \[12425]  & n3734;
  assign n4709 = ~preset & \[12410]  & (\[17999]  | ~\[18077] );
  assign n4710 = ~preset & \[12395]  & (~\[17427]  | \[17648] );
  assign n4711 = ~preset & \[12380]  & (~\[17427]  | \[17648] );
  assign n4712 = ~preset & \[12365]  & (~n3798 | ~n5732);
  assign n4713 = ~preset & \[12350]  & (~n3798 | ~n5732);
  assign n4714 = n3962 & (n3887 ? (n3912 ^ ~n3913_1) : (~n3912 ^ ~n3913_1));
  assign n4715 = n4427 & (n3890 ? (n3921 ^ ~n3922) : (~n3921 ^ ~n3922));
  assign n4716 = ~preset & ppeaki_2_2_ & (~n3857 | n5630);
  assign n4717 = \[11585]  & (n5628 | (~n3955 & n3963));
  assign n4718 = ~preset & ppeaki_13_13_ & (~n3857 | n5630);
  assign n4719 = ~preset & \[12275]  & (~\[17570]  | \[17635] );
  assign n4720 = ~preset & \[12260]  & (\[18142]  | ~\[18220] );
  assign n4721 = n3966 & ppeaka_13_13_ & n3756;
  assign n4722 = n3821 & \[14885]  & n3756;
  assign n4723 = n3802_1 & \[5210]  & n3756;
  assign n4724 = n3876 & \[13670]  & n3756;
  assign n4725 = n3800 & \[4460]  & n3756;
  assign n4726 = n3814 & n3796 & \[13595]  & n3756;
  assign n4727 = n3803 & \[7325]  & n3756;
  assign n4728 = n3815 & n3796 & \[14375]  & n3756;
  assign n4729 = n3801 & \[8570]  & n3756;
  assign n4730 = ppeakb_13_13_ & ((n3756 & n3960) | n3968);
  assign n4731 = \[15500]  & n3804 & (n5627 | n5628);
  assign n4732 = ~preset & \[12200]  & (~\[17570]  | \[17635] );
  assign n4733 = ~preset & \[12185]  & (~\[17570]  | \[17635] );
  assign n4734 = ~preset & \[12170]  & (\[18142]  | ~\[18220] );
  assign n4735 = ~preset & \[12155]  & (~\[17414]  | \[17505] );
  assign n4736 = ~preset & \[12140]  & (~\[17791]  | \[17843] );
  assign n4737 = ~preset & ppeaki_7_7_ & (~n3857 | n5630);
  assign n4738 = \[12065]  & (n5628 | (~n3955 & n3963));
  assign n4739 = ~preset & \[12080]  & (~\[17570]  | \[17635] );
  assign n4740 = ~preset & \[12065]  & (~\[17570]  | \[17635] );
  assign n4741 = ~preset & \[12050]  & (\[18142]  | ~\[18220] );
  assign n4742 = ~preset & \[12035]  & (~\[17414]  | \[17505] );
  assign n4743 = ~preset & \[12020]  & (~\[17791]  | \[17843] );
  assign n4744 = n3966 & ppeaka_15_15_ & n3756;
  assign n4745 = n3821 & \[15620]  & n3756;
  assign n4746 = n3802_1 & \[6590]  & n3756;
  assign n4747 = n3876 & \[4535]  & n3756;
  assign n4748 = n3800 & \[8450]  & n3756;
  assign n4749 = n3814 & n3796 & \[14390]  & n3756;
  assign n4750 = n3803 & \[8600]  & n3756;
  assign n4751 = n3815 & n3796 & \[13580]  & n3756;
  assign n4752 = n3801 & \[7295]  & n3756;
  assign n4753 = ppeakb_15_15_ & ((n3756 & n3960) | n3968);
  assign n4754 = \[13550]  & n3804 & (n5627 | n5628);
  assign n4755 = ~preset & ppeaki_8_8_ & (~n3857 | n5630);
  assign n4756 = \[12485]  & (n5628 | (~n3955 & n3963));
  assign n4757 = ~preset & \[11930]  & (~\[17570]  | \[17635] );
  assign n4758 = ~preset & \[11915]  & (\[18142]  | ~\[18220] );
  assign n4759 = ~preset & \[11900]  & (~\[17414]  | \[17505] );
  assign n4760 = ~preset & \[11885]  & (~\[17414]  | \[17505] );
  assign n4761 = n3966 & n3857 & ppeaka_14_14_ & n3756;
  assign n4762 = n3857 & n3812_1 & \[7250]  & n3756;
  assign n4763 = n3857 & n3801 & \[7925]  & n3756;
  assign n4764 = n3876 & n3857 & \[12770]  & n3756;
  assign n4765 = n3857 & n3821 & \[15965]  & n3756;
  assign n4766 = n3857 & n3802_1 & \[4505]  & n3756;
  assign n4767 = n3857 & n3803 & \[9260]  & n3756;
  assign n4768 = n3857 & \[15140]  & n3702;
  assign n4769 = n3857 & n3800 & \[5165]  & n3756;
  assign n4770 = ppeakb_14_14_ & ((n3756 & n3960) | n3968);
  assign n4771 = ~preset & ppeaki_9_9_ & (~n3857 | n5630);
  assign n4772 = \[12275]  & (n5628 | (~n3955 & n3963));
  assign n4773 = ~preset & \[11810]  & (~\[17570]  | \[17635] );
  assign n4774 = ~preset & \[11795]  & (\[18142]  | ~\[18220] );
  assign n4775 = ~preset & \[11780]  & (~\[17414]  | \[17505] );
  assign n4776 = ~preset & \[11765]  & (~\[17414]  | \[17505] );
  assign n4777 = ~preset & \[11750]  & (~\[17791]  | \[17843] );
  assign n4778 = ~preset & \[11675]  & (\[17037]  | ~\[18025] );
  assign n4779 = ~preset & \[11660]  & (\[17037]  | ~\[18025] );
  assign n4780 = ~preset & \[11615]  & (~n3798 | ~n5731);
  assign n4781 = ~preset & \[11600]  & (~\[17570]  | \[17635] );
  assign n4782 = ~preset & \[11585]  & (~\[17570]  | \[17635] );
  assign n4783 = ~preset & \[11570]  & (\[18142]  | ~\[18220] );
  assign n4784 = ~preset & \[11555]  & (\[18142]  | ~\[18220] );
  assign n4785 = ~preset & \[11540]  & (~\[17414]  | \[17505] );
  assign n4786 = ~preset & \[11525]  & (~\[17791]  | \[17843] );
  assign n4787 = ~preset & \[11450]  & (\[17037]  | ~\[18025] );
  assign n4788 = ~preset & \[11435]  & (\[17037]  | ~\[18025] );
  assign n4789 = n3723 & (n3890 ? (n3921 ^ ~n3922) : (~n3921 ^ ~n3922));
  assign n4790 = ~preset & \[11390]  & (~n3798 | ~n5731);
  assign n4791 = n4547 & (n3895 ? (n3904 ^ ~n3905) : (~n3904 ^ ~n3905));
  assign n4792 = ~preset & \[11345]  & (~\[17570]  | \[17635] );
  assign n4793 = ~preset & \[11330]  & (\[18142]  | ~\[18220] );
  assign n4794 = ~preset & \[11315]  & (\[18142]  | ~\[18220] );
  assign n4795 = ~preset & \[11300]  & (~\[17414]  | \[17505] );
  assign n4796 = ~preset & \[11285]  & (~\[17791]  | \[17843] );
  assign n4797 = ~preset & \[11240]  & (~\[17180]  | \[17232] );
  assign n4798 = ~preset & \[11210]  & (\[17037]  | ~\[18025] );
  assign n4799 = ~preset & \[11195]  & (\[17037]  | ~\[18025] );
  assign n4800 = ~preset & \[11150]  & (~n3798 | ~n5731);
  assign n4801 = n4160 & (n3887 ? (n3912 ^ ~n3913_1) : (~n3912 ^ ~n3913_1));
  assign n4802 = ~preset & \[11090]  & (~\[17570]  | \[17635] );
  assign n4803 = ~preset & \[11075]  & (\[18142]  | ~\[18220] );
  assign n4804 = ~preset & \[11060]  & (\[18142]  | ~\[18220] );
  assign n4805 = ~preset & \[11045]  & (~\[17414]  | \[17505] );
  assign n4806 = ~preset & \[11030]  & (~\[17791]  | \[17843] );
  assign n4807 = ~preset & \[10955]  & (\[17037]  | ~\[18025] );
  assign n4808 = ~preset & \[10940]  & (\[17037]  | ~\[18025] );
  assign n4809 = n3723 & (n3889 ? (n3907 ^ ~n3908_1) : (~n3907 ^ ~n3908_1));
  assign n4810 = ~preset & \[10880]  & (~n3798 | ~n5731);
  assign n4811 = n4547 & (n3888_1 ? (n3901 ^ ~n3918_1) : (~n3901 ^ ~n3918_1));
  assign n4812 = n3718 & (n3886 ? (n3923_1 ^ ~n3941) : (~n3923_1 ^ ~n3941));
  assign n4813 = ~preset & \[10850]  & (\[17310]  | ~\[17388] );
  assign n4814 = ~preset & \[10820]  & (~\[17570]  | \[17635] );
  assign n4815 = ~preset & \[10805]  & (~\[17570]  | \[17635] );
  assign n4816 = ~preset & \[10790]  & (\[18142]  | ~\[18220] );
  assign n4817 = ~preset & \[10775]  & (~\[17414]  | \[17505] );
  assign n4818 = ~preset & \[10760]  & (~\[17791]  | \[17843] );
  assign n4819 = ~preset & \[10730]  & (~\[17180]  | \[17232] );
  assign n4820 = ~preset & \[10715]  & (~\[17180]  | \[17232] );
  assign n4821 = ~preset & \[10655]  & (~\[17635]  | \[17986] );
  assign n4822 = ~preset & \[10625]  & (\[18311]  | ~\[18506] );
  assign n4823 = ~preset & \[10610]  & (\[18311]  | ~\[18506] );
  assign n4824 = n3709 & (n3895 ? (n3904 ^ ~n3905) : (~n3904 ^ ~n3905));
  assign n4825 = ~preset & \[10580]  & (~\[18285]  | \[18363] );
  assign n4826 = ~preset & \[10565]  & (~\[18285]  | \[18363] );
  assign n4827 = ~preset & \[10550]  & (\[17310]  | ~\[17388] );
  assign n4828 = ~preset & ppeaki_5_5_ & (~n3857 | n5630);
  assign n4829 = \[11810]  & (n5628 | (~n3955 & n3963));
  assign n4830 = ~preset & ppeaki_14_14_ & (~n3857 | n5630);
  assign n4831 = ~preset & \[10505]  & (\[18142]  | ~\[18220] );
  assign n4832 = ~preset & \[10490]  & (~\[17414]  | \[17505] );
  assign n4833 = ~preset & \[10475]  & (~\[17414]  | \[17505] );
  assign n4834 = ~preset & \[10445]  & (~\[17180]  | \[17232] );
  assign n4835 = ~preset & \[10430]  & (~\[17180]  | \[17232] );
  assign n4836 = ~preset & \[10370]  & (~\[17635]  | \[17986] );
  assign n4837 = ~preset & \[10355]  & (\[17999]  | ~\[18077] );
  assign n4838 = n3721_1 & (n3885 ? (n3903_1 ^ ~n3920) : (~n3903_1 ^ ~n3920));
  assign n4839 = ~preset & \[10340]  & (\[18311]  | ~\[18506] );
  assign n4840 = n3721_1 & (n3888_1 ? (n3901 ^ ~n3918_1) : (~n3901 ^ ~n3918_1));
  assign n4841 = ~preset & \[10325]  & (\[18311]  | ~\[18506] );
  assign n4842 = ~preset & \[10280]  & (~\[18285]  | \[18363] );
  assign n4843 = n3716_1 & (n3889 ? (n3907 ^ ~n3908_1) : (~n3907 ^ ~n3908_1));
  assign n4844 = ~preset & ppeaki_4_4_ & (~n3857 | n5630);
  assign n4845 = \[11930]  & (n5628 | (~n3955 & n3963));
  assign n4846 = ~preset & ppeaki_15_15_ & (~n3857 | n5630);
  assign n4847 = ~preset & \[10220]  & (\[18142]  | ~\[18220] );
  assign n4848 = ~preset & \[10205]  & (~\[17414]  | \[17505] );
  assign n4849 = ~preset & \[10145]  & (~\[17180]  | \[17232] );
  assign n4850 = ~preset & \[10085]  & (~\[17635]  | \[17986] );
  assign n4851 = ~preset & \[10070]  & (\[17999]  | ~\[18077] );
  assign n4852 = ~preset & \[10055]  & (\[18311]  | ~\[18506] );
  assign n4853 = \[10025]  & n3710;
  assign n4854 = ~preset & \[9950]  & (\[18142]  | ~\[18220] );
  assign n4855 = ~preset & \[9935]  & (~\[17414]  | \[17505] );
  assign n4856 = ~preset & \[9890]  & (~\[17180]  | \[17232] );
  assign n4857 = ~preset & \[9875]  & (~\[17180]  | \[17232] );
  assign n4858 = ~preset & \[9815]  & (~\[17635]  | \[17986] );
  assign n4859 = ~preset & \[9800]  & (\[17999]  | ~\[18077] );
  assign n4860 = n3721_1 & (n3887 ? (n3912 ^ ~n3913_1) : (~n3912 ^ ~n3913_1));
  assign n4861 = ~preset & \[9785]  & (\[18311]  | ~\[18506] );
  assign n4862 = n3709 & (n3897 ? (n3910 ^ ~n3911) : (~n3910 ^ ~n3911));
  assign n4863 = n3706_1 & (n3885 ? (n3903_1 ^ ~n3920) : (~n3903_1 ^ ~n3920));
  assign n4864 = n3706_1 & (n3888_1 ? (n3901 ^ ~n3918_1) : (~n3901 ^ ~n3918_1));
  assign n4865 = ~preset & ppeaki_6_6_ & (~n3857 | n5630);
  assign n4866 = \[12185]  & (n5628 | (~n3955 & n3963));
  assign n4867 = ~preset & \[9680]  & (~\[17414]  | \[17505] );
  assign n4868 = ~preset & \[9665]  & (~\[17414]  | \[17505] );
  assign n4869 = ~preset & \[9620]  & (~\[17180]  | \[17232] );
  assign n4870 = ~preset & \[9605]  & (~\[17180]  | \[17232] );
  assign n4871 = ~preset & \[9575]  & (\[17037]  | ~\[18025] );
  assign n4872 = ~preset & \[9530]  & (~\[17635]  | \[17986] );
  assign n4873 = ~preset & \[9515]  & (~\[17635]  | \[17986] );
  assign n4874 = ~preset & \[9500]  & (\[17999]  | ~\[18077] );
  assign n4875 = \[9455]  & n3722;
  assign n4876 = n3721_1 & (n3886 ? (n3923_1 ^ ~n3941) : (~n3923_1 ^ ~n3941));
  assign n4877 = ~preset & \[9440]  & (\[18311]  | ~\[18506] );
  assign n4878 = n3709 & (n3890 ? (n3921 ^ ~n3922) : (~n3921 ^ ~n3922));
  assign n4879 = ~preset & \[9395]  & (~n3798 | ~n5733);
  assign n4880 = ~preset & \[9380]  & (~n3798 | ~n5731);
  assign n4881 = n4547 & (n3887 ? (n3912 ^ ~n3913_1) : (~n3912 ^ ~n3913_1));
  assign n4882 = ~preset & \[9335]  & (~\[18285]  | \[18363] );
  assign n4883 = n3716_1 & (n3895 ? (n3904 ^ ~n3905) : (~n3904 ^ ~n3905));
  assign n4884 = ~preset & \[9320]  & (~\[18285]  | \[18363] );
  assign n4885 = n3716_1 & (n3888_1 ? (n3901 ^ ~n3918_1) : (~n3901 ^ ~n3918_1));
  assign n4886 = n3706_1 & (n3897 ? (n3910 ^ ~n3911) : (~n3910 ^ ~n3911));
  assign n4887 = n4160 & (n3890 ? (n3921 ^ ~n3922) : (~n3921 ^ ~n3922));
  assign n4888 = ~preset & \[9260]  & (\[17310]  | ~\[17388] );
  assign n4889 = ~preset & \[9245]  & (\[17310]  | ~\[17388] );
  assign n4890 = ~preset & \[9170]  & (~n3798 | ~n5731);
  assign n4891 = n5731 & n3798 & ~preset & pdata_4_4_;
  assign n4892 = ~preset & \[9155]  & (~\[17284]  | \[18376] );
  assign n4893 = ~preset & \[9140]  & (~\[17284]  | \[18376] );
  assign n4894 = ~preset & \[9125]  & (~\[17167]  | \[17362] );
  assign n4895 = ~preset & \[9110]  & (~\[17167]  | \[17362] );
  assign n4896 = ~preset & \[9050]  & (~\[17453]  | \[18246] );
  assign n4897 = ppeaka_0_0_ & (n5577 | n5720);
  assign n4898 = n3963 & \[5675]  & n3874_1;
  assign n4899 = ppeakp_0_0_ & (n5722 | n5723 | n5725);
  assign n4900 = n3801 & ppeakb_0_0_ & n3756;
  assign n4901 = ppeaka_9_9_ & (n5577 | n5720);
  assign n4902 = n3963 & \[11750]  & n3874_1;
  assign n4903 = ppeakp_9_9_ & (n5722 | n5723 | n5725);
  assign n4904 = n3801 & ppeakb_9_9_ & n3756;
  assign n4905 = n3857 & n3827_1 & \[12680]  & n3756;
  assign n4906 = n3963 & n3874_1 & \[10475]  & n3857;
  assign n4907 = n3857 & n3826 & \[15425]  & n3756;
  assign n4908 = n3857 & n3808 & \[6980]  & n3756;
  assign n4909 = n3857 & n3806 & \[10100]  & n3756;
  assign n4910 = n3857 & n3812_1 & \[14600]  & n3756;
  assign n4911 = n3857 & n3801 & \[10325]  & n3756;
  assign n4912 = n3876 & n3857 & \[14150]  & n3756;
  assign n4913 = n3857 & n3821 & \[10880]  & n3756;
  assign n4914 = n3857 & n3802_1 & \[8690]  & n3756;
  assign n4915 = n3857 & n3803 & \[5510]  & n3756;
  assign n4916 = n3857 & \[13100]  & n3702;
  assign n4917 = n3857 & n3800 & \[9320]  & n3756;
  assign n4918 = ppeaks_2_2_ & (n5708 | n5709);
  assign n4919 = n3857 & n3827_1 & \[10130]  & n3756;
  assign n4920 = n3963 & n3874_1 & \[10490]  & n3857;
  assign n4921 = n3857 & n3826 & \[12125]  & n3756;
  assign n4922 = n3857 & n3808 & \[13490]  & n3756;
  assign n4923 = n3857 & n3806 & \[10115]  & n3756;
  assign n4924 = n3857 & n3812_1 & \[6830]  & n3756;
  assign n4925 = n3857 & n3801 & \[7505]  & n3756;
  assign n4926 = n3876 & n3857 & \[13415]  & n3756;
  assign n4927 = n3857 & n3821 & \[11390]  & n3756;
  assign n4928 = n3857 & n3802_1 & \[7430]  & n3756;
  assign n4929 = n3857 & n3803 & \[5525]  & n3756;
  assign n4930 = n3857 & \[13115]  & n3702;
  assign n4931 = n3857 & n3800 & \[9335]  & n3756;
  assign n4932 = ppeaks_11_11_ & (n5708 | n5709);
  assign n4933 = ~preset & \[8945]  & (~\[17180]  | \[17232] );
  assign n4934 = ~preset & \[8930]  & (~\[17180]  | \[17232] );
  assign n4935 = ~preset & \[8900]  & (\[17037]  | ~\[18025] );
  assign n4936 = ~preset & \[8855]  & (~\[17635]  | \[17986] );
  assign n4937 = ~preset & \[8840]  & (~\[17635]  | \[17986] );
  assign n4938 = ~preset & \[8825]  & (\[17999]  | ~\[18077] );
  assign n4939 = n3723 & (n3897 ? (n3910 ^ ~n3911) : (~n3910 ^ ~n3911));
  assign n4940 = ~preset & \[8780]  & (\[18311]  | ~\[18506] );
  assign n4941 = n3709 & (n3886 ? (n3923_1 ^ ~n3941) : (~n3923_1 ^ ~n3941));
  assign n4942 = ~preset & \[8735]  & (~n3798 | ~n5733);
  assign n4943 = ~preset & \[8720]  & (~n3798 | ~n5731);
  assign n4944 = n3718 & (n3885 ? (n3903_1 ^ ~n3920) : (~n3903_1 ^ ~n3920));
  assign n4945 = n3718 & (n3888_1 ? (n3901 ^ ~n3918_1) : (~n3901 ^ ~n3918_1));
  assign n4946 = ~preset & \[8675]  & (~\[18285]  | \[18363] );
  assign n4947 = ~preset & \[8660]  & (~\[18285]  | \[18363] );
  assign n4948 = n3706_1 & (n3895 ? (n3904 ^ ~n3905) : (~n3904 ^ ~n3905));
  assign n4949 = \[8630]  & n3707;
  assign n4950 = ~preset & \[8600]  & (\[17310]  | ~\[17388] );
  assign n4951 = ~preset & \[8585]  & (\[17310]  | ~\[17388] );
  assign n4952 = ~preset & \[8510]  & (~n3798 | ~n5731);
  assign n4953 = n5731 & n3798 & ~preset & pdata_3_3_;
  assign n4954 = ~preset & \[8495]  & (~\[17284]  | \[18376] );
  assign n4955 = ~preset & \[8480]  & (~\[17284]  | \[18376] );
  assign n4956 = ~preset & \[8465]  & (~\[17167]  | \[17362] );
  assign n4957 = ~preset & \[8390]  & (~\[17453]  | \[18246] );
  assign n4958 = ppeaka_1_1_ & (n5577 | n5720);
  assign n4959 = n3963 & \[4970]  & n3874_1;
  assign n4960 = ppeakp_1_1_ & (n5722 | n5723 | n5725);
  assign n4961 = n3801 & ppeakb_1_1_ & n3756;
  assign n4962 = ppeaka_8_8_ & (n5577 | n5720);
  assign n4963 = n3963 & \[13895]  & n3874_1;
  assign n4964 = ppeakp_8_8_ & (n5722 | n5723 | n5725);
  assign n4965 = n3801 & ppeakb_8_8_ & n3756;
  assign n4966 = n3857 & n3827_1 & \[12455]  & n3756;
  assign n4967 = n3963 & n3874_1 & \[12155]  & n3857;
  assign n4968 = n3857 & n3826 & \[14255]  & n3756;
  assign n4969 = n3857 & n3808 & \[4910]  & n3756;
  assign n4970 = n3857 & n3806 & \[5570]  & n3756;
  assign n4971 = n3857 & n3812_1 & \[14180]  & n3756;
  assign n4972 = n3857 & n3801 & \[10610]  & n3756;
  assign n4973 = n3876 & n3857 & \[12575]  & n3756;
  assign n4974 = n3857 & n3821 & \[8720]  & n3756;
  assign n4975 = n3857 & n3802_1 & \[9350]  & n3756;
  assign n4976 = n3857 & n3803 & \[6200]  & n3756;
  assign n4977 = n3857 & \[12845]  & n3702;
  assign n4978 = n3857 & n3800 & \[7385]  & n3756;
  assign n4979 = ppeaks_3_3_ & (n5708 | n5709);
  assign n4980 = n3801 & \[4565]  & n3756;
  assign n4981 = \[8330]  & (n3968 | n5701 | n5702);
  assign n4982 = \[12635]  & n3804 & (n5627 | n5628);
  assign n4983 = ~preset & \[8285]  & (~\[17180]  | \[17232] );
  assign n4984 = ~preset & \[8210]  & (~\[17635]  | \[17986] );
  assign n4985 = ~preset & \[8195]  & (~\[17635]  | \[17986] );
  assign n4986 = ~preset & \[8180]  & (\[17999]  | ~\[18077] );
  assign n4987 = ~preset & \[8150]  & (\[18311]  | ~\[18506] );
  assign n4988 = n3721_1 & (n3897 ? (n3910 ^ ~n3911) : (~n3910 ^ ~n3911));
  assign n4989 = ~preset & \[8135]  & (\[18311]  | ~\[18506] );
  assign n4990 = ~preset & \[8120]  & (\[18311]  | ~\[18506] );
  assign n4991 = n3709 & (n3889 ? (n3907 ^ ~n3908_1) : (~n3907 ^ ~n3908_1));
  assign n4992 = ~preset & \[8090]  & (~n3798 | ~n5733);
  assign n4993 = n4106 & (n3885 ? (n3903_1 ^ ~n3920) : (~n3903_1 ^ ~n3920));
  assign n4994 = ~preset & \[8075]  & (~n3798 | ~n5731);
  assign n4995 = n3718 & (n3897 ? (n3910 ^ ~n3911) : (~n3910 ^ ~n3911));
  assign n4996 = ~preset & \[8030]  & (~\[18285]  | \[18363] );
  assign n4997 = n3716_1 & (n3885 ? (n3903_1 ^ ~n3920) : (~n3903_1 ^ ~n3920));
  assign n4998 = ~preset & \[8015]  & (~\[18285]  | \[18363] );
  assign n4999 = n3716_1 & (n3887 ? (n3912 ^ ~n3913_1) : (~n3912 ^ ~n3913_1));
  assign n5000 = n3706_1 & (n3886 ? (n3923_1 ^ ~n3941) : (~n3923_1 ^ ~n3941));
  assign n5001 = ~preset & \[7955]  & (\[17310]  | ~\[17388] );
  assign n5002 = ~preset & \[7940]  & (\[17310]  | ~\[17388] );
  assign n5003 = ~preset & \[7880]  & (~n3798 | ~n5733);
  assign n5004 = n5733 & n3798 & ~preset & pdata_15_15_;
  assign n5005 = ~preset & \[7865]  & (~n3798 | ~n5731);
  assign n5006 = n5731 & n3798 & ~preset & pdata_6_6_;
  assign n5007 = ~preset & \[7850]  & (~\[17284]  | \[18376] );
  assign n5008 = ~preset & \[7835]  & (~\[17284]  | \[18376] );
  assign n5009 = ~preset & \[7820]  & (~\[17167]  | \[17362] );
  assign n5010 = ~preset & \[7805]  & (~\[17167]  | \[17362] );
  assign n5011 = ~preset & \[7745]  & (~\[17453]  | \[18246] );
  assign n5012 = ppeaka_2_2_ & (n5577 | n5720);
  assign n5013 = n3963 & ndout & n3874_1;
  assign n5014 = ppeakp_2_2_ & (n5722 | n5723 | n5725);
  assign n5015 = n3801 & ppeakb_2_2_ & n3756;
  assign n5016 = ppeaka_7_7_ & (n5577 | n5720);
  assign n5017 = n3963 & \[14285]  & n3874_1;
  assign n5018 = ppeakp_7_7_ & (n5722 | n5723 | n5725);
  assign n5019 = n3801 & ppeakb_7_7_ & n3756;
  assign n5020 = n3857 & n3827_1 & \[10700]  & n3756;
  assign n5021 = n3963 & n3874_1 & \[12035]  & n3857;
  assign n5022 = n3857 & n3826 & \[14690]  & n3756;
  assign n5023 = n3857 & n3808 & \[14240]  & n3756;
  assign n5024 = n3857 & n3806 & \[8885]  & n3756;
  assign n5025 = n3857 & n3812_1 & \[8090]  & n3756;
  assign n5026 = n3857 & n3801 & \[10340]  & n3756;
  assign n5027 = n3876 & n3857 & \[12815]  & n3756;
  assign n5028 = n3857 & n3821 & \[14990]  & n3756;
  assign n5029 = n3857 & n3802_1 & \[8705]  & n3756;
  assign n5030 = n3857 & n3803 & \[6890]  & n3756;
  assign n5031 = n3857 & \[12620]  & n3702;
  assign n5032 = n3857 & n3800 & \[8030]  & n3756;
  assign n5033 = ppeaks_13_13_ & (n5708 | n5709);
  assign n5034 = n3801 & \[6635]  & n3756;
  assign n5035 = \[7685]  & (n3968 | n5701 | n5702);
  assign n5036 = \[12410]  & n3804 & (n5627 | n5628);
  assign n5037 = ~preset & \[7655]  & (~\[17180]  | \[17232] );
  assign n5038 = ~preset & \[7640]  & (~\[17180]  | \[17232] );
  assign n5039 = ~preset & \[7580]  & (~\[17635]  | \[17986] );
  assign n5040 = ~preset & \[7565]  & (~\[17635]  | \[17986] );
  assign n5041 = ~preset & \[7550]  & (\[17999]  | ~\[18077] );
  assign n5042 = n3723 & (n3886 ? (n3923_1 ^ ~n3941) : (~n3923_1 ^ ~n3941));
  assign n5043 = n3721_1 & (n3895 ? (n3904 ^ ~n3905) : (~n3904 ^ ~n3905));
  assign n5044 = ~preset & \[7505]  & (\[18311]  | ~\[18506] );
  assign n5045 = ~preset & \[7490]  & (\[18311]  | ~\[18506] );
  assign n5046 = ~preset & \[7460]  & (~n3798 | ~n5733);
  assign n5047 = ~preset & \[7445]  & (~n3798 | ~n5731);
  assign n5048 = n4547 & (n3889 ? (n3907 ^ ~n3908_1) : (~n3907 ^ ~n3908_1));
  assign n5049 = n3718 & (n3895 ? (n3904 ^ ~n3905) : (~n3904 ^ ~n3905));
  assign n5050 = \[7415]  & n3717;
  assign n5051 = ~preset & \[7400]  & (~\[18285]  | \[18363] );
  assign n5052 = ~preset & \[7385]  & (~\[18285]  | \[18363] );
  assign n5053 = ~preset & \[7355]  & (\[18103]  | ~\[18168] );
  assign n5054 = n4160 & (n3886 ? (n3923_1 ^ ~n3941) : (~n3923_1 ^ ~n3941));
  assign n5055 = ~preset & \[7325]  & (\[17310]  | ~\[17388] );
  assign n5056 = ~preset & \[7310]  & (\[17310]  | ~\[17388] );
  assign n5057 = ~preset & \[7250]  & (~n3798 | ~n5733);
  assign n5058 = n5733 & n3798 & ~preset & pdata_14_14_;
  assign n5059 = ~preset & \[7235]  & (~n3798 | ~n5731);
  assign n5060 = n5731 & n3798 & ~preset & pdata_5_5_;
  assign n5061 = ~preset & \[7220]  & (~\[17284]  | \[18376] );
  assign n5062 = ~preset & \[7205]  & (~\[17167]  | \[17362] );
  assign n5063 = ~preset & \[7190]  & (~\[17167]  | \[17362] );
  assign n5064 = ~preset & \[7175]  & (~\[17167]  | \[17362] );
  assign n5065 = ~preset & \[7115]  & (~\[17453]  | \[18246] );
  assign n5066 = ppeaka_3_3_ & (n5577 | n5720);
  assign n5067 = n3963 & \[15785]  & n3874_1;
  assign n5068 = ppeakp_3_3_ & (n5722 | n5723 | n5725);
  assign n5069 = n3801 & ppeakb_3_3_ & n3756;
  assign n5070 = n3857 & n3827_1 & \[12920]  & n3756;
  assign n5071 = n3963 & n3874_1 & \[9665]  & n3857;
  assign n5072 = n3857 & n3826 & \[12005]  & n3756;
  assign n5073 = n3857 & n3808 & \[6305]  & n3756;
  assign n5074 = n3857 & n3806 & \[9830]  & n3756;
  assign n5075 = n3857 & n3812_1 & \[15020]  & n3756;
  assign n5076 = n3857 & n3801 & \[8120]  & n3756;
  assign n5077 = n3876 & n3857 & \[14570]  & n3756;
  assign n5078 = n3857 & n3821 & \[11150]  & n3756;
  assign n5079 = n3857 & n3802_1 & \[8045]  & n3756;
  assign n5080 = n3857 & n3803 & \[4805]  & n3756;
  assign n5081 = n3857 & \[12380]  & n3702;
  assign n5082 = n3857 & n3800 & \[8660]  & n3756;
  assign n5083 = ppeaks_1_1_ & (n5708 | n5709);
  assign n5084 = n3857 & n3827_1 & \[10415]  & n3756;
  assign n5085 = n3963 & n3874_1 & \[9680]  & n3857;
  assign n5086 = n3857 & n3826 & \[15065]  & n3756;
  assign n5087 = n3857 & n3808 & \[14660]  & n3756;
  assign n5088 = n3857 & n3806 & \[9845]  & n3756;
  assign n5089 = n3857 & n3812_1 & \[7460]  & n3756;
  assign n5090 = n3857 & n3801 & \[10625]  & n3756;
  assign n5091 = n3876 & n3857 & \[13775]  & n3756;
  assign n5092 = n3857 & n3821 & \[11615]  & n3756;
  assign n5093 = n3857 & n3802_1 & \[9365]  & n3756;
  assign n5094 = n3857 & n3803 & \[4820]  & n3756;
  assign n5095 = n3857 & \[12395]  & n3702;
  assign n5096 = n3857 & n3800 & \[8675]  & n3756;
  assign n5097 = ppeaks_12_12_ & (n5708 | n5709);
  assign n5098 = n3801 & \[5960]  & n3756;
  assign n5099 = \[7055]  & (n3968 | n5701 | n5702);
  assign n5100 = \[6245]  & n3804 & (n5627 | n5628);
  assign n5101 = \[7010]  & n3722;
  assign n5102 = ~preset & \[6965]  & (\[17037]  | ~\[18025] );
  assign n5103 = ~preset & \[6950]  & (\[17037]  | ~\[18025] );
  assign n5104 = ~preset & \[6935]  & (~\[17635]  | \[17986] );
  assign n5105 = ~preset & \[6920]  & (\[17999]  | ~\[18077] );
  assign n5106 = n3723 & (n3885 ? (n3903_1 ^ ~n3920) : (~n3903_1 ^ ~n3920));
  assign n5107 = n3723 & (n3887 ? (n3912 ^ ~n3913_1) : (~n3912 ^ ~n3913_1));
  assign n5108 = ~preset & \[6830]  & (~n3798 | ~n5733);
  assign n5109 = n4106 & (n3895 ? (n3904 ^ ~n3905) : (~n3904 ^ ~n3905));
  assign n5110 = ~preset & \[6815]  & (~n3798 | ~n5731);
  assign n5111 = n4547 & (n3886 ? (n3923_1 ^ ~n3941) : (~n3923_1 ^ ~n3941));
  assign n5112 = n3718 & (n3890 ? (n3921 ^ ~n3922) : (~n3921 ^ ~n3922));
  assign n5113 = ~preset & \[6770]  & (~\[18285]  | \[18363] );
  assign n5114 = n3716_1 & (n3890 ? (n3921 ^ ~n3922) : (~n3921 ^ ~n3922));
  assign n5115 = ~preset & \[6725]  & (\[18103]  | ~\[18168] );
  assign n5116 = n4160 & (n3895 ? (n3904 ^ ~n3905) : (~n3904 ^ ~n3905));
  assign n5117 = n4160 & (n3888_1 ? (n3901 ^ ~n3918_1) : (~n3901 ^ ~n3918_1));
  assign n5118 = ~preset & \[6680]  & (\[17310]  | ~\[17388] );
  assign n5119 = ~preset & \[6620]  & (~n3798 | ~n5733);
  assign n5120 = n5733 & n3798 & ~preset & pdata_13_13_;
  assign n5121 = ~preset & \[6605]  & (~n3798 | ~n5731);
  assign n5122 = n5731 & n3798 & ~preset & pdata_8_8_;
  assign n5123 = ~preset & \[6590]  & (~\[17284]  | \[18376] );
  assign n5124 = ~preset & \[6575]  & (~\[17284]  | \[18376] );
  assign n5125 = ~preset & \[6560]  & (~\[17167]  | \[17362] );
  assign n5126 = ~preset & \[6470]  & (~\[17453]  | \[18246] );
  assign n5127 = ppeaka_13_13_ & (n5577 | n5720);
  assign n5128 = n3963 & \[10760]  & n3874_1;
  assign n5129 = ppeakp_13_13_ & (n5722 | n5723 | n5725);
  assign n5130 = n3801 & ppeakb_13_13_ & n3756;
  assign n5131 = n3857 & n3827_1 & \[7625]  & n3756;
  assign n5132 = n3963 & n3874_1 & \[11300]  & n3857;
  assign n5133 = n3857 & n3826 & \[13865]  & n3756;
  assign n5134 = n3857 & n3808 & \[11690]  & n3756;
  assign n5135 = n3857 & n3806 & \[8870]  & n3756;
  assign n5136 = n3857 & n3812_1 & \[13085]  & n3756;
  assign n5137 = n3857 & n3801 & \[5495]  & n3756;
  assign n5138 = n3876 & n3857 & \[16085]  & n3756;
  assign n5139 = n3857 & n3821 & \[8075]  & n3756;
  assign n5140 = n3857 & n3802_1 & \[6110]  & n3756;
  assign n5141 = n3857 & n3803 & \[11165]  & n3756;
  assign n5142 = n3857 & \[14210]  & n3702;
  assign n5143 = n3857 & n3800 & \[10565]  & n3756;
  assign n5144 = ppeaks_6_6_ & (n5708 | n5709);
  assign n5145 = n3857 & n3827_1 & \[6320]  & n3756;
  assign n5146 = n3963 & n3874_1 & \[11780]  & n3857;
  assign n5147 = n3857 & n3826 & \[13880]  & n3756;
  assign n5148 = n3857 & n3808 & \[12425]  & n3756;
  assign n5149 = n3857 & n3806 & \[4880]  & n3756;
  assign n5150 = n3857 & n3812_1 & \[9395]  & n3756;
  assign n5151 = n3857 & n3801 & \[8150]  & n3756;
  assign n5152 = n3876 & n3857 & \[12365]  & n3756;
  assign n5153 = n3857 & n3821 & \[15725]  & n3756;
  assign n5154 = n3857 & n3802_1 & \[4730]  & n3756;
  assign n5155 = n3857 & n3803 & \[11180]  & n3756;
  assign n5156 = n3857 & \[15050]  & n3702;
  assign n5157 = n3857 & n3800 & \[10580]  & n3756;
  assign n5158 = ppeaks_15_15_ & (n5708 | n5709);
  assign n5159 = n3801 & \[7895]  & n3756;
  assign n5160 = \[6410]  & (n3968 | n5701 | n5702);
  assign n5161 = \[6920]  & n3804 & (n5627 | n5628);
  assign n5162 = n3966 & n3857 & ppeaka_2_2_ & n3756;
  assign n5163 = n3857 & n3812_1 & \[15290]  & n3756;
  assign n5164 = n3857 & n3801 & \[8555]  & n3756;
  assign n5165 = n3876 & n3857 & \[14465]  & n3756;
  assign n5166 = n3857 & n3821 & \[13640]  & n3756;
  assign n5167 = n3857 & n3802_1 & \[9140]  & n3756;
  assign n5168 = n3857 & n3803 & \[7310]  & n3756;
  assign n5169 = n3857 & \[15515]  & n3702;
  assign n5170 = n3857 & n3800 & \[4445]  & n3756;
  assign n5171 = ppeakb_2_2_ & ((n3756 & n3960) | n3968);
  assign n5172 = n3966 & n3857 & ppeaka_11_11_ & n3756;
  assign n5173 = n3857 & n3812_1 & \[5255]  & n3756;
  assign n5174 = n3857 & n3801 & \[4595]  & n3756;
  assign n5175 = n3876 & n3857 & \[14480]  & n3756;
  assign n5176 = n3857 & n3821 & \[5930]  & n3756;
  assign n5177 = n3857 & n3802_1 & \[9155]  & n3756;
  assign n5178 = n3857 & n3803 & \[14090]  & n3756;
  assign n5179 = n3857 & \[4295]  & n3702;
  assign n5180 = n3857 & n3800 & \[5855]  & n3756;
  assign n5181 = ppeakb_11_11_ & ((n3756 & n3960) | n3968);
  assign n5182 = \[6365]  & n3738;
  assign n5183 = \[6320]  & n3751;
  assign n5184 = ~preset & \[6290]  & (\[17037]  | ~\[18025] );
  assign n5185 = ~preset & \[6275]  & (\[17037]  | ~\[18025] );
  assign n5186 = ~preset & \[6260]  & (~\[17635]  | \[17986] );
  assign n5187 = ~preset & \[6245]  & (\[17999]  | ~\[18077] );
  assign n5188 = n3721_1 & (n3889 ? (n3907 ^ ~n3908_1) : (~n3907 ^ ~n3908_1));
  assign n5189 = ~preset & \[6185]  & (\[18311]  | ~\[18506] );
  assign n5190 = n3709 & (n3887 ? (n3912 ^ ~n3913_1) : (~n3912 ^ ~n3913_1));
  assign n5191 = ~preset & \[6155]  & (~n3798 | ~n5733);
  assign n5192 = n4106 & (n3897 ? (n3910 ^ ~n3911) : (~n3910 ^ ~n3911));
  assign n5193 = ~preset & \[6140]  & (~n3798 | ~n5731);
  assign n5194 = n4547 & (n3890 ? (n3921 ^ ~n3922) : (~n3921 ^ ~n3922));
  assign n5195 = ~preset & \[6125]  & (~n3798 | ~n5731);
  assign n5196 = ~preset & \[6095]  & (~\[18285]  | \[18363] );
  assign n5197 = n3716_1 & (n3886 ? (n3923_1 ^ ~n3941) : (~n3923_1 ^ ~n3941));
  assign n5198 = n3706_1 & (n3890 ? (n3921 ^ ~n3922) : (~n3921 ^ ~n3922));
  assign n5199 = ~preset & \[6050]  & (\[18103]  | ~\[18168] );
  assign n5200 = n3715 & (n3885 ? (n3903_1 ^ ~n3920) : (~n3903_1 ^ ~n3920));
  assign n5201 = n4160 & (n3897 ? (n3910 ^ ~n3911) : (~n3910 ^ ~n3911));
  assign n5202 = ~preset & \[6005]  & (\[17310]  | ~\[17388] );
  assign n5203 = ~preset & \[5945]  & (~n3798 | ~n5733);
  assign n5204 = n5733 & n3798 & ~preset & pdata_12_12_;
  assign n5205 = ~preset & \[5930]  & (~n3798 | ~n5731);
  assign n5206 = n5731 & n3798 & ~preset & pdata_11_11_;
  assign n5207 = ~preset & \[5915]  & (~n3798 | ~n5731);
  assign n5208 = n5731 & n3798 & ~preset & pdata_7_7_;
  assign n5209 = ~preset & \[5900]  & (~n3798 | ~n5731);
  assign n5210 = n5731 & n3798 & ~preset & pdata_0_0_;
  assign n5211 = ~preset & \[5885]  & (~\[17284]  | \[18376] );
  assign n5212 = ~preset & \[5870]  & (~\[17167]  | \[17362] );
  assign n5213 = ~preset & \[5780]  & (~\[17453]  | \[18246] );
  assign n5214 = ppeaka_12_12_ & (n5577 | n5720);
  assign n5215 = n3963 & \[11030]  & n3874_1;
  assign n5216 = ppeakp_12_12_ & (n5722 | n5723 | n5725);
  assign n5217 = n3801 & ppeakb_12_12_ & n3756;
  assign n5218 = n3857 & n3827_1 & \[8255]  & n3756;
  assign n5219 = n3963 & n3874_1 & \[11540]  & n3857;
  assign n5220 = n3857 & n3826 & \[12905]  & n3756;
  assign n5221 = n3857 & n3808 & \[10970]  & n3756;
  assign n5222 = n3857 & n3806 & \[8225]  & n3756;
  assign n5223 = n3857 & n3812_1 & \[12830]  & n3756;
  assign n5224 = n3857 & n3801 & \[4790]  & n3756;
  assign n5225 = n3876 & n3857 & \[15005]  & n3756;
  assign n5226 = n3857 & n3821 & \[6140]  & n3756;
  assign n5227 = n3857 & n3802_1 & \[6785]  & n3756;
  assign n5228 = n3857 & n3803 & \[11405]  & n3756;
  assign n5229 = n3857 & \[14630]  & n3702;
  assign n5230 = n3857 & n3800 & \[6770]  & n3756;
  assign n5231 = ppeaks_7_7_ & (n5708 | n5709);
  assign n5232 = n3857 & n3827_1 & \[10985]  & n3756;
  assign n5233 = n3963 & n3874_1 & \[11900]  & n3857;
  assign n5234 = n3857 & n3826 & \[14270]  & n3756;
  assign n5235 = n3857 & n3808 & \[12650]  & n3756;
  assign n5236 = n3857 & n3806 & \[9560]  & n3756;
  assign n5237 = n3857 & n3812_1 & \[8735]  & n3756;
  assign n5238 = n3857 & n3801 & \[10055]  & n3756;
  assign n5239 = n3876 & n3857 & \[13070]  & n3756;
  assign n5240 = n3857 & n3821 & \[16070]  & n3756;
  assign n5241 = n3857 & n3802_1 & \[5435]  & n3756;
  assign n5242 = n3857 & n3803 & \[6215]  & n3756;
  assign n5243 = n3857 & \[15410]  & n3702;
  assign n5244 = n3857 & n3800 & \[7400]  & n3756;
  assign n5245 = ppeaks_14_14_ & (n5708 | n5709);
  assign n5246 = n3801 & \[7265]  & n3756;
  assign n5247 = \[5720]  & (n3968 | n5701 | n5702);
  assign n5248 = \[7550]  & n3804 & (n5627 | n5628);
  assign n5249 = n3857 & n3811 & \[6350]  & n3756;
  assign n5250 = n3857 & n3819 & \[4475]  & n3756;
  assign n5251 = n3957_1 & n3857 & \[6410]  & n3756;
  assign n5252 = n3857 & n3808 & \[11225]  & n3756;
  assign n5253 = n3857 & n3806 & \[14405]  & n3756;
  assign n5254 = n3857 & n3803 & \[10175]  & n3756;
  assign n5255 = n3857 & n3800 & \[5135]  & n3756;
  assign n5256 = ppeaka_8_8_ & ((n3756 & n3801) | n3968);
  assign n5257 = n3966 & n3857 & ppeaka_10_10_ & n3756;
  assign n5258 = n3857 & n3812_1 & \[4550]  & n3756;
  assign n5259 = n3857 & n3801 & \[5300]  & n3756;
  assign n5260 = n3876 & n3857 & \[14060]  & n3756;
  assign n5261 = n3857 & n3821 & \[5225]  & n3756;
  assign n5262 = n3857 & n3802_1 & \[7220]  & n3756;
  assign n5263 = n3857 & n3803 & \[10850]  & n3756;
  assign n5264 = n3857 & \[5015]  & n3702;
  assign n5265 = n3857 & n3800 & \[15230]  & n3756;
  assign n5266 = ppeakb_10_10_ & ((n3756 & n3960) | n3968);
  assign n5267 = ~preset & \[5675]  & (~\[17791]  | \[17843] );
  assign n5268 = ~preset & \[5630]  & (~\[17180]  | \[17232] );
  assign n5269 = ~preset & \[5600]  & (\[17037]  | ~\[18025] );
  assign n5270 = ~preset & \[5555]  & (~\[17635]  | \[17986] );
  assign n5271 = n3723 & (n3895 ? (n3904 ^ ~n3905) : (~n3904 ^ ~n3905));
  assign n5272 = n3723 & (n3888_1 ? (n3901 ^ ~n3918_1) : (~n3901 ^ ~n3918_1));
  assign n5273 = ~preset & \[5495]  & (\[18311]  | ~\[18506] );
  assign n5274 = ~preset & \[5465]  & (~n3798 | ~n5733);
  assign n5275 = ~preset & \[5450]  & (~n3798 | ~n5731);
  assign n5276 = n4547 & (n3897 ? (n3910 ^ ~n3911) : (~n3910 ^ ~n3911));
  assign n5277 = n3718 & (n3889 ? (n3907 ^ ~n3908_1) : (~n3907 ^ ~n3908_1));
  assign n5278 = ~preset & \[5405]  & (~\[18285]  | \[18363] );
  assign n5279 = ~preset & \[5390]  & (~\[18285]  | \[18363] );
  assign n5280 = n3706_1 & (n3887 ? (n3912 ^ ~n3913_1) : (~n3912 ^ ~n3913_1));
  assign n5281 = ~preset & \[5360]  & (\[18103]  | ~\[18168] );
  assign n5282 = n4160 & (n3885 ? (n3903_1 ^ ~n3920) : (~n3903_1 ^ ~n3920));
  assign n5283 = \[5330]  & n3713;
  assign n5284 = ~preset & \[5315]  & (\[17310]  | ~\[17388] );
  assign n5285 = ~preset & \[5255]  & (~n3798 | ~n5733);
  assign n5286 = n5733 & n3798 & ~preset & pdata_11_11_;
  assign n5287 = ~preset & \[5240]  & (~n3798 | ~n5732);
  assign n5288 = n5732 & n3798 & ~preset & pdata_5_5_;
  assign n5289 = ~preset & \[5225]  & (~n3798 | ~n5731);
  assign n5290 = n5731 & n3798 & ~preset & pdata_10_10_;
  assign n5291 = ~preset & \[5210]  & (~\[17284]  | \[18376] );
  assign n5292 = ~preset & \[5195]  & (~\[17284]  | \[18376] );
  assign n5293 = ~preset & \[5180]  & (~\[17167]  | \[17362] );
  assign n5294 = ~preset & \[5120]  & (~\[17102]  | \[17154] );
  assign n5295 = ~preset & \[5105]  & (~\[17102]  | \[17154] );
  assign n5296 = ~preset & \[5090]  & (~\[17453]  | \[18246] );
  assign n5297 = ~preset & \[5075]  & (~\[17453]  | \[18246] );
  assign n5298 = ppeaka_11_11_ & (n5577 | n5720);
  assign n5299 = n3963 & \[12020]  & n3874_1;
  assign n5300 = ppeakp_11_11_ & (n5722 | n5723 | n5725);
  assign n5301 = n3801 & ppeakb_11_11_ & n3756;
  assign n5302 = n3857 & n3827_1 & \[12245]  & n3756;
  assign n5303 = n3963 & n3874_1 & \[11765]  & n3857;
  assign n5304 = n3857 & n3826 & \[14675]  & n3756;
  assign n5305 = n3857 & n3808 & \[5615]  & n3756;
  assign n5306 = n3857 & n3806 & \[4865]  & n3756;
  assign n5307 = n3857 & n3812_1 & \[13790]  & n3756;
  assign n5308 = n3857 & n3801 & \[9785]  & n3756;
  assign n5309 = n3876 & n3857 & \[12350]  & n3756;
  assign n5310 = n3857 & n3821 & \[9380]  & n3756;
  assign n5311 = n3857 & n3802_1 & \[4715]  & n3756;
  assign n5312 = n3857 & n3803 & \[6875]  & n3756;
  assign n5313 = n3857 & \[15035]  & n3702;
  assign n5314 = n3857 & n3800 & \[8015]  & n3756;
  assign n5315 = ppeaks_4_4_ & (n5708 | n5709);
  assign n5316 = n3801 & \[9185]  & n3756;
  assign n5317 = \[5030]  & (n3968 | n5701 | n5702);
  assign n5318 = \[13835]  & n3804 & (n5627 | n5628);
  assign n5319 = n3801 & \[9200]  & n3756;
  assign n5320 = \[5015]  & (n3968 | n5701 | n5702);
  assign n5321 = \[8180]  & n3804 & (n5627 | n5628);
  assign n5322 = n3857 & n3811 & \[7025]  & n3756;
  assign n5323 = n3857 & n3819 & \[5180]  & n3756;
  assign n5324 = n3957_1 & n3857 & \[7055]  & n3756;
  assign n5325 = n3857 & n3808 & \[10970]  & n3756;
  assign n5326 = n3857 & n3806 & \[13985]  & n3756;
  assign n5327 = n3857 & n3803 & \[10460]  & n3756;
  assign n5328 = n3857 & n3800 & \[4430]  & n3756;
  assign n5329 = ppeaka_7_7_ & ((n3756 & n3801) | n3968);
  assign n5330 = n3966 & n3857 & ppeaka_0_0_ & n3756;
  assign n5331 = n3857 & n3812_1 & \[15995]  & n3756;
  assign n5332 = n3857 & n3801 & \[4580]  & n3756;
  assign n5333 = n3876 & n3857 & \[13655]  & n3756;
  assign n5334 = n3857 & n3821 & \[5900]  & n3756;
  assign n5335 = n3857 & n3802_1 & \[7835]  & n3756;
  assign n5336 = n3857 & n3803 & \[10550]  & n3756;
  assign n5337 = n3857 & \[4310]  & n3702;
  assign n5338 = n3857 & n3800 & \[15605]  & n3756;
  assign n5339 = ppeakb_0_0_ & ((n3756 & n3960) | n3968);
  assign n5340 = ~preset & \[4970]  & (~\[17791]  | \[17843] );
  assign n5341 = ~preset & \[4895]  & (\[17037]  | ~\[18025] );
  assign n5342 = \[4880]  & n3729;
  assign n5343 = n3804 & ~\[17986]  & \[11915]  & \[17635] ;
  assign n5344 = ppeakp_11_11_ & (n3807_1 | (~n3804 & n3805));
  assign n5345 = ~\[17648]  & \[16100]  & \[17427] ;
  assign n5346 = ~\[17232]  & \[10130]  & \[17180] ;
  assign n5347 = n3811 & n3798 & ppeaka_11_11_ & ~\[17245] ;
  assign n5348 = \[18077]  & \[13115]  & ~\[17999] ;
  assign n5349 = n3803 & n3798 & ppeakb_11_11_ & ~\[16933] ;
  assign n5350 = n3804 & ~\[17986]  & \[12050]  & \[17635] ;
  assign n5351 = ppeakp_12_12_ & (n3807_1 | (~n3804 & n3805));
  assign n5352 = ~\[17648]  & \[15755]  & \[17427] ;
  assign n5353 = ~\[17232]  & \[10415]  & \[17180] ;
  assign n5354 = n3811 & n3798 & ppeaka_12_12_ & ~\[17245] ;
  assign n5355 = \[18077]  & \[12395]  & ~\[17999] ;
  assign n5356 = n3803 & n3798 & ppeakb_12_12_ & ~\[16933] ;
  assign n5357 = n3804 & ~\[17986]  & \[12170]  & \[17635] ;
  assign n5358 = ppeakp_13_13_ & (n3807_1 | (~n3804 & n3805));
  assign n5359 = ~\[17648]  & \[13805]  & \[17427] ;
  assign n5360 = ~\[17232]  & \[10700]  & \[17180] ;
  assign n5361 = n3811 & n3798 & ppeaka_13_13_ & ~\[17245] ;
  assign n5362 = \[18077]  & \[12620]  & ~\[17999] ;
  assign n5363 = n3803 & n3798 & ppeakb_13_13_ & ~\[16933] ;
  assign n5364 = n3804 & ~\[17986]  & \[12260]  & \[17635] ;
  assign n5365 = ppeakp_14_14_ & (n3807_1 | (~n3804 & n3805));
  assign n5366 = ~\[17648]  & \[13445]  & \[17427] ;
  assign n5367 = ~\[17232]  & \[10985]  & \[17180] ;
  assign n5368 = n3811 & n3798 & ppeaka_14_14_ & ~\[17245] ;
  assign n5369 = \[18077]  & \[15410]  & ~\[17999] ;
  assign n5370 = n3803 & n3798 & ppeakb_14_14_ & ~\[16933] ;
  assign n5371 = n3804 & ~\[17986]  & \[12470]  & \[17635] ;
  assign n5372 = ppeakp_15_15_ & (n3807_1 | (~n3804 & n3805));
  assign n5373 = ~\[17648]  & \[14615]  & \[17427] ;
  assign n5374 = ~\[17232]  & \[6320]  & \[17180] ;
  assign n5375 = n3811 & n3798 & ppeaka_15_15_ & ~\[17245] ;
  assign n5376 = \[18077]  & \[15050]  & ~\[17999] ;
  assign n5377 = n3803 & n3798 & ppeakb_15_15_ & ~\[16933] ;
  assign n5378 = ~preset & \[4850]  & (~\[17635]  | \[17986] );
  assign n5379 = n3804 & ~\[17986]  & \[11075]  & \[17635] ;
  assign n5380 = ppeakp_7_7_ & (n3807_1 | (~n3804 & n3805));
  assign n5381 = ~\[17648]  & \[5540]  & \[17427] ;
  assign n5382 = ~\[17232]  & \[8255]  & \[17180] ;
  assign n5383 = n3811 & n3798 & ppeaka_7_7_ & ~\[17245] ;
  assign n5384 = \[18077]  & \[14630]  & ~\[17999] ;
  assign n5385 = n3803 & n3798 & ppeakb_7_7_ & ~\[16933] ;
  assign n5386 = n3804 & ~\[17986]  & \[11330]  & \[17635] ;
  assign n5387 = ppeakp_8_8_ & (n3807_1 | (~n3804 & n3805));
  assign n5388 = ~\[17648]  & \[11420]  & \[17427] ;
  assign n5389 = ~\[17232]  & \[8915]  & \[17180] ;
  assign n5390 = n3811 & n3798 & ppeaka_8_8_ & ~\[17245] ;
  assign n5391 = \[18077]  & \[13460]  & ~\[17999] ;
  assign n5392 = n3803 & n3798 & ppeakb_8_8_ & ~\[16933] ;
  assign n5393 = n3804 & ~\[17986]  & \[11570]  & \[17635] ;
  assign n5394 = ppeakp_9_9_ & (n3807_1 | (~n3804 & n3805));
  assign n5395 = ~\[17648]  & \[11645]  & \[17427] ;
  assign n5396 = ~\[17232]  & \[9590]  & \[17180] ;
  assign n5397 = n3811 & n3798 & ppeaka_9_9_ & ~\[17245] ;
  assign n5398 = \[18077]  & \[13820]  & ~\[17999] ;
  assign n5399 = n3803 & n3798 & ppeakb_9_9_ & ~\[16933] ;
  assign n5400 = n3804 & ~\[17986]  & \[11795]  & \[17635] ;
  assign n5401 = ppeakp_10_10_ & (n3807_1 | (~n3804 & n3805));
  assign n5402 = ~\[17648]  & \[10925]  & \[17427] ;
  assign n5403 = ~\[17232]  & \[9860]  & \[17180] ;
  assign n5404 = n3811 & n3798 & ppeaka_10_10_ & ~\[17245] ;
  assign n5405 = \[18077]  & \[12860]  & ~\[17999] ;
  assign n5406 = n3803 & n3798 & ppeakb_10_10_ & ~\[16933] ;
  assign n5407 = n3803 & n3798 & ppeaka_0_0_ & ~\[16933] ;
  assign n5408 = n3804 & ~\[17986]  & \[11555]  & \[17635] ;
  assign n5409 = ppeakp_0_0_ & (n3807_1 | (~n3804 & n3805));
  assign n5410 = ~\[17648]  & \[11630]  & \[17427] ;
  assign n5411 = ~\[17232]  & \[13175]  & \[17180] ;
  assign n5412 = n3811 & n3798 & ppeaka_0_0_ & ~\[17245] ;
  assign n5413 = \[18077]  & \[12605]  & ~\[17999] ;
  assign n5414 = n3803 & n3798 & ppeakb_0_0_ & ~\[16933] ;
  assign n5415 = n3804 & ~\[17986]  & \[11315]  & \[17635] ;
  assign n5416 = ppeakp_1_1_ & (n3807_1 | (~n3804 & n3805));
  assign n5417 = ~\[17648]  & \[9485]  & \[17427] ;
  assign n5418 = ~\[17232]  & \[12920]  & \[17180] ;
  assign n5419 = n3811 & n3798 & ppeaka_1_1_ & ~\[17245] ;
  assign n5420 = \[18077]  & \[12380]  & ~\[17999] ;
  assign n5421 = n3803 & n3798 & ppeakb_1_1_ & ~\[16933] ;
  assign n5422 = n3804 & ~\[17986]  & \[11060]  & \[17635] ;
  assign n5423 = ppeakp_2_2_ & (n3807_1 | (~n3804 & n3805));
  assign n5424 = ~\[17648]  & \[7535]  & \[17427] ;
  assign n5425 = ~\[17232]  & \[12680]  & \[17180] ;
  assign n5426 = n3811 & n3798 & ppeaka_2_2_ & ~\[17245] ;
  assign n5427 = \[18077]  & \[13100]  & ~\[17999] ;
  assign n5428 = n3803 & n3798 & ppeakb_2_2_ & ~\[16933] ;
  assign n5429 = n3804 & ~\[17986]  & \[10790]  & \[17635] ;
  assign n5430 = ppeakp_3_3_ & (n3807_1 | (~n3804 & n3805));
  assign n5431 = ~\[17648]  & \[8165]  & \[17427] ;
  assign n5432 = ~\[17232]  & \[12455]  & \[17180] ;
  assign n5433 = n3811 & n3798 & ppeaka_3_3_ & ~\[17245] ;
  assign n5434 = \[18077]  & \[12845]  & ~\[17999] ;
  assign n5435 = n3803 & n3798 & ppeakb_3_3_ & ~\[16933] ;
  assign n5436 = n3804 & ~\[17986]  & \[10505]  & \[17635] ;
  assign n5437 = ppeakp_4_4_ & (n3807_1 | (~n3804 & n3805));
  assign n5438 = ~\[17648]  & \[6230]  & \[17427] ;
  assign n5439 = ~\[17232]  & \[12245]  & \[17180] ;
  assign n5440 = n3811 & n3798 & ppeaka_4_4_ & ~\[17245] ;
  assign n5441 = \[18077]  & \[15035]  & ~\[17999] ;
  assign n5442 = n3803 & n3798 & ppeakb_4_4_ & ~\[16933] ;
  assign n5443 = n3804 & ~\[17986]  & \[10220]  & \[17635] ;
  assign n5444 = ppeakp_5_5_ & (n3807_1 | (~n3804 & n3805));
  assign n5445 = ~\[17648]  & \[6905]  & \[17427] ;
  assign n5446 = ~\[17232]  & \[6995]  & \[17180] ;
  assign n5447 = n3811 & n3798 & ppeaka_5_5_ & ~\[17245] ;
  assign n5448 = \[18077]  & \[15395]  & ~\[17999] ;
  assign n5449 = n3803 & n3798 & ppeakb_5_5_ & ~\[16933] ;
  assign n5450 = n3804 & ~\[17986]  & \[9950]  & \[17635] ;
  assign n5451 = ppeakp_6_6_ & (n3807_1 | (~n3804 & n3805));
  assign n5452 = ~\[17648]  & \[4835]  & \[17427] ;
  assign n5453 = ~\[17232]  & \[7625]  & \[17180] ;
  assign n5454 = n3811 & n3798 & ppeaka_6_6_ & ~\[17245] ;
  assign n5455 = \[18077]  & \[14210]  & ~\[17999] ;
  assign n5456 = n3803 & n3798 & ppeakb_6_6_ & ~\[16933] ;
  assign n5457 = n3721_1 & (n3890 ? (n3921 ^ ~n3922) : (~n3921 ^ ~n3922));
  assign n5458 = ~preset & \[4790]  & (\[18311]  | ~\[18506] );
  assign n5459 = n3709 & (n3885 ? (n3903_1 ^ ~n3920) : (~n3903_1 ^ ~n3920));
  assign n5460 = n3709 & (n3888_1 ? (n3901 ^ ~n3918_1) : (~n3901 ^ ~n3918_1));
  assign n5461 = ~preset & \[4745]  & (~n3798 | ~n5731);
  assign n5462 = n5788 & ~n5468 & ~n5784;
  assign n5463 = ~ppeaka_15_15_ & (~n3950 | (~n5532 & ~n5533));
  assign n5464 = ~\[18363]  & \[6755]  & \[18285] ;
  assign n5465 = n3800 & n3798 & ppeaka_15_15_ & ~\[18285] ;
  assign n5466 = n5730 & n5729 & ppeakb_15_15_ & n3798;
  assign n5467 = n3801 & n3798 & \[13550]  & ~\[18506] ;
  assign n5468 = ~ppeaka_14_14_ & (~n3950 | (~n5532 & ~n5533));
  assign n5469 = ~\[18363]  & \[9740]  & \[18285] ;
  assign n5470 = n3800 & n3798 & ppeaka_13_13_ & ~\[18285] ;
  assign n5471 = n5730 & n5729 & ppeakb_13_13_ & n3798;
  assign n5472 = n3801 & n3798 & \[15500]  & ~\[18506] ;
  assign n5473 = ~\[18363]  & \[6080]  & \[18285] ;
  assign n5474 = n3800 & n3798 & ppeaka_14_14_ & ~\[18285] ;
  assign n5475 = n5730 & n5729 & ppeakb_14_14_ & n3798;
  assign n5476 = n3801 & n3798 & \[15140]  & ~\[18506] ;
  assign n5477 = n3718 & (n3887 ? (n3912 ^ ~n3913_1) : (~n3912 ^ ~n3913_1));
  assign n5478 = ~preset & \[4700]  & (~\[18285]  | \[18363] );
  assign n5479 = n3716_1 & (n3897 ? (n3910 ^ ~n3911) : (~n3910 ^ ~n3911));
  assign n5480 = n3706_1 & (n3889 ? (n3907 ^ ~n3908_1) : (~n3907 ^ ~n3908_1));
  assign n5481 = ~preset & \[4655]  & (\[18103]  | ~\[18168] );
  assign n5482 = n3715 & (n3895 ? (n3904 ^ ~n3905) : (~n3904 ^ ~n3905));
  assign n5483 = n3906 & ((n3910 & n3911) | (n3897 & (n3910 | n3911)));
  assign n5484 = n3895 & (n5534 | n5535 | n5536);
  assign n5485 = n3942 & ((n3921 & n3922) | (n3890 & (n3921 | n3922)));
  assign n5486 = n3886 & n3941;
  assign n5487 = n3909 & ((n3912 & n3913_1) | (n3887 & (n3912 | n3913_1)));
  assign n5488 = n3889 & (n5539 | n5749);
  assign n5489 = ~\[18363]  & \[9725]  & \[18285] ;
  assign n5490 = n3800 & n3798 & ppeaka_2_2_ & ~\[18285] ;
  assign n5491 = n5730 & n5729 & ppeakb_2_2_ & n3798;
  assign n5492 = n3801 & n3798 & \[15515]  & ~\[18506] ;
  assign n5493 = ~ppeaka_3_3_ & ~n5541 & (n3792_1 | n3900);
  assign n5494 = ~\[18363]  & \[9995]  & \[18285] ;
  assign n5495 = n3800 & n3798 & ppeaka_3_3_ & ~\[18285] ;
  assign n5496 = n5730 & n5729 & ppeakb_3_3_ & n3798;
  assign n5497 = n3801 & n3798 & \[15860]  & ~\[18506] ;
  assign n5498 = ~\[18363]  & \[5375]  & \[18285] ;
  assign n5499 = n3800 & n3798 & ppeaka_4_4_ & ~\[18285] ;
  assign n5500 = n5730 & n5729 & ppeakb_4_4_ & n3798;
  assign n5501 = n3801 & n3798 & \[14765]  & ~\[18506] ;
  assign n5502 = ~\[18363]  & \[4670]  & \[18285] ;
  assign n5503 = n3800 & n3798 & ppeaka_5_5_ & ~\[18285] ;
  assign n5504 = n5730 & n5729 & ppeakb_5_5_ & n3798;
  assign n5505 = n3801 & n3798 & \[8330]  & ~\[18506] ;
  assign n5506 = ~\[18363]  & \[6740]  & \[18285] ;
  assign n5507 = n3800 & n3798 & ppeaka_6_6_ & ~\[18285] ;
  assign n5508 = n5730 & n5729 & ppeakb_6_6_ & n3798;
  assign n5509 = n3801 & n3798 & \[7685]  & ~\[18506] ;
  assign n5510 = ~\[18363]  & \[6065]  & \[18285] ;
  assign n5511 = n3800 & n3798 & ppeaka_7_7_ & ~\[18285] ;
  assign n5512 = n5730 & n5729 & ppeakb_7_7_ & n3798;
  assign n5513 = n3801 & n3798 & \[7055]  & ~\[18506] ;
  assign n5514 = ~\[18363]  & \[8000]  & \[18285] ;
  assign n5515 = n3800 & n3798 & ppeaka_8_8_ & ~\[18285] ;
  assign n5516 = n5730 & n5729 & ppeakb_8_8_ & n3798;
  assign n5517 = n3801 & n3798 & \[6410]  & ~\[18506] ;
  assign n5518 = ~n5537 & ~n3941 & ~ppeaka_8_8_ & ppeaka_9_9_;
  assign n5519 = ~ppeaka_9_9_ & ~n5537 & (ppeaka_8_8_ | n3941);
  assign n5520 = ~\[18363]  & \[7370]  & \[18285] ;
  assign n5521 = n3800 & n3798 & ppeaka_9_9_ & ~\[18285] ;
  assign n5522 = n5730 & n5729 & ppeakb_9_9_ & n3798;
  assign n5523 = n3801 & n3798 & \[5720]  & ~\[18506] ;
  assign n5524 = ~\[18363]  & \[9305]  & \[18285] ;
  assign n5525 = n3800 & n3798 & ppeaka_10_10_ & ~\[18285] ;
  assign n5526 = n5730 & n5729 & ppeakb_10_10_ & n3798;
  assign n5527 = n3801 & n3798 & \[5015]  & ~\[18506] ;
  assign n5528 = ~\[18363]  & \[8645]  & \[18285] ;
  assign n5529 = n3800 & n3798 & ppeaka_11_11_ & ~\[18285] ;
  assign n5530 = n5730 & n5729 & ppeakb_11_11_ & n3798;
  assign n5531 = n3801 & n3798 & \[4295]  & ~\[18506] ;
  assign n5532 = ~n5536 & ~n5534 & ~n5535 & n5753;
  assign n5533 = ~n3792_1 & (n3949 | (~n3941 & n5751));
  assign n5534 = n5752 & (n5537 | (~n3941 & n5751));
  assign n5535 = n3954 & ~n5537 & (n3941 | ~n5751);
  assign n5536 = ~ppeaka_11_11_ & ~n3952;
  assign n5537 = n3949 & (~n3798 | ~n5729 | ~n5730);
  assign n5538 = ~n3792_1 & (~n3900 | n5541);
  assign n5539 = n3948_1 & (n3792_1 | n3900) & ~n5541;
  assign n5540 = ~ppeaka_5_5_ & ~n3947;
  assign n5541 = ~n5545 & ~n5543 & ~n5544 & n5747;
  assign n5542 = ~n3900 & (~n3798 | ~n5729 | ~n5730);
  assign n5543 = ~n5739 & ~n3878_1 & ~n5737 & n5746;
  assign n5544 = n3946 & (n3878_1 | n5737 | n5739);
  assign n5545 = ~ppeaka_2_2_ & ~n3945;
  assign n5546 = ~\[18363]  & \[10010]  & \[18285] ;
  assign n5547 = n3800 & n3798 & ppeaka_12_12_ & ~\[18285] ;
  assign n5548 = n5730 & n5729 & ppeakb_12_12_ & n3798;
  assign n5549 = n3801 & n3798 & \[15845]  & ~\[18506] ;
  assign n5550 = n5730 & n5729 & ppeaka_0_0_ & n3798;
  assign n5551 = ~\[18363]  & \[8630]  & \[18285] ;
  assign n5552 = n3800 & n3798 & ppeaka_0_0_ & ~\[18285] ;
  assign n5553 = n5730 & n5729 & ppeakb_0_0_ & n3798;
  assign n5554 = n3801 & n3798 & \[4310]  & ~\[18506] ;
  assign n5555 = ~\[18363]  & \[9290]  & \[18285] ;
  assign n5556 = n3800 & n3798 & ppeaka_1_1_ & ~\[18285] ;
  assign n5557 = n5730 & n5729 & ppeakb_1_1_ & n3798;
  assign n5558 = n3801 & n3798 & \[5030]  & ~\[18506] ;
  assign n5559 = ~preset & \[4610]  & (\[17310]  | ~\[17388] );
  assign n5560 = ~preset & \[4550]  & (~n3798 | ~n5733);
  assign n5561 = n5733 & n3798 & ~preset & pdata_10_10_;
  assign n5562 = ~preset & \[4535]  & (~n3798 | ~n5732);
  assign n5563 = n5732 & n3798 & ~preset & pdata_15_15_;
  assign n5564 = ~preset & \[4520]  & (~n3798 | ~n5731);
  assign n5565 = n5731 & n3798 & ~preset & pdata_9_9_;
  assign n5566 = ~preset & \[4505]  & (~\[17284]  | \[18376] );
  assign n5567 = ~preset & \[4490]  & (~\[17284]  | \[18376] );
  assign n5568 = ~preset & \[4475]  & (~\[17167]  | \[17362] );
  assign n5569 = ~preset & \[4415]  & (~\[17102]  | \[17154] );
  assign n5570 = ~preset & \[4400]  & (~\[17102]  | \[17154] );
  assign n5571 = ~preset & \[4370]  & (~\[17453]  | \[18246] );
  assign n5572 = ~preset & \[4355]  & (~\[17453]  | \[18246] );
  assign n5573 = ppeaka_10_10_ & (n5577 | n5720);
  assign n5574 = n3963 & \[12140]  & n3874_1;
  assign n5575 = ppeakp_10_10_ & (n5722 | n5723 | n5725);
  assign n5576 = n3801 & ppeakb_10_10_ & n3756;
  assign n5577 = n3899 & n3756 & n3876;
  assign n5578 = ~n3899 & n3756 & n3876;
  assign n5579 = n3857 & n3827_1 & \[6995]  & n3756;
  assign n5580 = n3963 & n3874_1 & \[11885]  & n3857;
  assign n5581 = n3857 & n3826 & \[13505]  & n3756;
  assign n5582 = n3857 & n3808 & \[11465]  & n3756;
  assign n5583 = n3857 & n3806 & \[9545]  & n3756;
  assign n5584 = n3857 & n3812_1 & \[13430]  & n3756;
  assign n5585 = n3857 & n3801 & \[6185]  & n3756;
  assign n5586 = n3876 & n3857 & \[13055]  & n3756;
  assign n5587 = n3857 & n3821 & \[7445]  & n3756;
  assign n5588 = n3857 & n3802_1 & \[5420]  & n3756;
  assign n5589 = n3857 & n3803 & \[10895]  & n3756;
  assign n5590 = n3857 & \[15395]  & n3702;
  assign n5591 = n3857 & n3800 & \[10280]  & n3756;
  assign n5592 = ppeaks_5_5_ & (n5708 | n5709);
  assign n5593 = n3801 & \[8525]  & n3756;
  assign n5594 = \[4310]  & (n3968 | n5701 | n5702);
  assign n5595 = \[14225]  & n3804 & (n5627 | n5628);
  assign n5596 = n3801 & \[8540]  & n3756;
  assign n5597 = \[4295]  & (n3968 | n5701 | n5702);
  assign n5598 = \[8825]  & n3804 & (n5627 | n5628);
  assign n5599 = n3857 & n3811 & \[4955]  & n3756;
  assign n5600 = n3857 & n3819 & \[5870]  & n3756;
  assign n5601 = n3957_1 & n3857 & \[7685]  & n3756;
  assign n5602 = n3857 & n3808 & \[11690]  & n3756;
  assign n5603 = n3857 & n3806 & \[15200]  & n3756;
  assign n5604 = n3857 & n3803 & \[10745]  & n3756;
  assign n5605 = n3857 & n3800 & \[15935]  & n3756;
  assign n5606 = ppeaka_6_6_ & ((n3756 & n3801) | n3968);
  assign n5607 = n3966 & n3857 & ppeaka_1_1_ & n3756;
  assign n5608 = n3857 & n3812_1 & \[15650]  & n3756;
  assign n5609 = n3857 & n3801 & \[5285]  & n3756;
  assign n5610 = n3876 & n3857 & \[13310]  & n3756;
  assign n5611 = n3857 & n3821 & \[13295]  & n3756;
  assign n5612 = n3857 & n3802_1 & \[8480]  & n3756;
  assign n5613 = n3857 & n3803 & \[14510]  & n3756;
  assign n5614 = n3857 & \[5030]  & n3702;
  assign n5615 = n3857 & n3800 & \[5150]  & n3756;
  assign n5616 = ppeakb_1_1_ & ((n3756 & n3960) | n3968);
  assign n5617 = n3966 & n3857 & ppeaka_12_12_ & n3756;
  assign n5618 = n3857 & n3812_1 & \[5945]  & n3756;
  assign n5619 = n3857 & n3801 & \[9230]  & n3756;
  assign n5620 = n3876 & n3857 & \[13325]  & n3756;
  assign n5621 = n3857 & n3821 & \[15260]  & n3756;
  assign n5622 = n3857 & n3802_1 & \[8495]  & n3756;
  assign n5623 = n3857 & n3803 & \[7955]  & n3756;
  assign n5624 = n3857 & \[15845]  & n3702;
  assign n5625 = n3857 & n3800 & \[6545]  & n3756;
  assign n5626 = ppeakb_12_12_ & ((n3756 & n3960) | n3968);
  assign n5627 = ~n3955 & ~\[17089]  & ~preset & pdn;
  assign n5628 = n3790 & ~preset & ~\[17596] ;
  assign n5629 = n5686 & (n3799 | (~\[17596]  & n3790));
  assign n5630 = n3955 & pdn & ~\[17089] ;
  assign n5631 = ~\[17856]  & \[18207] ;
  assign n5632 = ~preset & ndout & (~\[17791]  | \[17843] );
  assign n5633 = ~\[17752]  & ~ppeaki_6_6_ & ~ppeaki_7_7_;
  assign n5634 = \[17752]  & ~\[17544]  & \[17713] ;
  assign n5635 = \[17674]  & \[17609] ;
  assign n5636 = \[17752]  & \[17544]  & \[17713] ;
  assign n5637 = ppeaki_6_6_ & ~ppeaki_4_4_;
  assign n5638 = ~\[17713]  & ~\[17674] ;
  assign n5639 = ~ppeaki_5_5_ & ppeaki_4_4_;
  assign n5640 = \[17713]  & \[17609] ;
  assign n5641 = \[17713]  & ~\[17609]  & \[17674] ;
  assign n5642 = ~\[17752]  & ppeaki_6_6_ & ~ppeaki_7_7_;
  assign n5643 = ~\[17713]  & \[17674] ;
  assign n5644 = ~ppeaki_5_5_ & ~ppeaki_4_4_;
  assign n5645 = ~\[17713]  & \[17609] ;
  assign n5646 = \[17674]  & \[17609] ;
  assign n5647 = \[17752]  & \[17544]  & ~\[17713] ;
  assign n5648 = ~ppeaki_5_5_ & ~ppeaki_4_4_;
  assign n5649 = ~\[17713]  & ~\[17609] ;
  assign n5650 = ppeaki_6_6_ & ppeaki_4_4_;
  assign n5651 = \[17713]  & ~\[17674] ;
  assign n5652 = ~ppeaki_5_5_ & ppeaki_4_4_;
  assign n5653 = \[17713]  & ~\[17609] ;
  assign n5654 = ~\[17752]  & ppeaki_6_6_ & ~ppeaki_7_7_;
  assign n5655 = \[17713]  & \[17674] ;
  assign n5656 = ~\[17713]  & ~\[17609]  & \[17674] ;
  assign n5657 = ~\[17752]  & ~ppeaki_6_6_ & ~ppeaki_7_7_;
  assign n5658 = \[17752]  & ~\[17544]  & ~\[17713] ;
  assign n5659 = n3843 | n3842_1;
  assign n5660 = n3830 | n3831 | n3832_1 | n3833;
  assign n5661 = n3834 | n3835 | n3836 | n3837_1;
  assign n5662 = n3838 | n3839 | n3840 | n3841;
  assign n5663 = ~\[18636]  & ~\[18597]  & \[17596]  & ~\[17661] ;
  assign n5664 = ~n3828 & n5663 & (n3875 | n3881);
  assign n5665 = ~\[18636]  & ~\[18597]  & \[17596]  & ~\[17661] ;
  assign n5666 = n5665 & (n3875 | n3881);
  assign n5667 = ~\[18636]  & ~\[18597]  & \[17596]  & ~\[17661] ;
  assign n5668 = ~n3828 & n5667 & (n3829 | n3862);
  assign n5669 = ~\[18636]  & ~\[18597]  & \[17596]  & ~\[17661] ;
  assign n5670 = n5669 & (n3829 | n3862);
  assign n5671 = ~n3796 & ~n3828 & (n5666 | n5670);
  assign n5672 = ~\[18597]  & \[17596]  & ~\[17661] ;
  assign n5673 = ~\[18207]  & ~\[10805]  & ~\[10820] ;
  assign n5674 = ~\[11585]  & ~\[11090]  & ~\[11345]  & ~\[11600] ;
  assign n5675 = ~\[12065]  & ~\[11810]  & ~\[11930]  & ~\[12080] ;
  assign n5676 = ~\[12275]  & ~\[12185]  & ~\[12200]  & ~\[12485] ;
  assign n5677 = n5675 & n5674;
  assign n5678 = n5676 & n5673 & ~\[12695]  & ~\[12935] ;
  assign n5679 = \[17986]  & ~\[17804] ;
  assign n5680 = ~\[17674]  & ~\[17609] ;
  assign n5681 = \[17752]  & ~\[17544]  & \[17713] ;
  assign n5682 = ~ppeaki_6_6_ & ppeaki_4_4_;
  assign n5683 = ~\[17674]  & ~\[17609] ;
  assign n5684 = \[17752]  & ~\[17544]  & ~\[17713] ;
  assign n5685 = ~ppeaki_6_6_ & ~ppeaki_4_4_;
  assign n5686 = ~preset & ((\[18064]  & ~\[18129] ) | (~pirq_0_0_ & (~\[18064]  | ~\[18129] )));
  assign n5687 = n5625 | (\[15545]  & n3698);
  assign n5688 = n5617 | (\[6470]  & n3697) | n5624;
  assign n5689 = n5618 | n5619 | n5620 | n5621;
  assign n5690 = n5622 | n5623 | n5626 | n5689;
  assign n5691 = n5615 | (\[9065]  & n3698);
  assign n5692 = n5607 | (\[5075]  & n3697) | n5614;
  assign n5693 = n5608 | n5609 | n5610 | n5611;
  assign n5694 = n5612 | n5613 | n5616 | n5693;
  assign n5695 = n5605 | n5604;
  assign n5696 = (ppeakp_6_6_ & n3699) | (ppeaka_7_7_ & n3700);
  assign n5697 = (\[12560]  & n3698) | (~ppeaka_6_6_ & n3697);
  assign n5698 = n5599 | (ppeakb_6_6_ & n3701_1) | (~ppeakb_6_6_ & n3697);
  assign n5699 = n5600 | n5601 | n5602 | n5603;
  assign n5700 = n5606 | n5695 | n5696 | n5697;
  assign n5701 = n3756 & (n3964 | n3967_1);
  assign n5702 = n3756 & (n3826 | n3961);
  assign n5703 = n5598 | (\[7655]  & n3756 & n3827_1);
  assign n5704 = n5595 | (\[7640]  & n3756 & n3827_1);
  assign n5705 = ~n3874_1 & ~\[17089]  & ~preset & pdn;
  assign n5706 = ~n5631 & (~n5677 | ~n5678) & n5705;
  assign n5707 = ~n3804 & (n5628 | (~n3955 & n3963));
  assign n5708 = n3857 & (n5706 | n5707);
  assign n5709 = ~preset & (n3783 ? n3960 : ~n3856_1);
  assign n5710 = n5589 | n5588;
  assign n5711 = n5591 | n5580 | n5590;
  assign n5712 = (\[14555]  & n3698) | (\[13700]  & n3697);
  assign n5713 = n5579 | n5581 | n5582 | n5583;
  assign n5714 = n5584 | n5585 | n5586 | n5587;
  assign n5715 = n5592 | n5710 | n5711 | n5712;
  assign n5716 = ppeakb_7_7_ | ppeakb_14_14_ | ppeakb_10_10_ | ppeakb_8_8_;
  assign n5717 = ppeakb_9_9_ | ppeakb_15_15_ | ppeakb_11_11_ | ppeakb_0_0_;
  assign n5718 = ppeakb_1_1_ | ppeakb_12_12_ | ppeakb_2_2_ | ppeakb_3_3_;
  assign n5719 = ppeakb_13_13_ | ppeakb_4_4_ | ppeakb_5_5_ | ppeakb_6_6_;
  assign n5720 = n3756 & (n3821 | n3828);
  assign n5721 = n3963 & (\[17024]  ? ~\[18545]  : ~preset_0_0_);
  assign n5722 = (n3756 & n3808) | (n3955 & n5721);
  assign n5723 = n3756 & (n3957_1 | n3964);
  assign n5724 = n3756 & (n3956 | n3958);
  assign n5725 = n5724 | n5578 | (~preset & ~n3857);
  assign n5726 = n5574 | (\[4850]  & (n5627 | n5628));
  assign n5727 = n5726 | (\[6965]  & n3756 & n3806);
  assign n5728 = n3796 & ~\[18610] ;
  assign n5729 = ~n3797_1 & ~\[18610]  & n3796;
  assign n5730 = n3814 & ~\[18168] ;
  assign n5731 = n3821 & ~\[18493] ;
  assign n5732 = n3876 & ~\[16920] ;
  assign n5733 = n3812_1 & ~\[17297] ;
  assign n5734 = n3815 & ~\[17453] ;
  assign n5735 = n3798 & (n5733 | (~\[16920]  & n3876));
  assign n5736 = n3798 & (n5731 | (n5729 & n5734));
  assign n5737 = n3810 | (~\[17284]  & n3798 & n3802_1);
  assign n5738 = (\[18285]  & ~\[18363] ) | (~\[18311]  & \[18506] );
  assign n5739 = n3813 | n3817_1 | n5550 | n5738;
  assign n5740 = n5551 | (\[10025]  & ~\[18311]  & \[18506] );
  assign n5741 = n5552 | n5553 | n5554 | n5740;
  assign n5742 = n5555 | (\[10310]  & ~\[18311]  & \[18506] );
  assign n5743 = n5556 | n5557 | n5558 | n5742;
  assign n5744 = n5546 | (\[6860]  & ~\[18311]  & \[18506] );
  assign n5745 = n5547 | n5548 | n5549 | n5744;
  assign n5746 = ~n3946 & ~ppeaka_1_1_;
  assign n5747 = ~ppeaka_3_3_ & ~ppeaka_2_2_;
  assign n5748 = ~n3948_1 & ~ppeaka_4_4_;
  assign n5749 = n5540 | (n5748 & (n5541 | n5542));
  assign n5750 = ~ppeaka_6_6_ & ~ppeaka_5_5_;
  assign n5751 = ~ppeaka_9_9_ & ~ppeaka_8_8_;
  assign n5752 = ~n3954 & ~ppeaka_10_10_;
  assign n5753 = ~ppeaka_12_12_ & ~ppeaka_11_11_;
  assign n5754 = ~ppeaka_11_11_ & n3951 & (~ppeaka_10_10_ | ~n3792_1);
  assign n5755 = (~n3951 & (~n3792_1 | (~n5532 & n5754))) | (n3792_1 & ~n5532 & n5754);
  assign n5756 = n5489 | (\[4760]  & ~\[18311]  & \[18506] );
  assign n5757 = n5490 | n5491 | n5492 | n5756;
  assign n5758 = n5494 | (\[6845]  & ~\[18311]  & \[18506] );
  assign n5759 = n5495 | n5496 | n5497 | n5758;
  assign n5760 = ~ppeaka_2_2_ & ~n3893_1 & (~ppeaka_1_1_ | ~n3792_1);
  assign n5761 = ~n5541 & ((n3792_1 & n5760) | (n3900 & (~n3792_1 | n5760)));
  assign n5762 = n5498 | (\[6170]  & ~\[18311]  & \[18506] );
  assign n5763 = n5499 | n5500 | n5501 | n5762;
  assign n5764 = n5502 | (\[8105]  & ~\[18311]  & \[18506] );
  assign n5765 = n5503 | n5504 | n5505 | n5764;
  assign n5766 = n5506 | (\[7475]  & ~\[18311]  & \[18506] );
  assign n5767 = n5507 | n5508 | n5509 | n5766;
  assign n5768 = ~n5749 & ~ppeaka_5_5_ & ~n5539;
  assign n5769 = n5510 | (\[9410]  & ~\[18311]  & \[18506] );
  assign n5770 = n5511 | n5512 | n5513 | n5769;
  assign n5771 = n5514 | (\[8750]  & ~\[18311]  & \[18506] );
  assign n5772 = n5515 | n5516 | n5517 | n5771;
  assign n5773 = n5520 | (\[10040]  & ~\[18311]  & \[18506] );
  assign n5774 = n5521 | n5522 | n5523 | n5773;
  assign n5775 = n5524 | (\[9770]  & ~\[18311]  & \[18506] );
  assign n5776 = n5525 | n5526 | n5527 | n5775;
  assign n5777 = n5528 | (\[10595]  & ~\[18311]  & \[18506] );
  assign n5778 = n5529 | n5530 | n5531 | n5777;
  assign n5779 = n5469 | (\[4775]  & ~\[18311]  & \[18506] );
  assign n5780 = n5470 | n5471 | n5472 | n5779;
  assign n5781 = n5473 | (\[5480]  & ~\[18311]  & \[18506] );
  assign n5782 = n5474 | n5475 | n5476 | n5781;
  assign n5783 = ~ppeaka_13_13_ & ppeaka_14_14_;
  assign n5784 = n3792_1 ? (n5532 & n5783) : (~n3951 & ~n5532);
  assign n5785 = n5464 | (\[8765]  & ~\[18311]  & \[18506] );
  assign n5786 = n5465 | n5466 | n5467 | n5785;
  assign n5787 = ppeaka_15_15_ & ~ppeaka_14_14_;
  assign n5788 = n5787 & n5730 & n3798 & n5729;
  assign n5789 = ~ppeaka_15_15_ & ppeaka_14_14_;
  assign n5790 = n3792_1 ? n5789 : (~n3951 & ~n5532);
  assign n5791 = n3825 | (~\[18025]  & n3798 & n3806);
  assign n5792 = n5455 | n5452 | n5453;
  assign n5793 = n5792 | n5450 | n5451;
  assign n5794 = n5793 | n5454 | n5456;
  assign n5795 = n5448 | n5445 | n5446;
  assign n5796 = n5795 | n5443 | n5444;
  assign n5797 = n5796 | n5447 | n5449;
  assign n5798 = n5441 | n5438 | n5439;
  assign n5799 = n5798 | n5436 | n5437;
  assign n5800 = n5799 | n5440 | n5442;
  assign n5801 = n5434 | n5431 | n5432;
  assign n5802 = n5801 | n5429 | n5430;
  assign n5803 = n5802 | n5433 | n5435;
  assign n5804 = n5427 | n5424 | n5425;
  assign n5805 = n5804 | n5422 | n5423;
  assign n5806 = n5805 | n5426 | n5428;
  assign n5807 = (\[17635]  & ~\[17986] ) | (~\[17037]  & \[18025] );
  assign n5808 = (\[17427]  & ~\[17648] ) | (~\[17999]  & \[18077] );
  assign n5809 = n5808 | n5807;
  assign n5810 = n5809 | (~\[17245]  & n3798 & n3811);
  assign n5811 = n5810 | n5407;
  assign n5812 = n5413 | n5410 | n5411;
  assign n5813 = n5812 | n5408 | n5409;
  assign n5814 = n5813 | n5412 | n5414;
  assign n5815 = n5420 | n5417 | n5418;
  assign n5816 = n5815 | n5415 | n5416;
  assign n5817 = n5816 | n5419 | n5421;
  assign n5818 = (n5811 & n5814) | (n3848 & (ppeaks_0_0_ | n5814));
  assign n5819 = n3803 & n3798 & ppeaka_2_2_ & ~\[16933] ;
  assign n5820 = n3803 & n3798 & ppeaka_3_3_ & ~\[16933] ;
  assign n5821 = n3803 & n3798 & ppeaka_4_4_ & ~\[16933] ;
  assign n5822 = n3803 & n3798 & ppeaka_5_5_ & ~\[16933] ;
  assign n5823 = n3803 & n3798 & ppeaka_6_6_ & ~\[16933] ;
  assign n5824 = n5405 | n5402 | n5403;
  assign n5825 = n5824 | n5400 | n5401;
  assign n5826 = n5825 | n5404 | n5406;
  assign n5827 = n5398 | n5395 | n5396;
  assign n5828 = n5827 | n5393 | n5394;
  assign n5829 = n5828 | n5397 | n5399;
  assign n5830 = n5391 | n5388 | n5389;
  assign n5831 = n5830 | n5386 | n5387;
  assign n5832 = n5831 | n5390 | n5392;
  assign n5833 = n5384 | n5381 | n5382;
  assign n5834 = n5833 | n5379 | n5380;
  assign n5835 = n5834 | n5383 | n5385;
  assign n5836 = n3803 & n3798 & ppeaka_7_7_ & ~\[16933] ;
  assign n5837 = n3803 & n3798 & ppeaka_8_8_ & ~\[16933] ;
  assign n5838 = n3803 & n3798 & ppeaka_9_9_ & ~\[16933] ;
  assign n5839 = n3803 & n3798 & ppeaka_10_10_ & ~\[16933] ;
  assign n5840 = n5376 | n5373 | n5374;
  assign n5841 = n5840 | n5371 | n5372;
  assign n5842 = n5841 | n5375 | n5377;
  assign n5843 = n5369 | n5366 | n5367;
  assign n5844 = n5843 | n5364 | n5365;
  assign n5845 = n5844 | n5368 | n5370;
  assign n5846 = n5362 | n5359 | n5360;
  assign n5847 = n5846 | n5357 | n5358;
  assign n5848 = n5847 | n5361 | n5363;
  assign n5849 = n5355 | n5352 | n5353;
  assign n5850 = n5849 | n5350 | n5351;
  assign n5851 = n5850 | n5354 | n5356;
  assign n5852 = n5348 | n5345 | n5346;
  assign n5853 = n5852 | n5343 | n5344;
  assign n5854 = n5853 | n5347 | n5349;
  assign n5855 = n3803 & n3798 & ppeaka_11_11_ & ~\[16933] ;
  assign n5856 = n3803 & n3798 & ppeaka_12_12_ & ~\[16933] ;
  assign n5857 = n3803 & n3798 & ppeaka_13_13_ & ~\[16933] ;
  assign n5858 = n3803 & n3798 & ppeaka_14_14_ & ~\[16933] ;
  assign n5859 = n5338 | (\[8405]  & n3698);
  assign n5860 = n5330 | (\[4355]  & n3697) | n5337;
  assign n5861 = n5331 | n5332 | n5333 | n5334;
  assign n5862 = n5335 | n5336 | n5339 | n5861;
  assign n5863 = n5328 | n5327;
  assign n5864 = (ppeakp_7_7_ & n3699) | (ppeaka_8_8_ & n3700);
  assign n5865 = (\[12335]  & n3698) | (~ppeaka_7_7_ & n3697);
  assign n5866 = n5322 | (ppeakb_7_7_ & n3701_1) | (~ppeakb_7_7_ & n3697);
  assign n5867 = n5323 | n5324 | n5325 | n5326;
  assign n5868 = n5329 | n5863 | n5864 | n5865;
  assign n5869 = n5321 | (\[9620]  & n3756 & n3827_1);
  assign n5870 = n5318 | (\[9605]  & n3756 & n3827_1);
  assign n5871 = n5312 | n5311;
  assign n5872 = n5314 | n5303 | n5313;
  assign n5873 = (\[14975]  & n3698) | (\[11120]  & n3697);
  assign n5874 = n5302 | n5304 | n5305 | n5306;
  assign n5875 = n5307 | n5308 | n5309 | n5310;
  assign n5876 = n5315 | n5871 | n5872 | n5873;
  assign n5877 = n5299 | (\[5555]  & (n5627 | n5628));
  assign n5878 = n5877 | (\[6290]  & n3756 & n3806);
  assign n5879 = n5265 | (\[14810]  & n3698);
  assign n5880 = n5257 | (\[5090]  & n3697) | n5264;
  assign n5881 = n5258 | n5259 | n5260 | n5261;
  assign n5882 = n5262 | n5263 | n5266 | n5881;
  assign n5883 = n5255 | n5254;
  assign n5884 = (ppeakp_8_8_ & n3699) | (ppeaka_9_9_ & n3700);
  assign n5885 = (\[15695]  & n3698) | (~ppeaka_8_8_ & n3697);
  assign n5886 = n5249 | (ppeakb_8_8_ & n3701_1) | (~ppeakb_8_8_ & n3697);
  assign n5887 = n5250 | n5251 | n5252 | n5253;
  assign n5888 = n5256 | n5883 | n5884 | n5885;
  assign n5889 = n5248 | (\[8945]  & n3756 & n3827_1);
  assign n5890 = n5242 | n5241;
  assign n5891 = n5244 | n5233 | n5243;
  assign n5892 = (\[11375]  & n3697) | (\[6725]  & n3698);
  assign n5893 = n5232 | n5234 | n5235 | n5236;
  assign n5894 = n5237 | n5238 | n5239 | n5240;
  assign n5895 = n5245 | n5890 | n5891 | n5892;
  assign n5896 = n5228 | n5227;
  assign n5897 = n5230 | n5219 | n5229;
  assign n5898 = (\[13745]  & n3698) | (\[9275]  & n3697);
  assign n5899 = n5218 | n5220 | n5221 | n5222;
  assign n5900 = n5223 | n5224 | n5225 | n5226;
  assign n5901 = n5231 | n5896 | n5897 | n5898;
  assign n5902 = n5215 | (\[8855]  & (n5627 | n5628));
  assign n5903 = n5902 | (\[11210]  & n3756 & n3806);
  assign n5904 = n5180 | (\[15890]  & n3698);
  assign n5905 = n5172 | (\[4370]  & n3697) | n5179;
  assign n5906 = n5173 | n5174 | n5175 | n5176;
  assign n5907 = n5177 | n5178 | n5181 | n5906;
  assign n5908 = n5170 | (\[7130]  & n3698);
  assign n5909 = n5162 | (\[5780]  & n3697) | n5169;
  assign n5910 = n5163 | n5164 | n5165 | n5166;
  assign n5911 = n5167 | n5168 | n5171 | n5910;
  assign n5912 = n5161 | (\[5630]  & n3756 & n3827_1);
  assign n5913 = n5155 | n5154;
  assign n5914 = n5157 | n5146 | n5156;
  assign n5915 = (\[15320]  & n3697) | (\[7355]  & n3698);
  assign n5916 = n5145 | n5147 | n5148 | n5149;
  assign n5917 = n5150 | n5151 | n5152 | n5153;
  assign n5918 = n5158 | n5913 | n5914 | n5915;
  assign n5919 = n5141 | n5140;
  assign n5920 = n5143 | n5132 | n5142;
  assign n5921 = (\[14135]  & n3698) | (\[8615]  & n3697);
  assign n5922 = n5131 | n5133 | n5134 | n5135;
  assign n5923 = n5136 | n5137 | n5138 | n5139;
  assign n5924 = n5144 | n5919 | n5920 | n5921;
  assign n5925 = n5128 | (\[9530]  & (n5627 | n5628));
  assign n5926 = n5925 | (\[10955]  & n3756 & n3806);
  assign n5927 = n5100 | (\[11240]  & n3756 & n3827_1);
  assign n5928 = n5094 | n5093;
  assign n5929 = n5096 | n5085 | n5095;
  assign n5930 = (\[5360]  & n3698) | (\[4640]  & n3697);
  assign n5931 = n5084 | n5086 | n5087 | n5088;
  assign n5932 = n5089 | n5090 | n5091 | n5092;
  assign n5933 = n5097 | n5928 | n5929 | n5930;
  assign n5934 = n5080 | n5079;
  assign n5935 = n5082 | n5071 | n5081;
  assign n5936 = (\[16055]  & n3698) | (\[4625]  & n3697);
  assign n5937 = n5070 | n5072 | n5073 | n5074;
  assign n5938 = n5075 | n5076 | n5077 | n5078;
  assign n5939 = n5083 | n5934 | n5935 | n5936;
  assign n5940 = n5067 | (\[7565]  & (n5627 | n5628));
  assign n5941 = n5940 | (\[11195]  & n3756 & n3806);
  assign n5942 = n5036 | (\[10430]  & n3756 & n3827_1);
  assign n5943 = n5030 | n5029;
  assign n5944 = n5032 | n5021 | n5031;
  assign n5945 = (\[6050]  & n3698) | (\[5345]  & n3697);
  assign n5946 = n5020 | n5022 | n5023 | n5024;
  assign n5947 = n5025 | n5026 | n5027 | n5028;
  assign n5948 = n5033 | n5943 | n5944 | n5945;
  assign n5949 = n5017 | (\[9815]  & (n5627 | n5628));
  assign n5950 = n5949 | (\[8900]  & n3756 & n3806);
  assign n5951 = n5013 | (\[8195]  & (n5627 | n5628));
  assign n5952 = n5951 | (\[10940]  & n3756 & n3806);
  assign n5953 = n4982 | (\[10715]  & n3756 & n3827_1);
  assign n5954 = n4976 | n4975;
  assign n5955 = n4978 | n4967 | n4977;
  assign n5956 = (\[15350]  & n3698) | (\[6020]  & n3697);
  assign n5957 = n4966 | n4968 | n4969 | n4970;
  assign n5958 = n4971 | n4972 | n4973 | n4974;
  assign n5959 = n4979 | n5954 | n5955 | n5956;
  assign n5960 = n4963 | (\[10655]  & (n5627 | n5628));
  assign n5961 = n5960 | (\[5600]  & n3756 & n3806);
  assign n5962 = n4959 | (\[6260]  & (n5627 | n5628));
  assign n5963 = n5962 | (\[6950]  & n3756 & n3806);
  assign n5964 = n4929 | n4928;
  assign n5965 = n4931 | n4920 | n4930;
  assign n5966 = (\[6710]  & n3697) | (\[4655]  & n3698);
  assign n5967 = n4919 | n4921 | n4922 | n4923;
  assign n5968 = n4924 | n4925 | n4926 | n4927;
  assign n5969 = n4932 | n5964 | n5965 | n5966;
  assign n5970 = n4915 | n4914;
  assign n5971 = n4917 | n4906 | n4916;
  assign n5972 = (\[15710]  & n3698) | (\[6695]  & n3697);
  assign n5973 = n4905 | n4907 | n4908 | n4909;
  assign n5974 = n4910 | n4911 | n4912 | n4913;
  assign n5975 = n4918 | n5970 | n5971 | n5972;
  assign n5976 = n4902 | (\[10370]  & (n5627 | n5628));
  assign n5977 = n5976 | (\[4895]  & n3756 & n3806);
  assign n5978 = n4898 | (\[6935]  & (n5627 | n5628));
  assign n5979 = n5978 | (\[6275]  & n3756 & n3806);
  assign n5980 = n4769 | (\[13250]  & n3698);
  assign n5981 = n4761 | (\[13235]  & n3697) | n4768;
  assign n5982 = n4762 | n4763 | n4764 | n4765;
  assign n5983 = n4766 | n4767 | n4770 | n5982;
  assign n5984 = n4754 | (\[7880]  & n3756 & n3812_1);
  assign n5985 = n5984 | n4751;
  assign n5986 = n4744 | n4745 | n4746 | n4747;
  assign n5987 = n4748 | n4749 | n4750 | n4752;
  assign n5988 = n4731 | (\[6620]  & n3756 & n3812_1);
  assign n5989 = n5988 | n4728;
  assign n5990 = n4721 | n4722 | n4723 | n4724;
  assign n5991 = n4725 | n4726 | n4727 | n4729;
  assign n5992 = n4661 | (\[5795]  & n3698);
  assign n5993 = n4653 | (\[14360]  & n3697) | n4660;
  assign n5994 = n4654 | n4655 | n4656 | n4657;
  assign n5995 = n4658 | n4659 | n4662 | n5994;
  assign n5996 = n4651 | n4650;
  assign n5997 = (ppeakp_9_9_ & n3699) | (ppeaka_10_10_ & n3700);
  assign n5998 = (\[16040]  & n3698) | (~ppeaka_9_9_ & n3697);
  assign n5999 = n4645 | (ppeakb_9_9_ & n3701_1) | (~ppeakb_9_9_ & n3697);
  assign n6000 = n4646 | n4647 | n4648 | n4649;
  assign n6001 = n4652 | n5996 | n5997 | n5998;
  assign n6002 = n4623 | (\[6485]  & n3698);
  assign n6003 = n4615 | (\[13955]  & n3697) | n4622;
  assign n6004 = n4616 | n4617 | n4618 | n4619;
  assign n6005 = n4620 | n4621 | n4624 | n6004;
  assign n6006 = n4614 | (\[9890]  & n3756 & n3827_1);
  assign n6007 = n4609 | (\[10085]  & (n5627 | n5628));
  assign n6008 = n6007 | (\[9575]  & n3756 & n3806);
  assign n6009 = n4585 | n4584_1;
  assign n6010 = (ppeakp_11_11_ & n3699) | (ppeaka_12_12_ & n3700);
  assign n6011 = (\[15335]  & n3698) | (~ppeakb_11_11_ & n3697);
  assign n6012 = n4579_1 | n4578 | (~ppeaka_11_11_ & n3697);
  assign n6013 = n4580 | n4581 | n4582 | n4583;
  assign n6014 = n4586 | n6009 | n6010 | n6011;
  assign n6015 = n4575 | n4565_1 | n4566;
  assign n6016 = n4567 | n4568 | n4569 | n4570_1;
  assign n6017 = n4564 | n4571 | n4572 | n4576;
  assign n6018 = n4573 | n4574_1 | n6015 | n6017;
  assign n6019 = n4561_1 | (\[8840]  & (n5627 | n5628));
  assign n6020 = n6019 | (\[11660]  & n3756 & n3806);
  assign n6021 = n4538 | (\[14915]  & n3756 & n3812_1);
  assign n6022 = n6021 | n4535;
  assign n6023 = n4528_1 | n4529 | n4530 | n4531;
  assign n6024 = n4532 | n4533_1 | n4534 | n4536;
  assign n6025 = n4525 | n4515 | n4516;
  assign n6026 = n4517 | n4518_1 | n4519 | n4520;
  assign n6027 = n4514_1 | n4521 | n4522 | n4526;
  assign n6028 = n4523_1 | n4524 | n6025 | n6027;
  assign n6029 = n4511 | n4501 | n4502;
  assign n6030 = n4503 | n4504_1 | n4505 | n4506;
  assign n6031 = n4500 | n4507 | n4508 | n4512;
  assign n6032 = n4509_1 | n4510 | n6029 | n6031;
  assign n6033 = n4497 | (\[9515]  & (n5627 | n5628));
  assign n6034 = n6033 | (\[11435]  & n3756 & n3806);
  assign n6035 = n4471 | (\[13010]  & n3756 & n3812_1);
  assign n6036 = n6035 | n4468;
  assign n6037 = n4461 | n4462_1 | n4463 | n4464;
  assign n6038 = n4465 | n4466_1 | n4467 | n4469;
  assign n6039 = n4459 | n4458;
  assign n6040 = (ppeakp_13_13_ & n3699) | (ppeaka_14_14_ & n3700);
  assign n6041 = (\[14540]  & n3698) | (~ppeakb_13_13_ & n3697);
  assign n6042 = n4453 | n4452_1 | (~ppeaka_13_13_ & n3697);
  assign n6043 = n4454 | n4455 | n4456 | n4457_1;
  assign n6044 = n4460 | n6039 | n6040 | n6041;
  assign n6045 = n4449 | n4439 | n4440;
  assign n6046 = n4441 | n4442_1 | n4443 | n4444;
  assign n6047 = n4438 | n4445 | n4446 | n4450;
  assign n6048 = n4447_1 | n4448 | n6045 | n6047;
  assign n6049 = n4437_1 | (\[9875]  & n3756 & n3827_1);
  assign n6050 = n4431 | n4430;
  assign n6051 = n4433 | n4422_1 | n4432_1;
  assign n6052 = (\[13040]  & n3698) | (\[7970]  & n3697);
  assign n6053 = n4421 | n4423 | n4424 | n4425;
  assign n6054 = n4426 | n4427_1 | n4428 | n4429;
  assign n6055 = n4434 | n6050 | n6051 | n6052;
  assign n6056 = n4418 | (\[7580]  & (n5627 | n5628));
  assign n6057 = n6056 | (\[11675]  & n3756 & n3806);
  assign n6058 = n4397_1 | (\[16010]  & n3756 & n3812_1);
  assign n6059 = n6058 | n4394;
  assign n6060 = n4387_1 | n4388 | n4389 | n4390;
  assign n6061 = n4391 | n4392_1 | n4393 | n4395;
  assign n6062 = n4385 | n4384;
  assign n6063 = (ppeaka_13_13_ & n3700) | (ppeakp_12_12_ & n3699);
  assign n6064 = (\[14120]  & n3698) | (~ppeaka_12_12_ & n3697);
  assign n6065 = n4379 | (ppeakb_12_12_ & n3701_1) | (~ppeakb_12_12_ & n3697);
  assign n6066 = n4380 | n4381 | n4382 | n4383_1;
  assign n6067 = n4386 | n6062 | n6063 | n6064;
  assign n6068 = n4376 | n4366 | n4367;
  assign n6069 = n4368_1 | n4369 | n4370 | n4371;
  assign n6070 = n4365 | n4372 | n4373_1 | n4377;
  assign n6071 = n4374 | n4375 | n6068 | n6070;
  assign n6072 = n4364 | (\[10730]  & n3756 & n3827_1);
  assign n6073 = n4358_1 | n4357;
  assign n6074 = n4360 | n4349 | n4359;
  assign n6075 = (\[13385]  & n3698) | (\[7340]  & n3697);
  assign n6076 = n4348_1 | n4350 | n4351 | n4352;
  assign n6077 = n4353_1 | n4354 | n4355 | n4356;
  assign n6078 = n4361 | n6073 | n6074 | n6075;
  assign n6079 = n4345 | (\[8210]  & (n5627 | n5628));
  assign n6080 = n6079 | (\[11450]  & n3756 & n3806);
  assign n6081 = n4326 | (\[13685]  & n3756 & n3812_1);
  assign n6082 = n6081 | n4323;
  assign n6083 = n4316 | n4317 | n4318 | n4319_1;
  assign n6084 = n4320 | n4321 | n4322 | n4324_1;
  assign n6085 = n4303 | n4304_1 | n4305 | n4306;
  assign n6086 = n4307 | n4308 | n4310 | n4314_1;
  assign n6087 = n4309_1 | n4311 | n4312 | n4313;
  assign n6088 = n4300_1 | n4290_1 | n4291;
  assign n6089 = n4292 | n4293 | n4294 | n4295_1;
  assign n6090 = n4289 | n4296 | n4297 | n4301;
  assign n6091 = n4298 | n4299 | n6088 | n6090;
  assign n6092 = n4288 | (\[10445]  & n3756 & n3827_1);
  assign n6093 = n4285_1 | (\[8930]  & n3756 & n3827_1);
  assign n6094 = n4279 | n4278;
  assign n6095 = n4281 | n4270_1 | n4280_1;
  assign n6096 = (\[13025]  & n3698) | (\[5330]  & n3697);
  assign n6097 = n4269 | n4271 | n4272 | n4273;
  assign n6098 = n4274 | n4275_1 | n4276 | n4277;
  assign n6099 = n4282 | n6094 | n6095 | n6096;
  assign n6100 = n4254 | (\[6500]  & n3698);
  assign n6101 = n4246 | (\[7115]  & n3697) | n4253;
  assign n6102 = n4247_1 | n4248 | n4249 | n4250;
  assign n6103 = n4251_1 | n4252 | n4255 | n6102;
  assign n6104 = n4244 | n4243;
  assign n6105 = (ppeakp_14_14_ & n3699) | (ppeaka_15_15_ & n3700);
  assign n6106 = (\[13370]  & n3698) | (~ppeaka_14_14_ & n3697);
  assign n6107 = n4238 | (ppeakb_14_14_ & n3701_1) | (~ppeakb_14_14_ & n3697);
  assign n6108 = n4239 | n4240 | n4241 | n4242_1;
  assign n6109 = n4245 | n6104 | n6105 | n6106;
  assign n6110 = n4235 | n4225 | n4226;
  assign n6111 = n4227_1 | n4228 | n4229 | n4230;
  assign n6112 = n4224 | n4231 | n4232_1 | n4236;
  assign n6113 = n4233 | n4234 | n6110 | n6112;
  assign n6114 = n4223_1 | (\[8285]  & n3756 & n3827_1);
  assign n6115 = n4220 | (\[10145]  & n3756 & n3827_1);
  assign n6116 = n4214 | n4213_1;
  assign n6117 = n4216 | n4205 | n4215;
  assign n6118 = (\[12800]  & n3698) | (\[6035]  & n3697);
  assign n6119 = n4204 | n4206 | n4207 | n4208_1;
  assign n6120 = n4209 | n4210 | n4211 | n4212;
  assign n6121 = n4217 | n6116 | n6117 | n6118;
  assign n6122 = (\[17999]  & ~\[18220] ) | (~\[17791]  & n3788);
  assign n6123 = (\[17180]  & ~\[17232] ) | (~\[17050]  & \[17115] );
  assign n6124 = (\[17206]  & ~\[17271] ) | (\[16933]  & ~\[17388] );
  assign n6125 = (\[18311]  & ~\[18389] ) | (~\[17414]  & \[17843] );
  assign n6126 = n6125 | n6124;
  assign n6127 = n3789 | n3794 | n3879 | n6123;
  assign n6128 = n3816 | n6122 | n6126 | n6127;
  assign n6129 = n6128 | (~\[17167]  & n3798 & n3819);
  assign n6130 = n3858 | n3813 | n3817_1;
  assign n6131 = n3792_1 | n5735 | n5736 | n6129;
  assign n6132 = n4141 | (~preset & \[17284]  & ~\[18376] );
  assign n6133 = n6132 | (~preset & n3798 & n5732);
  assign n6134 = ~preset & n3798 & (n5731 | n5733);
  assign n6135 = n4182 | n4181;
  assign n6136 = n4183 | (ppeakb_8_8_ & n3777_1);
  assign n6137 = (\[13460]  & n3775) | (\[7595]  & n3776);
  assign n6138 = (\[11420]  & n3773) | (\[6410]  & n3774);
  assign n6139 = n4177 | n4178 | n4179_1 | n4180;
  assign n6140 = n4184_1 | n4185 | n6135 | n6136;
  assign n6141 = n4186 | n6137 | n6138 | n6139;
  assign n6142 = n4176 | (~preset & ppeakb_7_7_ & n3859);
  assign n6143 = ~\[17388]  & ~preset;
  assign n6144 = n4170 | n4169_1;
  assign n6145 = n4171 | (ppeakb_9_9_ & n3777_1);
  assign n6146 = (\[13820]  & n3775) | (\[10685]  & n3776);
  assign n6147 = (\[11645]  & n3773) | (\[5720]  & n3774);
  assign n6148 = n4165_1 | n4166 | n4167 | n4168;
  assign n6149 = n4172 | n4173 | n6144 | n6145;
  assign n6150 = n4174_1 | n6146 | n6147 | n6148;
  assign n6151 = n4164 | (~preset & ppeakb_8_8_ & n3859);
  assign n6152 = n4162 | (~preset & ppeakb_5_5_ & n3859);
  assign n6153 = n4160_1 | (~preset & ppeakb_6_6_ & n3859);
  assign n6154 = n4158 | (~preset & ppeakb_15_15_ & n3859);
  assign n6155 = ~\[17050]  & ~preset;
  assign n6156 = n4156 | (~preset & ppeakb_3_3_ & n3859);
  assign n6157 = ~\[17232]  & ~preset;
  assign n6158 = n4154 | (~preset & ppeakb_4_4_ & n3859);
  assign n6159 = ~\[17271]  & ~preset;
  assign n6160 = n4152 | (~preset & ppeakb_1_1_ & n3859);
  assign n6161 = ~\[18376]  & ~preset;
  assign n6162 = n4150_1 | (~preset & ppeakb_2_2_ & n3859);
  assign n6163 = n4144 | n4143;
  assign n6164 = n4145 | (ppeakb_11_11_ & n3777_1);
  assign n6165 = (\[13115]  & n3775) | (\[10115]  & n3776);
  assign n6166 = (\[16100]  & n3773) | (\[4295]  & n3774);
  assign n6167 = n4139 | n4140 | n4141_1 | n4142;
  assign n6168 = n4146_1 | n4147 | n6163 | n6164;
  assign n6169 = n4148 | n6165 | n6166 | n6167;
  assign n6170 = n4134 | n4133;
  assign n6171 = n4135 | (ppeakb_10_10_ & n3777_1);
  assign n6172 = (\[12860]  & n3775) | (\[10400]  & n3776);
  assign n6173 = (\[10925]  & n3773) | (\[5015]  & n3774);
  assign n6174 = n4129 | n4130 | n4131_1 | n4132;
  assign n6175 = n4136_1 | n4137 | n6170 | n6171;
  assign n6176 = n4138 | n6172 | n6173 | n6174;
  assign n6177 = n4128 | (~preset & ppeakb_13_13_ & n3859);
  assign n6178 = n4121_1 | n4120;
  assign n6179 = n4122 | (ppeakb_13_13_ & n3777_1);
  assign n6180 = (\[12620]  & n3775) | (\[8885]  & n3776);
  assign n6181 = (\[15500]  & n3774) | (\[13805]  & n3773);
  assign n6182 = n4116_1 | n4117 | n4118 | n4119;
  assign n6183 = n4123 | n4124 | n6178 | n6179;
  assign n6184 = n4125 | n6180 | n6181 | n6182;
  assign n6185 = ~n3883_1 | (~ppeaki_13_13_ & ~ppeaki_12_12_);
  assign n6186 = ~n3883_1 | (~ppeaki_15_15_ & ~ppeaki_14_14_);
  assign n6187 = n6185 & (~n3883_1 | (~ppeaki_15_15_ & ~ppeaki_14_14_));
  assign n6188 = ~n3759 & ~n3755 & ~n3758_1 & ~n3765;
  assign n6189 = ~n3770 & ~n3766 & ~n3768_1 & ~n3772_1;
  assign n6190 = n6188 & n6185 & n6186;
  assign n6191 = n6189 & (\[18636]  | (~n3798 & n5672));
  assign n6192 = \[17986]  & \[17596] ;
  assign n6193 = n4115 | \[17804]  | (\[17986]  & \[18597] );
  assign n6194 = ~\[18597]  & ~preset & \[17596] ;
  assign n6195 = n3790 & ~preset & ~\[17596] ;
  assign n6196 = n4109 | n4108;
  assign n6197 = n4110 | (ppeakb_12_12_ & n3777_1);
  assign n6198 = (\[12395]  & n3775) | (\[9845]  & n3776);
  assign n6199 = (\[15845]  & n3774) | (\[15755]  & n3773);
  assign n6200 = n4104 | n4105 | n4106_1 | n4107;
  assign n6201 = n4111_1 | n4112 | n6196 | n6197;
  assign n6202 = n4113 | n6198 | n6199 | n6200;
  assign n6203 = n4099 | n4098;
  assign n6204 = n4100 | (ppeakb_15_15_ & n3777_1);
  assign n6205 = (\[15050]  & n3775) | (\[4880]  & n3776);
  assign n6206 = (\[14615]  & n3773) | (\[13550]  & n3774);
  assign n6207 = n4094 | n4095 | n4096_1 | n4097;
  assign n6208 = n4101_1 | n4102 | n6203 | n6204;
  assign n6209 = n4103 | n6205 | n6206 | n6207;
  assign n6210 = n4089 | n4088;
  assign n6211 = n4090 | (ppeakb_14_14_ & n3777_1);
  assign n6212 = (\[15410]  & n3775) | (\[9560]  & n3776);
  assign n6213 = (\[15140]  & n3774) | (\[13445]  & n3773);
  assign n6214 = n4084 | n4085 | n4086_1 | n4087;
  assign n6215 = n4091_1 | n4092 | n6210 | n6211;
  assign n6216 = n4093 | n6212 | n6213 | n6214;
  assign n6217 = n4083 | (~preset & ppeakb_9_9_ & n3859);
  assign n6218 = n4081_1 | (~preset & ppeakb_14_14_ & n3859);
  assign n6219 = (\[17180]  & ~\[17232] ) | (~\[17050]  & \[17115] );
  assign n6220 = (\[17206]  & ~\[17271] ) | (\[17232]  & ~\[18441] );
  assign n6221 = (\[17583]  & ~\[18077] ) | (~\[17427]  & \[17518] );
  assign n6222 = (\[17050]  & ~\[17219] ) | (\[17271]  & ~\[17349] );
  assign n6223 = n3789 | n3879 | n6219 | n6220;
  assign n6224 = n6223 | n6221 | n6222;
  assign n6225 = n3789 & ~preset;
  assign n6226 = pwr_0_0_ & ~preset;
  assign n6227 = (~n3858 & ~n6224 & n6226) | (n6225 & (n3858 | n6224));
  assign n6228 = ~preset & (n3858 | (n3781 & n6224));
  assign n6229 = (n4011 | n4081) & (n3858 | n6224);
  assign n6230 = (\[16933]  & ~\[17388] ) | (~\[17414]  & \[17843] );
  assign n6231 = (\[18311]  & ~\[18389] ) | (\[18363]  & ~\[18415] );
  assign n6232 = (\[17791]  & ~\[17843] ) | (\[17453]  & ~\[18246] );
  assign n6233 = (\[17102]  & ~\[17154] ) | (\[17167]  & ~\[17362] );
  assign n6234 = (\[17414]  & ~\[17505] ) | (~\[17310]  & \[17388] );
  assign n6235 = (~\[18142]  & \[18220] ) | (~\[18311]  & \[18506] );
  assign n6236 = (\[17570]  & ~\[17635] ) | (\[18285]  & ~\[18363] );
  assign n6237 = (\[18415]  & ~\[18480] ) | (~\[18428]  & \[18493] );
  assign n6238 = (~\[18298]  & \[18376] ) | (~\[16985]  & \[18389] );
  assign n6239 = (\[16920]  & ~\[16972] ) | (\[17297]  & ~\[17375] );
  assign n6240 = n6239 | n3879 | n6230;
  assign n6241 = n6231 | n6232 | n6233 | n6234;
  assign n6242 = n6235 | n6236 | n6237 | n6238;
  assign n6243 = n6242 | n6240 | n6241;
  assign n6244 = n6243 | n3816 | n6122;
  assign n6245 = n6244 | (~\[17167]  & n3798 & n3819);
  assign n6246 = n3792_1 | n3813 | n3817_1 | n6245;
  assign n6247 = ~preset & (n3816 | n6122);
  assign n6248 = prd_0_0_ & ~preset;
  assign n6249 = (~n3878_1 & ~n6246 & n6248) | (n6247 & (n3878_1 | n6246));
  assign n6250 = (n3706_1 | n3709) & (n3878_1 | n6246);
  assign n6251 = (n4518 | n3791) & (n3878_1 | n6246);
  assign n6252 = (n4150 | n4509) & (n3878_1 | n6246);
  assign n6253 = (n4031 | n4056) & (n3878_1 | n6246);
  assign n6254 = n6253 | n6249 | n6250;
  assign n6255 = n4078 | (~preset & ppeakb_10_10_ & n3859);
  assign n6256 = n4076_1 | (~preset & ppeakb_12_12_ & n3859);
  assign n6257 = \[18129]  & ~preset;
  assign n6258 = n4065 | (~preset & ppeakb_11_11_ & n3859);
  assign n6259 = n4057 | n4056_1;
  assign n6260 = (\[10670]  & n3776) | (ppeakb_0_0_ & n3777_1);
  assign n6261 = (\[12605]  & n3775) | (\[4310]  & n3774);
  assign n6262 = n4051_1 | (\[11630]  & n3773) | n4061_1;
  assign n6263 = n4052 | n4053 | n4054 | n4055;
  assign n6264 = n4058 | n4059 | n6259 | n6260;
  assign n6265 = n4060 | n6261 | n6262 | n6263;
  assign n6266 = ~\[18415]  & ~preset;
  assign n6267 = n4047 | n4043;
  assign n6268 = (\[9830]  & n3776) | (ppeakb_1_1_ & n3777_1);
  assign n6269 = (\[12380]  & n3775) | (\[5030]  & n3774);
  assign n6270 = n4037 | (\[9485]  & n3773) | n4038;
  assign n6271 = n4039 | n4040 | n4041_1 | n4042;
  assign n6272 = n4044 | n4045 | n6267 | n6268;
  assign n6273 = n4046_1 | n6269 | n6270 | n6271;
  assign n6274 = n4036_1 | (~preset & ppeakb_0_0_ & n3859);
  assign n6275 = n4030 | n4029;
  assign n6276 = n4031_1 | (ppeakb_2_2_ & n3777_1);
  assign n6277 = (\[13100]  & n3775) | (\[10100]  & n3776);
  assign n6278 = (\[15515]  & n3774) | (\[7535]  & n3773);
  assign n6279 = n4025 | n4026_1 | n4027 | n4028;
  assign n6280 = n4032 | n4033 | n6275 | n6276;
  assign n6281 = n4034 | n6277 | n6278 | n6279;
  assign n6282 = n4020 | n4019;
  assign n6283 = n4021_1 | (ppeakb_3_3_ & n3777_1);
  assign n6284 = (\[12845]  & n3775) | (\[5570]  & n3776);
  assign n6285 = (\[15860]  & n3774) | (\[8165]  & n3773);
  assign n6286 = n4015 | n4016_1 | n4017 | n4018;
  assign n6287 = n4022 | n4023 | n6282 | n6283;
  assign n6288 = n4024 | n6284 | n6285 | n6286;
  assign n6289 = \[17700]  & ~preset & ~pdn;
  assign n6290 = n4008 | n4007;
  assign n6291 = n4009 | (ppeakb_4_4_ & n3777_1);
  assign n6292 = (\[15035]  & n3775) | (\[4865]  & n3776);
  assign n6293 = (\[14765]  & n3774) | (\[6230]  & n3773);
  assign n6294 = n4003 | n4004 | n4005 | n4006_1;
  assign n6295 = n4010 | n4011_1 | n6290 | n6291;
  assign n6296 = n4012 | n6292 | n6293 | n6294;
  assign n6297 = n3998 | n3997;
  assign n6298 = n3999 | (ppeakb_5_5_ & n3777_1);
  assign n6299 = (\[15395]  & n3775) | (\[9545]  & n3776);
  assign n6300 = (\[8330]  & n3774) | (\[6905]  & n3773);
  assign n6301 = n3993 | n3994 | n3995 | n3996_1;
  assign n6302 = n4000 | n4001_1 | n6297 | n6298;
  assign n6303 = n4002 | n6299 | n6300 | n6301;
  assign n6304 = n3988 | n3987;
  assign n6305 = n3989 | (ppeakb_6_6_ & n3777_1);
  assign n6306 = (\[14210]  & n3775) | (\[8870]  & n3776);
  assign n6307 = (\[7685]  & n3774) | (\[4835]  & n3773);
  assign n6308 = n3983 | n3984 | n3985 | n3986_1;
  assign n6309 = n3990 | n3991_1 | n6304 | n6305;
  assign n6310 = n3992 | n6306 | n6307 | n6308;
  assign n6311 = \[17596]  & ~preset & ~pdn;
  assign n6312 = n3798 & ~preset & n3796;
  assign n6313 = n3798 & n3797_1 & ~preset & n3796;
  assign n6314 = n3798 & n3796 & ~preset & \[18168] ;
  assign n6315 = n3798 & n3796 & ~preset & \[17453] ;
  assign n6316 = ~n3783 & (n6313 | n6314);
  assign n6317 = ~n3783 & (n6315 | (~n3787_1 & n6312));
  assign n6318 = n3976_1 | n3975;
  assign n6319 = n3977 | (ppeakb_7_7_ & n3777_1);
  assign n6320 = (\[14630]  & n3775) | (\[8225]  & n3776);
  assign n6321 = (\[7055]  & n3774) | (\[5540]  & n3773);
  assign n6322 = n3971 | n3972_1 | n3973 | n3974;
  assign n6323 = n3978 | n3979 | n6318 | n6319;
  assign n6324 = n3980 | n6320 | n6321 | n6322;
  assign n6325 = ~preset & n3798 & (\[18493]  | n3811);
  assign n6326 = ~preset & n3798 & (\[18389]  | \[18415] );
  assign n6327 = ~preset & n3798 & (\[17388]  | \[18376] );
  assign n6328 = ~preset & n3798 & (\[17271]  | \[17297] );
  assign n6329 = ~preset & n3798 & (\[17167]  | \[17232] );
  assign n6330 = ~preset & n3798 & (\[17050]  | \[17102] );
  assign n6331 = n6330 | n3969 | n6325;
  assign n6332 = n6326 | n6327 | n6328 | n6329;
  always @ (posedge pclk) begin
    ndout <= n273;
    ppeakb_12_12_ <= n278;
    ppeakb_1_1_ <= n282;
    ppeaka_6_6_ <= n286;
    \[4295]  <= n290;
    \[4310]  <= n295;
    ppeaks_5_5_ <= n300;
    ppeakp_10_10_ <= n304;
    \[4355]  <= n308;
    \[4370]  <= n313;
    \[4385]  <= n318;
    \[4400]  <= n323;
    \[4415]  <= n328;
    \[4430]  <= n333;
    \[4445]  <= n338;
    \[4460]  <= n343;
    \[4475]  <= n348;
    \[4490]  <= n353;
    \[4505]  <= n358;
    \[4520]  <= n363;
    \[4535]  <= n368;
    \[4550]  <= n373;
    \[4565]  <= n378;
    \[4580]  <= n383;
    \[4595]  <= n388;
    \[4610]  <= n393;
    \[4625]  <= n398;
    \[4640]  <= n403;
    \[4655]  <= n408;
    \[4670]  <= n413;
    \[4700]  <= n418;
    \[4715]  <= n423;
    \[4730]  <= n428;
    \[4745]  <= n433;
    \[4760]  <= n438;
    \[4775]  <= n443;
    \[4790]  <= n448;
    \[4805]  <= n453;
    \[4820]  <= n458;
    \[4835]  <= n463;
    \[4850]  <= n468;
    \[4865]  <= n473;
    \[4880]  <= n478;
    \[4895]  <= n483;
    \[4910]  <= n488;
    \[4925]  <= n493;
    \[4940]  <= n498;
    \[4955]  <= n503;
    \[4970]  <= n508;
    ppeakb_0_0_ <= n513;
    ppeaka_7_7_ <= n517;
    \[5015]  <= n521;
    \[5030]  <= n526;
    ppeaks_4_4_ <= n531;
    ppeakp_11_11_ <= n535;
    \[5075]  <= n539;
    \[5090]  <= n544;
    \[5105]  <= n549;
    \[5120]  <= n554;
    \[5135]  <= n559;
    \[5150]  <= n564;
    \[5165]  <= n569;
    \[5180]  <= n574;
    \[5195]  <= n579;
    \[5210]  <= n584;
    \[5225]  <= n589;
    \[5240]  <= n594;
    \[5255]  <= n599;
    \[5270]  <= n604;
    \[5285]  <= n609;
    \[5300]  <= n614;
    \[5315]  <= n619;
    \[5330]  <= n624;
    \[5345]  <= n629;
    \[5360]  <= n634;
    \[5375]  <= n639;
    \[5390]  <= n644;
    \[5405]  <= n649;
    \[5420]  <= n654;
    \[5435]  <= n659;
    \[5450]  <= n664;
    \[5465]  <= n669;
    \[5480]  <= n674;
    \[5495]  <= n679;
    \[5510]  <= n684;
    \[5525]  <= n689;
    \[5540]  <= n694;
    \[5555]  <= n699;
    \[5570]  <= n704;
    \[5600]  <= n709;
    \[5615]  <= n714;
    \[5630]  <= n719;
    \[5645]  <= n724;
    \[5660]  <= n729;
    \[5675]  <= n734;
    ppeakb_10_10_ <= n739;
    ppeaka_8_8_ <= n743;
    \[5720]  <= n747;
    ppeaks_14_14_ <= n752;
    ppeaks_7_7_ <= n756;
    ppeakp_12_12_ <= n760;
    \[5780]  <= n764;
    \[5795]  <= n769;
    \[5810]  <= n774;
    \[5825]  <= n779;
    \[5840]  <= n784;
    \[5855]  <= n789;
    \[5870]  <= n794;
    \[5885]  <= n799;
    \[5900]  <= n804;
    \[5915]  <= n809;
    \[5930]  <= n814;
    \[5945]  <= n819;
    \[5960]  <= n824;
    \[5975]  <= n829;
    \[5990]  <= n834;
    \[6005]  <= n839;
    \[6020]  <= n844;
    \[6035]  <= n849;
    \[6050]  <= n854;
    \[6065]  <= n859;
    \[6080]  <= n864;
    \[6095]  <= n869;
    \[6110]  <= n874;
    \[6125]  <= n879;
    \[6140]  <= n884;
    \[6155]  <= n889;
    \[6170]  <= n894;
    \[6185]  <= n899;
    \[6200]  <= n904;
    \[6215]  <= n909;
    \[6230]  <= n914;
    \[6245]  <= n919;
    \[6260]  <= n924;
    \[6275]  <= n929;
    \[6290]  <= n934;
    \[6305]  <= n939;
    \[6320]  <= n944;
    \[6335]  <= n949;
    \[6350]  <= n954;
    \[6365]  <= n959;
    ppeakb_11_11_ <= n964;
    ppeakb_2_2_ <= n968;
    \[6410]  <= n972;
    ppeaks_15_15_ <= n977;
    ppeaks_6_6_ <= n981;
    ppeakp_13_13_ <= n985;
    \[6470]  <= n989;
    \[6485]  <= n994;
    \[6500]  <= n999;
    \[6515]  <= n1004;
    \[6530]  <= n1009;
    \[6545]  <= n1014;
    \[6560]  <= n1019;
    \[6575]  <= n1024;
    \[6590]  <= n1029;
    \[6605]  <= n1034;
    \[6620]  <= n1039;
    \[6635]  <= n1044;
    \[6650]  <= n1049;
    \[6665]  <= n1054;
    \[6680]  <= n1059;
    \[6695]  <= n1064;
    \[6710]  <= n1069;
    \[6725]  <= n1074;
    \[6740]  <= n1079;
    \[6755]  <= n1084;
    \[6770]  <= n1089;
    \[6785]  <= n1094;
    \[6815]  <= n1099;
    \[6830]  <= n1104;
    \[6845]  <= n1109;
    \[6860]  <= n1114;
    \[6875]  <= n1119;
    \[6890]  <= n1124;
    \[6905]  <= n1129;
    \[6920]  <= n1134;
    \[6935]  <= n1139;
    \[6950]  <= n1144;
    \[6965]  <= n1149;
    \[6980]  <= n1154;
    \[6995]  <= n1159;
    \[7010]  <= n1164;
    \[7025]  <= n1169;
    \[7055]  <= n1174;
    ppeaks_12_12_ <= n1179;
    ppeaks_1_1_ <= n1183;
    ppeakp_3_3_ <= n1187;
    \[7115]  <= n1191;
    \[7130]  <= n1196;
    \[7145]  <= n1201;
    \[7160]  <= n1206;
    \[7175]  <= n1211;
    \[7190]  <= n1216;
    \[7205]  <= n1221;
    \[7220]  <= n1226;
    \[7235]  <= n1231;
    \[7250]  <= n1236;
    \[7265]  <= n1241;
    \[7280]  <= n1246;
    \[7295]  <= n1251;
    \[7310]  <= n1256;
    \[7325]  <= n1261;
    \[7340]  <= n1266;
    \[7355]  <= n1271;
    \[7370]  <= n1276;
    \[7385]  <= n1281;
    \[7400]  <= n1286;
    \[7415]  <= n1291;
    \[7430]  <= n1296;
    \[7445]  <= n1301;
    \[7460]  <= n1306;
    \[7475]  <= n1311;
    \[7490]  <= n1316;
    \[7505]  <= n1321;
    \[7520]  <= n1326;
    \[7535]  <= n1331;
    \[7550]  <= n1336;
    \[7565]  <= n1341;
    \[7580]  <= n1346;
    \[7595]  <= n1351;
    \[7625]  <= n1356;
    \[7640]  <= n1361;
    \[7655]  <= n1366;
    \[7670]  <= n1371;
    \[7685]  <= n1376;
    ppeaks_13_13_ <= n1381;
    ppeakp_7_7_ <= n1385;
    ppeakp_2_2_ <= n1389;
    \[7745]  <= n1393;
    \[7760]  <= n1398;
    \[7775]  <= n1403;
    \[7790]  <= n1408;
    \[7805]  <= n1413;
    \[7820]  <= n1418;
    \[7835]  <= n1423;
    \[7850]  <= n1428;
    \[7865]  <= n1433;
    \[7880]  <= n1438;
    \[7895]  <= n1443;
    \[7910]  <= n1448;
    \[7925]  <= n1453;
    \[7940]  <= n1458;
    \[7955]  <= n1463;
    \[7970]  <= n1468;
    \[8000]  <= n1473;
    \[8015]  <= n1478;
    \[8030]  <= n1483;
    \[8045]  <= n1488;
    \[8060]  <= n1493;
    \[8075]  <= n1498;
    \[8090]  <= n1503;
    \[8105]  <= n1508;
    \[8120]  <= n1513;
    \[8135]  <= n1518;
    \[8150]  <= n1523;
    \[8165]  <= n1528;
    \[8180]  <= n1533;
    \[8195]  <= n1538;
    \[8210]  <= n1543;
    \[8225]  <= n1548;
    \[8240]  <= n1553;
    \[8255]  <= n1558;
    \[8285]  <= n1563;
    \[8300]  <= n1568;
    \[8315]  <= n1573;
    \[8330]  <= n1578;
    ppeaks_3_3_ <= n1583;
    ppeakp_8_8_ <= n1587;
    ppeakp_1_1_ <= n1591;
    \[8390]  <= n1595;
    \[8405]  <= n1600;
    \[8420]  <= n1605;
    \[8435]  <= n1610;
    \[8450]  <= n1615;
    \[8465]  <= n1620;
    \[8480]  <= n1625;
    \[8495]  <= n1630;
    \[8510]  <= n1635;
    \[8525]  <= n1640;
    \[8540]  <= n1645;
    \[8555]  <= n1650;
    \[8570]  <= n1655;
    \[8585]  <= n1660;
    \[8600]  <= n1665;
    \[8615]  <= n1670;
    \[8630]  <= n1675;
    \[8645]  <= n1680;
    \[8660]  <= n1685;
    \[8675]  <= n1690;
    \[8690]  <= n1695;
    \[8705]  <= n1700;
    \[8720]  <= n1705;
    \[8735]  <= n1710;
    \[8750]  <= n1715;
    \[8765]  <= n1720;
    \[8780]  <= n1725;
    \[8810]  <= n1730;
    \[8825]  <= n1735;
    \[8840]  <= n1740;
    \[8855]  <= n1745;
    \[8870]  <= n1750;
    \[8885]  <= n1755;
    \[8900]  <= n1760;
    \[8915]  <= n1765;
    \[8930]  <= n1770;
    \[8945]  <= n1775;
    \[8960]  <= n1780;
    \[8975]  <= n1785;
    ppeaks_11_11_ <= n1790;
    ppeaks_2_2_ <= n1794;
    ppeakp_9_9_ <= n1798;
    ppeakp_0_0_ <= n1802;
    \[9050]  <= n1806;
    \[9065]  <= n1811;
    \[9080]  <= n1816;
    \[9095]  <= n1821;
    \[9110]  <= n1826;
    \[9125]  <= n1831;
    \[9140]  <= n1836;
    \[9155]  <= n1841;
    \[9170]  <= n1846;
    \[9185]  <= n1851;
    \[9200]  <= n1856;
    \[9215]  <= n1861;
    \[9230]  <= n1866;
    \[9245]  <= n1871;
    \[9260]  <= n1876;
    \[9275]  <= n1881;
    \[9290]  <= n1886;
    \[9305]  <= n1891;
    \[9320]  <= n1896;
    \[9335]  <= n1901;
    \[9350]  <= n1906;
    \[9365]  <= n1911;
    \[9380]  <= n1916;
    \[9395]  <= n1921;
    \[9410]  <= n1926;
    \[9440]  <= n1931;
    \[9455]  <= n1936;
    \[9470]  <= n1941;
    \[9485]  <= n1946;
    \[9500]  <= n1951;
    \[9515]  <= n1956;
    \[9530]  <= n1961;
    \[9545]  <= n1966;
    \[9560]  <= n1971;
    \[9575]  <= n1976;
    \[9590]  <= n1981;
    \[9605]  <= n1986;
    \[9620]  <= n1991;
    \[9635]  <= n1996;
    \[9650]  <= n2001;
    \[9665]  <= n2006;
    \[9680]  <= n2011;
    ppeaki_6_6_ <= n2016;
    \[9710]  <= n2020;
    \[9725]  <= n2025;
    \[9740]  <= n2030;
    \[9770]  <= n2035;
    \[9785]  <= n2040;
    \[9800]  <= n2045;
    \[9815]  <= n2050;
    \[9830]  <= n2055;
    \[9845]  <= n2060;
    \[9860]  <= n2065;
    \[9875]  <= n2070;
    \[9890]  <= n2075;
    \[9905]  <= n2080;
    \[9920]  <= n2085;
    \[9935]  <= n2090;
    \[9950]  <= n2095;
    \[9980]  <= n2100;
    \[9995]  <= n2105;
    \[10010]  <= n2110;
    \[10025]  <= n2115;
    \[10040]  <= n2120;
    \[10055]  <= n2125;
    \[10070]  <= n2130;
    \[10085]  <= n2135;
    \[10100]  <= n2140;
    \[10115]  <= n2145;
    \[10130]  <= n2150;
    \[10145]  <= n2155;
    \[10175]  <= n2160;
    \[10190]  <= n2165;
    \[10205]  <= n2170;
    \[10220]  <= n2175;
    ppeaki_15_15_ <= n2180;
    ppeaki_4_4_ <= n2184;
    \[10265]  <= n2188;
    \[10280]  <= n2193;
    \[10310]  <= n2198;
    \[10325]  <= n2203;
    \[10340]  <= n2208;
    \[10355]  <= n2213;
    \[10370]  <= n2218;
    \[10400]  <= n2223;
    \[10415]  <= n2228;
    \[10430]  <= n2233;
    \[10445]  <= n2238;
    \[10460]  <= n2243;
    \[10475]  <= n2248;
    \[10490]  <= n2253;
    \[10505]  <= n2258;
    ppeaki_14_14_ <= n2263;
    ppeaki_5_5_ <= n2267;
    \[10550]  <= n2271;
    \[10565]  <= n2276;
    \[10580]  <= n2281;
    \[10595]  <= n2286;
    \[10610]  <= n2291;
    \[10625]  <= n2296;
    \[10655]  <= n2301;
    \[10670]  <= n2306;
    \[10685]  <= n2311;
    \[10700]  <= n2316;
    \[10715]  <= n2321;
    \[10730]  <= n2326;
    \[10745]  <= n2331;
    \[10760]  <= n2336;
    \[10775]  <= n2341;
    \[10790]  <= n2346;
    \[10805]  <= n2351;
    \[10820]  <= n2356;
    \[10850]  <= n2361;
    \[10865]  <= n2366;
    \[10880]  <= n2371;
    \[10895]  <= n2376;
    \[10925]  <= n2381;
    \[10940]  <= n2386;
    \[10955]  <= n2391;
    \[10970]  <= n2396;
    \[10985]  <= n2401;
    \[11015]  <= n2406;
    \[11030]  <= n2411;
    \[11045]  <= n2416;
    \[11060]  <= n2421;
    \[11075]  <= n2426;
    \[11090]  <= n2431;
    \[11120]  <= n2436;
    \[11135]  <= n2441;
    \[11150]  <= n2446;
    \[11165]  <= n2451;
    \[11180]  <= n2456;
    \[11195]  <= n2461;
    \[11210]  <= n2466;
    \[11225]  <= n2471;
    \[11240]  <= n2476;
    \[11255]  <= n2481;
    \[11270]  <= n2486;
    \[11285]  <= n2491;
    \[11300]  <= n2496;
    \[11315]  <= n2501;
    \[11330]  <= n2506;
    \[11345]  <= n2511;
    \[11375]  <= n2516;
    \[11390]  <= n2521;
    \[11405]  <= n2526;
    \[11420]  <= n2531;
    \[11435]  <= n2536;
    \[11450]  <= n2541;
    \[11465]  <= n2546;
    \[11480]  <= n2551;
    \[11495]  <= n2556;
    \[11510]  <= n2561;
    \[11525]  <= n2566;
    \[11540]  <= n2571;
    \[11555]  <= n2576;
    \[11570]  <= n2581;
    \[11585]  <= n2586;
    \[11600]  <= n2591;
    \[11615]  <= n2596;
    \[11630]  <= n2601;
    \[11645]  <= n2606;
    \[11660]  <= n2611;
    \[11675]  <= n2616;
    \[11690]  <= n2621;
    \[11705]  <= n2626;
    \[11720]  <= n2631;
    \[11735]  <= n2636;
    \[11750]  <= n2641;
    \[11765]  <= n2646;
    \[11780]  <= n2651;
    \[11795]  <= n2656;
    \[11810]  <= n2661;
    ppeaki_9_9_ <= n2666;
    ppeakb_14_14_ <= n2670;
    \[11885]  <= n2674;
    \[11900]  <= n2679;
    \[11915]  <= n2684;
    \[11930]  <= n2689;
    ppeaki_8_8_ <= n2694;
    ppeakb_15_15_ <= n2698;
    \[12005]  <= n2702;
    \[12020]  <= n2707;
    \[12035]  <= n2712;
    \[12050]  <= n2717;
    \[12065]  <= n2722;
    \[12080]  <= n2727;
    ppeaki_7_7_ <= n2732;
    \[12125]  <= n2736;
    \[12140]  <= n2741;
    \[12155]  <= n2746;
    \[12170]  <= n2751;
    \[12185]  <= n2756;
    \[12200]  <= n2761;
    ppeakb_13_13_ <= n2766;
    \[12245]  <= n2770;
    \[12260]  <= n2775;
    \[12275]  <= n2780;
    ppeaki_13_13_ <= n2785;
    ppeaki_2_2_ <= n2789;
    \[12335]  <= n2793;
    \[12350]  <= n2798;
    \[12365]  <= n2803;
    \[12380]  <= n2808;
    \[12395]  <= n2813;
    \[12410]  <= n2818;
    \[12425]  <= n2823;
    \[12440]  <= n2828;
    \[12455]  <= n2833;
    \[12470]  <= n2838;
    \[12485]  <= n2843;
    ppeaki_12_12_ <= n2848;
    ppeaki_3_3_ <= n2852;
    \[12545]  <= n2856;
    \[12560]  <= n2861;
    \[12575]  <= n2866;
    \[12590]  <= n2871;
    \[12605]  <= n2876;
    \[12620]  <= n2881;
    \[12635]  <= n2886;
    \[12650]  <= n2891;
    \[12665]  <= n2896;
    \[12680]  <= n2901;
    \[12695]  <= n2906;
    ppeaki_11_11_ <= n2911;
    ppeaki_0_0_ <= n2915;
    \[12770]  <= n2919;
    \[12800]  <= n2924;
    \[12815]  <= n2929;
    \[12830]  <= n2934;
    \[12845]  <= n2939;
    \[12860]  <= n2944;
    \[12875]  <= n2949;
    \[12890]  <= n2954;
    \[12905]  <= n2959;
    \[12920]  <= n2964;
    \[12935]  <= n2969;
    ppeaki_10_10_ <= n2974;
    ppeaki_1_1_ <= n2978;
    \[13010]  <= n2982;
    \[13025]  <= n2987;
    \[13040]  <= n2992;
    \[13055]  <= n2997;
    \[13070]  <= n3002;
    \[13085]  <= n3007;
    \[13100]  <= n3012;
    \[13115]  <= n3017;
    \[13130]  <= n3022;
    \[13160]  <= n3027;
    \[13175]  <= n3032;
    ppeakb_4_4_ <= n3037;
    ppeaka_9_9_ <= n3041;
    \[13220]  <= n3045;
    \[13235]  <= n3050;
    \[13250]  <= n3055;
    \[13265]  <= n3060;
    \[13280]  <= n3065;
    \[13295]  <= n3070;
    \[13310]  <= n3075;
    \[13325]  <= n3080;
    \[13340]  <= n3085;
    \[13355]  <= n3090;
    \[13370]  <= n3095;
    \[13385]  <= n3100;
    \[13400]  <= n3105;
    \[13415]  <= n3110;
    \[13430]  <= n3115;
    \[13445]  <= n3120;
    \[13460]  <= n3125;
    \[13475]  <= n3130;
    \[13490]  <= n3135;
    \[13505]  <= n3140;
    ppeakb_5_5_ <= n3145;
    \[13550]  <= n3149;
    ppeakp_6_6_ <= n3154;
    \[13580]  <= n3158;
    \[13595]  <= n3163;
    \[13610]  <= n3168;
    \[13625]  <= n3173;
    \[13640]  <= n3178;
    \[13655]  <= n3183;
    \[13670]  <= n3188;
    \[13685]  <= n3193;
    \[13700]  <= n3198;
    \[13715]  <= n3203;
    \[13730]  <= n3208;
    \[13745]  <= n3213;
    \[13775]  <= n3218;
    \[13790]  <= n3223;
    \[13805]  <= n3228;
    \[13820]  <= n3233;
    \[13835]  <= n3238;
    \[13850]  <= n3243;
    \[13865]  <= n3248;
    \[13880]  <= n3253;
    \[13895]  <= n3258;
    ppeaka_11_11_ <= n3263;
    ppeaka_0_0_ <= n3267;
    ppeakp_5_5_ <= n3271;
    \[13955]  <= n3275;
    \[13970]  <= n3280;
    \[13985]  <= n3285;
    \[14000]  <= n3290;
    \[14015]  <= n3295;
    \[14030]  <= n3300;
    \[14045]  <= n3305;
    \[14060]  <= n3310;
    \[14075]  <= n3315;
    \[14090]  <= n3320;
    \[14105]  <= n3325;
    \[14120]  <= n3330;
    \[14135]  <= n3335;
    \[14150]  <= n3340;
    \[14165]  <= n3345;
    \[14180]  <= n3350;
    \[14210]  <= n3355;
    \[14225]  <= n3360;
    \[14240]  <= n3365;
    \[14255]  <= n3370;
    \[14270]  <= n3375;
    \[14285]  <= n3380;
    ppeakb_3_3_ <= n3385;
    ppeaka_10_10_ <= n3389;
    ppeaka_1_1_ <= n3393;
    ppeakp_4_4_ <= n3397;
    \[14360]  <= n3401;
    \[14375]  <= n3406;
    \[14390]  <= n3411;
    \[14405]  <= n3416;
    \[14420]  <= n3421;
    \[14435]  <= n3426;
    \[14450]  <= n3431;
    \[14465]  <= n3436;
    \[14480]  <= n3441;
    \[14495]  <= n3446;
    \[14510]  <= n3451;
    \[14525]  <= n3456;
    \[14540]  <= n3461;
    \[14555]  <= n3466;
    \[14570]  <= n3471;
    \[14585]  <= n3476;
    \[14600]  <= n3481;
    \[14615]  <= n3486;
    \[14630]  <= n3491;
    \[14660]  <= n3496;
    \[14675]  <= n3501;
    \[14690]  <= n3506;
    \[14705]  <= n3511;
    ppeakb_8_8_ <= n3516;
    ppeaka_13_13_ <= n3520;
    ppeaka_2_2_ <= n3524;
    \[14765]  <= n3528;
    ppeaks_9_9_ <= n3533;
    ppeakp_14_14_ <= n3537;
    \[14810]  <= n3541;
    \[14825]  <= n3546;
    \[14840]  <= n3551;
    \[14855]  <= n3556;
    \[14870]  <= n3561;
    \[14885]  <= n3566;
    \[14900]  <= n3571;
    \[14915]  <= n3576;
    \[14930]  <= n3581;
    \[14960]  <= n3586;
    \[14975]  <= n3591;
    \[14990]  <= n3596;
    \[15005]  <= n3601;
    \[15020]  <= n3606;
    \[15035]  <= n3611;
    \[15050]  <= n3616;
    \[15065]  <= n3621;
    \[15080]  <= n3626;
    ppeakb_9_9_ <= n3631;
    ppeaka_12_12_ <= n3635;
    ppeaka_3_3_ <= n3639;
    \[15140]  <= n3643;
    ppeaks_8_8_ <= n3648;
    ppeakp_15_15_ <= n3652;
    \[15185]  <= n3656;
    \[15200]  <= n3661;
    \[15215]  <= n3666;
    \[15230]  <= n3671;
    \[15245]  <= n3676;
    \[15260]  <= n3681;
    \[15275]  <= n3686;
    \[15290]  <= n3691;
    \[15305]  <= n3696;
    \[15320]  <= n3701;
    \[15335]  <= n3706;
    \[15350]  <= n3711;
    \[15365]  <= n3716;
    \[15380]  <= n3721;
    \[15395]  <= n3726;
    \[15410]  <= n3731;
    \[15425]  <= n3736;
    \[15440]  <= n3741;
    ppeakb_6_6_ <= n3746;
    ppeaka_15_15_ <= n3750;
    ppeaka_4_4_ <= n3754;
    \[15500]  <= n3758;
    \[15515]  <= n3763;
    ppeaks_0_0_ <= n3768;
    \[15545]  <= n3772;
    \[15560]  <= n3777;
    \[15575]  <= n3782;
    \[15590]  <= n3787;
    \[15605]  <= n3792;
    \[15620]  <= n3797;
    \[15635]  <= n3802;
    \[15650]  <= n3807;
    \[15665]  <= n3812;
    \[15680]  <= n3817;
    \[15695]  <= n3822;
    \[15710]  <= n3827;
    \[15725]  <= n3832;
    \[15755]  <= n3837;
    \[15770]  <= n3842;
    \[15785]  <= n3847;
    ppeakb_7_7_ <= n3852;
    ppeaka_14_14_ <= n3856;
    ppeaka_5_5_ <= n3860;
    \[15845]  <= n3864;
    \[15860]  <= n3869;
    ppeaks_10_10_ <= n3874;
    \[15890]  <= n3878;
    \[15905]  <= n3883;
    \[15920]  <= n3888;
    \[15935]  <= n3893;
    \[15950]  <= n3898;
    \[15965]  <= n3903;
    \[15980]  <= n3908;
    \[15995]  <= n3913;
    \[16010]  <= n3918;
    \[16025]  <= n3923;
    \[16040]  <= n3928;
    \[16055]  <= n3933;
    \[16070]  <= n3938;
    \[16085]  <= n3943;
    \[16100]  <= n3948;
    paddress_8_8_ <= n3953;
    \[16907]  <= n3957;
    \[16920]  <= n3962;
    \[16933]  <= n3967;
    paddress_9_9_ <= n3972;
    \[16959]  <= n3976;
    \[16972]  <= n3981;
    \[16985]  <= n3986;
    \[16998]  <= n3991;
    \[17011]  <= n3996;
    \[17024]  <= n4001;
    \[17037]  <= n4006;
    \[17050]  <= n4011;
    \[17063]  <= n4016;
    \[17076]  <= n4021;
    \[17089]  <= n4026;
    \[17102]  <= n4031;
    \[17115]  <= n4036;
    \[17128]  <= n4041;
    \[17141]  <= n4046;
    \[17154]  <= n4051;
    \[17167]  <= n4056;
    \[17180]  <= n4061;
    \[17193]  <= n4066;
    \[17206]  <= n4071;
    \[17219]  <= n4076;
    \[17232]  <= n4081;
    \[17245]  <= n4086;
    \[17258]  <= n4091;
    \[17271]  <= n4096;
    \[17284]  <= n4101;
    \[17297]  <= n4106;
    \[17310]  <= n4111;
    \[17323]  <= n4116;
    \[17336]  <= n4121;
    \[17349]  <= n4126;
    \[17362]  <= n4131;
    \[17375]  <= n4136;
    \[17388]  <= n4141;
    paddress_11_11_ <= n4146;
    \[17414]  <= n4150;
    \[17427]  <= n4155;
    \[17453]  <= n4160;
    paddress_10_10_ <= n4165;
    \[17479]  <= n4169;
    \[17492]  <= n4174;
    \[17505]  <= n4179;
    \[17518]  <= n4184;
    \[17531]  <= n4189;
    \[17544]  <= n4194;
    paddress_13_13_ <= n4199;
    \[17570]  <= n4203;
    \[17583]  <= n4208;
    \[17596]  <= n4213;
    \[17609]  <= n4218;
    paddress_12_12_ <= n4223;
    \[17635]  <= n4227;
    \[17648]  <= n4232;
    \[17661]  <= n4237;
    \[17674]  <= n4242;
    paddress_15_15_ <= n4247;
    \[17700]  <= n4251;
    \[17713]  <= n4256;
    paddress_14_14_ <= n4261;
    \[17739]  <= n4265;
    \[17752]  <= n4270;
    \[17765]  <= n4275;
    \[17778]  <= n4280;
    \[17791]  <= n4285;
    \[17804]  <= n4290;
    \[17817]  <= n4295;
    pwr_0_0_ <= n4300;
    \[17843]  <= n4304;
    \[17856]  <= n4309;
    \[17869]  <= n4314;
    \[17882]  <= n4319;
    prd_0_0_ <= n4324;
    \[17908]  <= n4328;
    \[17921]  <= n4333;
    \[17934]  <= n4338;
    \[17947]  <= n4343;
    \[17960]  <= n4348;
    \[17973]  <= n4353;
    \[17986]  <= n4358;
    \[17999]  <= n4363;
    \[18012]  <= n4368;
    \[18025]  <= n4373;
    \[18038]  <= n4378;
    pdn <= n4383;
    \[18064]  <= n4387;
    \[18077]  <= n4392;
    \[18090]  <= n4397;
    \[18103]  <= n4402;
    \[18116]  <= n4407;
    \[18129]  <= n4412;
    \[18142]  <= n4417;
    \[18155]  <= n4422;
    \[18168]  <= n4427;
    \[18181]  <= n4432;
    \[18194]  <= n4437;
    \[18207]  <= n4442;
    \[18220]  <= n4447;
    \[18233]  <= n4452;
    \[18246]  <= n4457;
    paddress_0_0_ <= n4462;
    piack_0_0_ <= n4466;
    \[18285]  <= n4470;
    \[18298]  <= n4475;
    \[18311]  <= n4480;
    paddress_1_1_ <= n4485;
    \[18337]  <= n4489;
    \[18350]  <= n4494;
    \[18363]  <= n4499;
    \[18376]  <= n4504;
    \[18389]  <= n4509;
    paddress_2_2_ <= n4514;
    \[18415]  <= n4518;
    \[18428]  <= n4523;
    \[18441]  <= n4528;
    paddress_3_3_ <= n4533;
    \[18467]  <= n4537;
    \[18480]  <= n4542;
    \[18493]  <= n4547;
    \[18506]  <= n4552;
    paddress_4_4_ <= n4557;
    paddress_5_5_ <= n4561;
    \[18545]  <= n4565;
    paddress_6_6_ <= n4570;
    \[18571]  <= n4574;
    \[18584]  <= n4579;
    \[18597]  <= n4584;
    \[18610]  <= n4589;
    paddress_7_7_ <= n4594;
    \[18636]  <= n4598;
  end
endmodule


